 "Ams	t->1	
 "Att	 ->1	
 "Big	 ->1	
 "Det	 ->4	
 "EU-	k->1	
 "Equ	a->1	
 "Eur	o->2	
 "Ja,	 ->1	
 "Kul	t->4	
 "Kvi	n->3	
 "Lot	h->1	
 "Min	d->1	
 "Mis	t->1	
 "Olj	e->1	
 "Om 	d->1	
 "Por	t->1	
 "Tib	e->2	
 "Ty 	h->1	
 "Urb	a->1	
 "aff	ä->1	
 "ald	r->2	
 "all	m->1	
 "ang	i->3	
 "avg	ö->1	
 "ban	k->1	
 "cou	p->1	
 "den	 ->3	
 "det	t->1	
 "död	a->1	
 "ege	n->1	
 "eko	l->1	
 "en 	e->1	l->1	w->1	
 "ent	r->1	
 "eur	o->3	
 "for	t->1	
 "för	"->1	
 "gem	e->1	
 "gen	d->1	
 "hel	l->1	
 "her	o->1	
 "in 	s->1	
 "inl	e->1	
 "irr	e->1	
 "ja 	t->1	
 "kol	l->2	
 "kro	n->1	
 "kul	t->1	
 "län	d->1	
 "läs	 ->2	
 "mel	l->1	
 "nat	u->1	
 "ne 	j->1	
 "nor	m->1	
 "någ	o->1	
 "obe	r->1	
 "orm	e->1	
 "ovi	l->1	
 "par	t->1	
 "påp	e->1	
 "ref	u->1	
 "res	t->1	u->3	
 "rik	t->1	
 "se 	p->1	
 "sha	l->1	
 "ska	d->1	
 "spe	c->1	
 "sva	g->1	
 "til	l->1	
 "utv	e->1	
 "utå	t->1	
 "val	u->1	
 "var	j->1	
 "åte	r->1	
 "öpp	e->1	
 "öve	r->1	
 'Vad	 ->1	
 ("di	e->1	
 (140	9->2	
 (199	8->2	
 (571	3->1	
 (809	5->2	
 (961	4->1	
 (A5-	0->35	
 (B5-	0->4	
 (Ben	e->1	
 (Bry	s->2	
 (C5-	0->7	
 (CEN	)->2	
 (CER	N->1	
 (COD	)->1	
 (DE)	 ->1	
 (EG,	 ->1	
 (EIF	)->1	
 (EL)	 ->1	
 (EN)	 ->23	
 (EU-	f->1	
 (EUG	F->2	
 (FI)	 ->1	
 (FIP	O->1	
 (FPÖ	)->1	
 (FR)	 ->12	
 (FUF	)->1	
 (H-0	0->1	7->12	8->8	
 (How	i->1	
 (ICE	S->1	
 (IFO	P->1	
 (IMO	)->1	
 (Int	e->1	
 (KOM	(->8	
 (Kul	t->2	
 (PPE	-->1	
 (PT)	 ->15	
 (SEK	(->1	
 (SPÖ	)->1	
 (Uts	k->2	
 (art	.->1	i->6	
 (att	 ->1	
 (avs	n->1	
 (de 	n->1	
 (det	 ->1	
 (eft	e->1	
 (ell	e->1	
 (en 	i->1	m->1	
 (fis	k->4	
 (for	t->1	
 (för	e->3	
 (häl	s->1	
 (i d	e->1	
 (i s	å->1	
 (inf	ö->1	
 (inr	e->1	
 (kod	i->2	
 (kom	m->1	
 (kon	s->1	
 (kri	s->2	
 (mai	n->2	
 (mer	 ->1	
 (och	 ->1	
 (rec	o->1	
 (råd	e->1	
 (se 	a->1	
 (sås	o->1	
 (t.e	x->1	
 (tyv	ä->1	
 (ung	.->1	
 (ÖVP	)->1	
 (Öst	e->4	
 (åte	r->1	
 , at	t->1	
 , bo	r->1	
 , de	t->1	
 , me	n->1	
 , vi	 ->1	
 - "d	e->1	
 - 'V	a->1	
 - , 	v->1	
 - 19	9->26	
 - 2,	8->1	
 - 31	 ->1	
 - 6 	m->1	
 - 80	 ->1	
 - Al	t->2	
 - C4	-->6	
 - C5	-->14	
 - Ca	m->1	
 - Do	m->1	
 - EU	-->1	
 - He	r->1	
 - Ka	l->1	
 - Ko	m->1	
 - Pa	r->1	
 - Re	v->1	
 - Ri	k->1	
 - Rå	d->1	
 - Sa	v->2	
 - al	l->5	
 - an	s->1	v->1	
 - ar	b->1	
 - at	t->27	
 - av	 ->9	
 - be	t->1	
 - bi	d->1	
 - bl	i->1	
 - bö	r->1	
 - ce	n->1	
 - de	 ->10	l->2	n->5	s->1	t->33	
 - do	c->1	
 - dv	s->2	
 - dä	r->2	
 - då	 ->2	
 - ef	t->2	
 - ek	o->1	
 - el	l->5	
 - en	 ->8	a->1	d->1	h->1	l->1	
 - et	t->3	
 - ev	e->1	
 - ex	e->1	i->1	
 - fa	t->1	
 - fi	c->1	
 - fr	a->1	ä->1	å->1	
 - få	 ->1	r->1	t->1	
 - fö	r->15	
 - ge	n->1	r->1	
 - gä	l->1	
 - gö	r->2	
 - ha	n->1	r->9	
 - ho	s->1	
 - hu	r->3	
 - hä	r->1	
 - i 	K->1	a->1	d->1	f->1	m->1	r->1	s->3	u->1	v->1	
 - id	a->1	
 - in	f->2	n->1	o->2	s->1	t->10	
 - ja	 ->1	,->2	g->12	
 - ju	s->1	
 - ka	n->1	
 - kn	a->1	
 - ko	m->6	n->1	s->2	
 - kr	ä->1	
 - li	k->1	n->1	
 - ly	s->1	
 - lå	t->2	
 - ma	n->2	r->1	
 - me	d->5	n->8	r->1	
 - mi	n->1	s->1	
 - mo	n->1	t->1	
 - må	n->1	s->1	
 - na	t->1	
 - ny	 ->1	
 - nä	m->3	r->3	
 - nå	g->6	
 - oc	h->61	k->1	
 - of	f->1	
 - om	 ->8	r->1	
 - or	d->1	
 - pa	r->1	
 - pr	e->1	i->1	
 - på	 ->4	m->1	
 - ra	p->1	
 - re	g->1	s->1	
 - ri	s->1	
 - rå	d->1	
 - rö	r->1	
 - sa	d->1	m->4	
 - se	 ->1	r->2	
 - si	t->1	
 - sk	a->2	u->1	
 - sn	a->1	e->1	
 - so	m->25	
 - st	a->2	o->1	
 - sy	f->1	s->1	
 - sä	g->1	r->1	
 - så	 ->5	l->1	
 - sö	k->1	
 - ta	c->1	
 - te	k->1	
 - ti	l->3	
 - tr	o->3	
 - tv	e->1	
 - tä	n->1	
 - un	d->1	
 - ut	a->7	g->1	s->1	t->1	
 - va	r->2	
 - ve	r->1	t->1	
 - vi	 ->6	k->1	l->10	s->1	
 - vä	l->1	
 - Ös	t->2	
 - är	 ->7	
 - äv	e->10	
 - åt	m->2	
 - öp	p->1	
 - öv	e->4	
 -(EN	)->1	
 -, a	t->1	
 -, d	ä->1	
 -, f	ö->1	
 -, i	 ->1	n->1	
 -, m	e->1	
 -, s	k->1	
 -, u	t->1	
 -, ä	r->1	
 -er 	r->1	
 -org	a->3	
 0 pr	o->1	
 000 	a->1	b->1	f->2	h->1	i->1	k->4	m->1	p->1	s->1	t->11	
 000.	M->1	
 008 	t->2	
 0113	 ->1	
 0550	 ->1	
 0652	 ->1	
 1 00	0->2	
 1 40	0->1	
 1 fr	å->1	
 1 i 	k->1	
 1 ja	n->5	
 1 ju	n->1	
 1 ma	r->2	
 1 me	n->1	
 1 oc	h->7	
 1 pr	o->4	
 1 se	p->1	
 1 ur	 ->1	
 1 ut	a->1	
 1, 2	 ->1	
 1, 4	,->1	
 1, a	t->1	
 1, o	c->1	
 1, s	k->1	
 1,2 	o->1	p->1	
 1,4 	t->1	
 1-2 	d->1	
 1-om	r->4	
 1-re	g->5	
 1-st	a->2	
 1.Ja	g->1	
 1/3 	a->1	
 10 0	0->2	
 10 e	l->1	
 10 j	a->1	
 10 k	a->1	
 10 m	i->2	
 10 p	r->4	
 10 r	i->1	
 10 s	o->1	
 10 ä	n->1	r->1	
 10 å	r->1	
 10, 	1->1	
 10.K	o->1	
 100 	d->1	k->1	m->1	o->1	p->1	ä->4	
 105 	i->1	t->1	
 11 i	 ->1	
 11 j	a->2	
 11 m	i->1	
 11 o	c->1	
 11 s	t->1	
 11, 	1->2	f->1	
 11,3	 ->1	
 11.0	0->3	
 11.A	l->1	
 11.E	x->1	
 11.K	u->1	
 110 	i->1	
 115 	m->1	
 12 f	r->1	
 12 i	n->1	
 12 j	a->1	
 12 m	i->1	å->1	
 12 o	c->1	
 12 p	r->1	
 12 s	t->1	
 12, 	1->2	d->1	t->1	
 12.0	0->6	
 12/9	9->3	
 120 	m->1	
 123 	p->1	
 1244	 ->1	.->2	
 125 	m->1	
 1260	/->1	
 13 (	E->1	
 13 0	0->1	
 13 A	m->1	
 13 f	e->1	
 13 i	 ->2	
 13 j	a->1	
 13 n	y->1	
 13 o	k->1	
 13 p	r->2	
 13 s	a->1	
 13 ä	r->1	
 13, 	2->2	
 13.0	5->1	
 13.F	ö->1	
 130 	d->1	
 133.	2->1	
 138.	4->1	
 14 f	e->5	
 14 m	e->5	
 14 o	c->1	
 14 s	e->1	
 14 t	i->1	
 14, 	e->1	
 140 	j->1	
 143 	o->1	
 15 a	v->1	
 15 m	a->1	
 15 o	l->2	m->1	
 15 p	r->3	
 15 r	ä->1	
 15 s	e->1	t->1	
 15 å	r->1	
 15, 	1->2	
 15.0	0->2	
 150 	g->1	o->1	
 158 	-->1	i->1	
 158)	.->1	
 158.	1->1	
 16 0	0->1	
 16 o	c->3	
 16 p	e->1	r->1	
 16 r	a->1	
 16) 	s->1	
 16, 	2->1	
 164 	r->1	
 166 	e->1	
 167 	m->3	
 17 d	e->2	
 17 m	i->1	
 17 o	k->1	
 17 s	å->1	
 17, 	1->1	s->1	
 17.3	0->1	
 17.S	l->1	
 170 	m->1	
 174 	t->1	
 1762	 ->1	.->1	
 18 d	e->1	
 18 h	ä->1	
 18 i	 ->1	
 18 m	i->1	å->1	
 18 n	o->3	
 18, 	2->1	
 180 	m->1	
 19 d	e->1	
 19 m	a->1	
 19 p	r->1	
 19 s	o->1	
 19 ä	r->1	
 19.5	0->1	
 1917	 ->1	
 1923	,->1	
 193 	o->1	
 1930	-->1	
 194.	D->1	
 1945	.->1	
 1948	.->1	
 195 	m->1	
 1957	 ->1	.->1	
 1967	 ->5	,->1	
 1969	 ->1	
 1976	 ->1	
 1977	 ->1	
 1982	,->1	.->1	
 1986	 ->2	.->1	
 1989	,->1	
 1990	 ->1	.->1	
 1991	 ->3	
 1992	 ->3	,->1	
 1993	 ->3	,->1	-->2	.->1	?->1	
 1994	 ->4	,->1	-->1	
 1995	 ->5	,->1	-->1	
 1996	 ->11	,->2	.->5	
 1997	 ->20	,->1	.->10	/->7	?->1	N->1	
 1998	 ->17	,->1	.->3	/->4	
 1999	 ->42	"->1	,->7	-->2	.->13	/->13	:->1	
 2 - 	v->1	
 2 00	0->1	
 2 40	0->1	
 2 bl	a->1	i->1	
 2 de	c->1	
 2 el	l->1	
 2 i 	a->2	r->1	s->1	
 2 mi	l->1	
 2 oc	h->3	
 2 pr	o->2	
 2 pu	n->1	
 2 so	m->1	
 2, 1	1->1	
 2, i	 ->1	
 2, s	k->1	o->1	
 2, v	i->1	
 2,48	7->1	
 2,6 	p->1	
 2,8 	m->1	
 2-om	r->2	
 2-st	ö->1	
 2.1 	i->1	
 2.2 	i->1	
 2.De	t->1	
 2.Me	n->1	
 20 0	0->1	
 20 e	u->1	
 20 g	å->1	
 20 m	i->2	
 20 n	y->1	
 20 p	r->3	
 20 º	 ->1	
 20 ä	n->1	
 20 å	r->5	
 20, 	2->1	
 20.2	5->1	
 200 	0->4	å->1	
 2000	 ->22	"->5	,->7	-->26	.->9	N->1	
 2001	 ->1	,->1	
 2002	 ->2	,->2	.->5	
 2003	?->1	
 2004	.->1	
 2006	 ->5	,->2	.->1	
 2007	,->1	
 2010	 ->1	
 2012	 ->1	
 21 j	a->1	u->1	
 21 o	c->1	m->1	
 21 s	t->1	
 21 ä	r->1	
 21 å	r->1	
 21.0	0->1	
 21.5	5->1	
 21:a	 ->1	
 22 a	v->1	
 22 r	i->1	
 22, 	2->1	i->1	v->1	
 22,5	 ->1	
 22.Ä	v->1	
 226 	i->1	
 23 d	e->1	
 23 i	n->1	
 23,7	 ->1	
 24 n	y->2	
 24 o	c->1	k->1	
 24 p	r->1	
 245 	o->1	
 248,	 ->1	
 25 g	r->1	
 25 m	e->1	i->1	
 25 o	m->1	
 25 p	r->7	
 25 t	i->1	
 25.D	e->1	
 250 	m->1	
 255 	i->4	
 26 "	p->1	
 26 i	n->1	
 26 m	e->1	
 26 n	o->1	
 26 o	c->1	
 26 p	r->1	
 262 	e->1	
 27 d	e->1	
 27 f	a->1	
 27 l	ä->1	
 27 o	c->1	
 27 p	r->2	
 27, 	3->1	
 28 f	r->1	
 28 j	u->1	
 28 n	y->1	
 28 p	r->1	
 28, 	3->2	
 280 	i->4	
 280.	4->1	
 28:e	 ->1	
 29 d	ö->1	
 29 f	r->1	
 29 l	ä->1	
 29 m	i->1	
 29, 	3->1	
 299.	2->2	
 3 00	0->2	
 3 fe	b->1	
 3 ja	n->1	
 3 ma	j->1	
 3 oc	h->1	
 3 ok	t->1	
 3 pr	o->1	
 3 pu	n->1	
 3, 7	,->1	
 3,8 	m->1	t->1	
 3-4 	p->1	
 3-li	t->2	
 3.1)	 ->1	
 3.8 	i->1	
 3.I 	ö->1	
 30 f	r->1	
 30 i	 ->1	n->1	
 30 j	u->1	
 30 m	e->1	i->1	
 30 o	c->1	
 30 p	r->3	
 30, 	3->1	
 300 	s->1	
 31 f	r->1	
 31 j	a->1	
 31 m	a->2	
 31 o	c->2	
 314 	l->1	
 32 m	i->1	
 32, 	3->2	
 32.J	a->1	
 33 0	0->2	
 33 a	v->1	
 33 f	r->1	ö->1	
 33 i	 ->1	
 33 o	c->1	
 332,	 ->1	
 34 i	 ->1	
 34 s	k->1	
 34 t	i->1	
 34 å	r->1	
 34, 	3->1	
 34.1	.->1	
 344 	-->1	
 35 f	r->1	
 35 m	i->5	
 35.S	å->1	
 350 	m->1	
 36 f	r->1	
 36, 	3->1	
 367 	0->1	
 37 f	r->1	
 37 i	 ->1	
 37 p	r->1	
 37, 	4->2	
 37.2	 ->1	
 37/6	0->1	
 370 	m->1	
 38 f	r->1	ö->1	
 38 o	c->2	
 38, 	4->1	
 38: 	f->1	
 39 f	r->1	
 39 i	 ->1	
 39 p	r->1	
 39, 	4->1	
 3: f	ö->1	
 4 00	0->1	
 4 c 	i->1	
 4 en	 ->1	
 4 i 	E->2	d->3	
 4 ju	n->2	
 4 li	k->1	
 4 oc	h->1	
 4 pr	o->1	
 4, 1	1->2	
 4, 6	,->1	
 4, o	c->1	
 4.2)	.->1	
 4.I 	d->2	
 4.Ja	g->1	
 40 f	r->1	
 40 m	i->1	
 40 p	r->6	
 40 å	r->3	
 40, 	4->1	
 400 	0->1	k->3	m->2	
 41 f	r->1	
 41 p	r->1	
 41 r	i->1	
 41 u	r->1	
 410 	f->1	
 42 f	r->1	
 42 i	 ->1	
 42 o	c->2	
 43 h	ö->1	
 43.F	r->1	
 44 f	r->1	
 44 o	c->2	
 45 a	v->1	
 45 c	e->1	
 45 f	r->1	
 45 g	ä->1	
 45, 	d->1	
 45. 	D->1	
 45."	I->1	
 45.H	e->1	
 45.V	i->1	
 46 o	c->2	
 462 	u->1	
 47 g	ä->1	
 48 g	ä->1	
 48 i	 ->2	n->1	
 48 ä	n->1	
 5 00	0->3	8->2	
 5 fr	å->1	
 5 gä	l->1	
 5 mi	l->3	
 5 ok	t->1	
 5 vi	s->1	
 5 år	.->1	
 5, d	ä->1	
 5, o	c->1	
 5, u	t->1	
 5,5 	p->1	
 5,8 	m->1	
 5.4 	i->1	
 5.Em	e->1	
 50 0	0->1	
 50 i	 ->1	
 50 m	i->2	
 50 p	r->3	
 50, 	s->1	
 50- 	o->1	
 50-t	a->2	
 500 	0->1	
 519 	-->1	
 52 i	 ->1	
 520 	-->1	f->1	
 522 	-->1	
 53 p	r->1	
 540 	m->1	
 55 m	o->1	
 55 p	r->1	
 56 p	r->1	
 56, 	s->1	
 57,5	 ->1	
 5b k	a->1	
 5b-o	m->1	
 5b.D	e->1	
 6 de	c->1	
 6 fr	å->1	
 6 i 	f->5	u->1	
 6 mi	l->1	
 6 oc	h->6	
 6 om	 ->1	
 6, 7	,->1	
 6, t	a->1	
 6,07	 ->1	
 6.Så	 ->1	
 60 0	0->1	
 60 f	r->1	
 60-t	a->1	
 600 	b->1	
 62 i	 ->1	
 67 i	 ->1	
 68 a	t->1	
 685/	9->1	
 7 - 	d->1	
 7 de	c->1	
 7 fö	r->1	
 7 gr	a->1	
 7 i 	A->2	b->1	d->1	f->3	v->1	
 7 le	d->1	
 7 nä	m->1	
 7 oc	h->2	
 7 pr	o->1	
 7 på	 ->1	
 7)..	 ->1	
 7, 9	,->1	
 7, d	v->1	
 7, o	c->1	m->1	
 7, s	o->1	
 7,2 	m->1	
 7,42	 ->1	
 7.Fr	å->1	
 70 a	n->1	
 70 p	r->1	
 700 	a->1	h->1	o->2	
 73,9	 ->1	
 75 -	 ->1	
 75 m	i->2	
 76 p	r->1	
 77 m	i->1	
 79/4	0->1	
 8 46	2->1	
 8 be	h->1	
 8 fr	å->1	
 8 oc	h->3	
 8 re	s->1	
 8 ti	l->1	
 8 är	 ->1	
 8, 9	,->1	
 8, s	å->1	
 80 e	n->1	
 80 p	r->11	
 80 ä	n->1	
 80 å	t->1	
 81 o	c->5	
 81 p	r->1	
 81.1	 ->3	.->2	
 81.3	 ->3	,->1	;->1	
 82 h	a->1	
 82 i	n->1	
 82) 	f->1	
 82, 	e->1	f->1	l->1	t->1	
 82.I	 ->1	
 83 p	r->1	
 85 o	c->2	
 85 p	r->1	
 85 t	i->1	
 86 i	 ->2	
 86 p	r->1	
 87, 	8->1	
 87.1	 ->1	
 87.2	 ->1	
 88 i	 ->1	
 88 o	c->1	
 88 ä	r->1	
 88/5	9->2	
 89 i	 ->1	
 89 t	i->1	
 9 de	c->1	
 9 fa	l->1	
 9 fe	b->1	
 9 fr	å->1	
 9 in	t->1	
 9 mi	l->3	
 9, a	n->1	
 9, f	ö->1	
 9.1 	v->1	
 90 d	e->1	ö->1	
 90 p	r->3	
 90-t	a->1	
 91 p	r->1	
 92/4	3->1	
 93 p	e->1	
 93/7	5->1	
 94 n	ä->1	
 94 p	r->2	
 94, 	k->1	
 94/5	5->2	
 94/7	2->1	
 95 i	 ->1	
 95 m	i->2	
 95 t	i->1	
 95/3	5->1	
 96/3	5->3	
 96/7	1->2	
 97.S	e->1	
 97/9	9->1	
 98 m	i->1	
 : Pa	r->1	
 A. G	u->1	
 ABB 	A->1	
 ABB-	A->2	
 ABC 	d->1	
 ADR)	 ->1	
 AKTU	E->1	
 Act.	 ->1	
 Adan	a->1	
 Aden	a->1	
 Adol	f->2	
 Adri	a->1	
 Afri	k->4	
 Agri	f->1	
 Agus	t->1	
 Aher	n->7	
 Aids	,->1	
 Akku	y->2	
 Akkö	y->1	
 Alav	a->2	
 Alba	c->1	n->1	
 Albe	r->1	
 Albr	i->1	
 Alex	a->2	
 Alge	r->1	
 Alic	a->1	
 Alla	 ->4	
 Allt	s->1	
 Alpe	r->1	
 Alsa	c->3	
 Alst	h->1	
 Alte	n->16	
 Amer	i->1	
 Amoc	o->1	
 Amok	o->5	
 Amos	 ->1	
 Amst	e->36	
 Ange	l->1	
 Anka	r->1	
 Anlä	g->1	
 Anmä	l->1	
 Anna	 ->1	
 Antó	n->1	
 Anve	r->1	
 Apar	i->1	
 Arab	r->1	
 Araf	a->1	
 Arbe	t->1	
 Ari 	V->1	
 Aria	n->3	
 Arti	k->1	
 Asie	n->2	
 Assa	d->2	
 Astu	r->1	
 Atat	u->1	ü->1	
 Atla	n->3	
 Att 	F->1	d->1	g->1	
 Ausc	h->1	
 Auto	/->1	
 Auve	r->1	
 Av d	e->1	
 Av o	m->1	
 Avfa	l->1	
 Avia	n->1	
 Avse	v->1	
 Azor	e->2	
 B oc	h->1	
 B ta	 ->1	
 BNI 	b->1	i->1	o->2	p->2	
 BNI,	 ->1	
 BNP 	j->1	m->1	p->4	å->1	
 BNP,	 ->2	
 BP, 	e->1	
 BRÅD	S->1	
 BSE 	o->2	
 BSE-	k->3	t->1	
 Balf	o->1	
 Balk	a->7	
 Bank	 ->1	
 Bara	k->9	
 Barc	e->2	
 Bare	n->1	
 Barn	h->1	i->14	
 Baró	n->2	
 Bask	i->2	
 Bass	e->1	
 Belg	i->9	
 Bere	n->12	
 Berg	 ->1	e->12	
 Berl	i->7	
 Bern	a->1	d->3	i->1	
 Bert	h->1	i->1	
 Besl	u->1	
 Besq	u->1	
 Betr	ä->1	
 Bisc	a->6	
 Blak	 ->1	
 Blan	d->1	
 Blok	 ->1	
 Boet	t->1	
 Bolk	e->1	
 Bond	e->1	
 Bord	e->1	
 Bort	o->1	
 Bour	l->6	
 Bowe	.->2	
 Bowi	s->2	
 Bran	d->2	
 Bras	i->1	
 Brav	e->1	
 Brem	e->1	
 Bret	a->7	
 Brit	i->1	
 Brok	 ->6	,->3	
 Brun	o->1	
 Brys	s->16	
 Buda	p->1	
 Bulg	a->1	
 Bush	,->1	
 Busq	u->1	
 Byrn	e->2	
 Byrå	n->1	
 C. D	e->1	
 C. E	f->1	
 C4-0	0->1	2->1	3->3	7->1	
 C5-0	0->6	1->5	3->4	
 CECA	F->1	
 CEN 	e->1	h->1	k->1	o->1	
 CEN,	 ->2	
 CEN:	s->4	
 CSU-	g->1	
 CSU:	s->1	
 Cadi	z->5	
 Cado	u->1	
 Camr	e->1	
 Camu	s->1	
 Cana	d->1	
 Cand	u->1	
 Cany	o->3	
 Casa	b->1	c->1	
 Caud	r->1	
 Cava	l->1	
 Cent	r->11	
 Cerm	i->1	
 Ceyh	u->1	
 Cham	p->1	
 Chiq	u->1	
 Clin	t->1	
 Coca	 ->1	
 Coci	l->1	
 Cola	,->1	
 Cona	k->1	
 Cons	t->1	
 Corb	e->1	
 Cost	a->9	
 Coun	c->1	
 Cox 	o->1	s->1	
 Cox!	J->1	
 Cox,	 ->1	
 Cres	p->2	
 Curi	e->1	
 Cusí	 ->1	
 Cuxh	a->1	
 Cype	r->1	
 D kr	ä->1	
 DDR.	S->1	
 Da C	o->3	
 Dage	n->1	
 Dagm	a->1	
 Dala	i->6	
 Dam 	b->1	s->1	
 Dama	s->1	
 Danm	a->25	
 Darm	s->1	
 Davi	d->3	
 De G	r->1	
 De P	a->1	
 De R	o->1	
 De d	a->1	i->1	
 De g	r->6	
 De h	a->1	
 De k	o->1	
 De n	o->1	
 De o	l->1	
 De s	o->2	t->1	
 De t	v->1	
 Delo	r->3	
 Demi	n->1	
 Demo	k->1	
 Den 	1->1	f->5	g->1	h->1	i->3	o->2	r->1	s->5	t->1	
 Denn	a->8	
 Dera	s->1	
 Dess	a->3	u->1	
 Det 	b->4	d->2	f->10	g->8	h->4	i->1	k->2	m->5	p->1	r->2	s->6	v->4	ä->25	å->1	
 Dett	a->13	
 Deut	s->1	
 Dimi	t->5	
 Dire	k->2	
 Doms	t->1	
 Dori	s->1	
 Dubl	i->7	
 Duha	m->1	
 Duis	e->3	
 Dutr	o->1	
 Där 	d->1	h->1	j->1	v->1	
 Däre	m->1	
 Därf	ö->2	
 Då b	ö->1	
 Då t	a->1	
 Díez	 ->1	
 Dühr	k->1	
 E-ko	l->1	
 ECHO	 ->1	,->1	.->1	
 EDD,	 ->1	
 EDD-	g->2	
 EEG 	t->1	
 EEG,	 ->2	
 EG t	i->1	
 EG-d	i->2	o->19	
 EG-f	ö->8	
 EG-k	o->16	
 EG-r	ä->3	
 EG.V	i->1	
 EG:s	 ->3	
 EIF 	h->1	
 EKSG	-->5	
 ELDR	 ->1	-->1	:->1	
 EMU,	 ->1	
 EMU-	a->1	k->1	
 EMU:	s->3	
 EU "	c->1	
 EU I	 ->1	
 EU a	g->1	t->2	
 EU b	l->1	ö->1	
 EU d	ä->1	
 EU f	r->1	
 EU g	e->1	ö->1	
 EU h	a->2	
 EU i	 ->1	n->3	
 EU k	a->3	
 EU m	e->1	y->1	
 EU o	c->4	
 EU p	å->1	
 EU r	e->1	
 EU s	k->1	o->4	y->1	
 EU u	t->2	
 EU ä	r->1	
 EU, 	f->1	l->1	m->1	p->1	v->1	
 EU-b	i->1	u->1	
 EU-e	n->1	
 EU-f	o->1	ö->4	
 EU-g	e->1	
 EU-i	n->5	
 EU-k	o->3	
 EU-l	a->2	ä->3	
 EU-m	a->1	e->5	
 EU-n	i->1	
 EU-p	r->2	
 EU-r	e->1	ä->1	
 EU-s	t->1	ä->2	
 EU-t	e->1	
 EU-u	t->1	
 EU-v	ä->1	
 EU..	 ->1	
 EU.A	l->1	
 EU.D	a->1	e->2	
 EU.F	r->1	
 EU.N	u->1	
 EU.R	o->1	
 EU.V	i->3	
 EU:s	 ->44	
 EU?H	e->1	
 EUGF	J->1	
 Ecem	i->1	
 Edin	b->1	
 Efta	r->2	
 Efte	r->9	
 Egyp	t->2	
 Ehud	 ->2	
 Eiec	k->1	
 Ekof	i->2	
 Ekon	o->1	
 Elis	a->1	
 Elle	s->3	
 Elma	r->2	
 Elst	.->1	
 Emil	i->1	
 En a	v->1	
 En b	e->1	
 En d	e->1	
 En p	e->1	r->1	
 En v	ä->1	
 Enda	s->1	
 Enli	g->5	
 Equa	l->7	
 Equq	a->2	
 Era 	t->1	
 Erik	a->24	
 Erit	r->1	
 Erkk	i->2	
 Ert 	b->1	
 Etio	p->3	
 Ett 	a->1	n->1	
 Eura	t->4	
 Euro	-->1	d->4	j->4	p->780	s->1	
 Evan	s->7	
 Exxo	n->3	
 FBI 	-->1	
 FEO 	b->1	ä->1	
 FMI 	d->1	
 FN, 	s->1	
 FN-u	p->1	
 FN.H	e->1	
 FN:s	 ->8	
 FPÖ 	(->2	f->1	i->1	m->1	o->3	s->1	v->1	
 FPÖ-	l->1	m->1	
 FPÖ:	s->2	
 FRÅG	O->1	
 Fact	o->1	
 Faro	u->1	
 Feir	a->2	
 Finl	a->6	
 Finn	s->1	
 Firm	a->1	
 Fisc	h->4	
 Flau	t->2	
 Flor	e->16	
 Fléc	h->1	
 FoU,	 ->1	
 FoU-	r->1	
 Fog 	f->1	
 Folk	f->1	r->2	
 Font	a->1	
 Ford	,->1	
 Fore	s->1	
 Frag	a->1	
 Fram	l->1	
 Fran	c->1	k->39	o->1	z->3	ç->1	
 Fras	s->1	
 Frih	e->2	
 Fru 	A->1	S->1	t->7	
 Frut	e->2	
 Främ	j->1	s->1	
 Fråg	a->2	
 Fund	 ->1	
 Fäst	n->1	
 Får 	j->2	
 Följ	a->1	
 För 	1->1	a->2	d->5	e->1	l->1	m->1	n->1	
 Förb	u->3	
 Före	n->40	
 Förh	i->1	
 Föri	n->2	
 Förs	l->1	t->10	ä->1	
 GA-s	t->1	
 GASP	 ->1	
 GUE/	N->2	
 GUSP	 ->1	
 Gale	o->1	
 Gali	c->2	
 Gama	 ->3	
 Garg	a->5	
 Gaza	 ->1	,->1	.->2	r->2	
 Geme	l->1	n->1	
 Gene	r->9	
 Geno	m->1	
 Genè	v->3	
 Gil-	D->1	R->1	
 Gino	,->1	
 Goeb	b->1	
 Gola	n->8	
 Golf	s->3	
 Goll	n->1	
 Gome	s->1	
 Gonz	á->1	
 Good	w->1	
 Gors	e->1	
 Gott	 ->1	
 Grac	a->3	o->1	
 Graç	a->5	
 Grek	l->12	
 Gros	s->3	
 Grup	p->8	
 Grön	a->1	i->1	
 Guat	e->1	
 Guig	o->1	
 Gulf	k->1	
 Gusp	"->1	
 Gute	r->2	
 Göte	b->1	
 Haar	d->1	
 Hade	r->1	
 Hagu	e->1	
 Haid	e->36	
 Hamb	u->1	
 Han 	k->1	
 Hand	i->1	
 Hans	 ->1	
 Har 	k->3	m->1	
 Hatz	i->2	
 Have	n->1	
 Hebr	o->1	
 Hedg	e->1	
 Hedk	v->1	
 Hein	z->1	
 Heli	g->1	
 Hels	i->20	
 Henr	y->1	
 Herr	 ->30	
 Hick	s->1	
 Hilt	o->1	
 Hima	l->1	
 Hitl	e->6	
 Hitt	i->1	
 Holl	y->1	
 Holz	m->2	
 Hon 	l->1	
 Huhn	e->1	
 Hult	e->18	h->6	
 Hur 	s->1	
 Häns	c->2	
 Här 	b->1	n->1	t->1	
 Håll	e->1	
 I - 	P->1	
 I Sc	h->1	
 I Tu	r->1	
 I be	t->1	
 I bu	d->1	
 I bö	r->2	
 I da	g->5	
 I de	n->3	t->3	
 I eg	e->3	
 I en	l->1	
 I gå	r->1	
 I li	k->1	
 I mo	r->1	t->1	
 I oc	h->2	
 I re	s->1	
 I si	t->1	
 I sl	u->1	
 I st	ä->1	
 I ut	s->1	
 I-pr	o->1	
 ICES	-->3	
 II -	 ->1	
 II h	a->1	
 II i	 ->1	
 II, 	h->1	
 II-p	r->2	
 III 	-->1	s->1	
 IMO.	D->1	
 IMO:	s->1	
 INTE	 ->1	R->3	
 IRA 	h->1	
 ISPA	-->1	
 IV -	 ->1	
 IV i	 ->2	
 IX o	c->1	
 IX, 	f->1	
 Ile-	d->1	
 Imbe	n->3	
 Indi	e->5	
 Inga	 ->1	
 Inge	n->1	r->1	t->1	
 Ingl	e->2	
 Init	i->1	
 Inte	 ->3	r->19	
 Irla	n->21	
 Isab	e->2	
 Isla	n->1	
 Isra	e->36	
 Ista	n->1	
 Ital	i->17	
 Izqu	i->1	
 Ja, 	h->1	v->1	
 Jack	s->1	
 Jaco	b->2	
 Jacq	u->2	
 Jag 	a->11	b->3	d->1	f->1	g->3	h->8	i->1	k->6	m->3	r->1	s->24	t->13	u->5	v->50	ä->9	ö->1	
 Jan-	K->1	
 Japa	n->3	
 Jave	t->1	
 Jean	-->1	
 Jeru	s->2	
 Jona	s->2	
 Jonc	k->13	
 Jord	a->2	b->1	
 Josp	i->1	
 Jugo	s->1	
 Junk	e->1	
 Jämf	ö->1	
 Jörg	 ->14	
 Kale	i->2	j->1	
 Kan 	r->1	
 Kana	d->1	
 Kant	a->3	
 Kara	s->3	
 Karl	 ->3	-->1	s->2	
 Kart	e->2	
 Kasp	i->1	
 Kauf	m->1	
 Kauk	a->3	
 Kaza	k->1	
 Kfor	 ->1	
 Kina	 ->7	,->1	.->1	s->1	
 Kinn	o->21	
 Kirg	i->5	
 Koch	 ->5	)->1	,->5	.->1	I->1	s->1	
 Komm	e->4	i->8	
 Konk	u->1	
 Konv	e->1	
 Kore	a->2	
 Koso	v->59	
 Kost	n->1	
 Kouc	h->12	
 Kult	u->11	
 Kuma	r->1	
 Kung	l->1	
 Kvin	n->1	
 Kväk	a->1	
 Kyot	o->7	
 Känn	e->1	
 Kära	 ->1	
 Kärn	k->1	t->1	
 Köln	 ->2	
 Köpe	n->1	
 LTCM	.->1	
 La R	é->1	
 Laan	 ->1	.->1	s->5	
 Lama	 ->3	.->2	s->2	
 Land	i->1	
 Lang	e->29	
 Lank	a->3	
 Lapp	l->2	
 Lead	e->5	
 Leda	m->1	
 Lein	e->6	s->2	
 Leon	i->1	
 Liba	n->5	
 Libe	r->2	
 Liby	e->1	
 Liik	a->3	
 Liks	o->2	
 Lill	e->1	
 Liss	a->8	
 Lita	u->1	
 Lloy	d->1	
 Loir	e->2	
 Lomé	a->1	k->1	
 Lond	o->4	
 Lord	 ->2	
 Lorr	a->2	
 Loth	a->2	
 Lous	e->1	
 Loyo	l->2	
 Lutt	e->1	
 Luxe	m->6	
 Lynn	e->3	
 Låt 	m->9	o->3	
 Lööw	 ->1	
 MARP	O->1	
 Maas	t->6	
 Maca	o->1	
 Mada	g->1	
 Made	i->2	
 Madr	i->3	
 Main	s->1	
 Malt	a->5	
 Man 	k->1	m->2	
 Marg	o->1	
 Mari	a->1	e->1	n->6	
 Mark	o->1	
 Marp	o->1	
 Mars	e->1	
 Mart	i->1	
 McCa	r->1	
 McNa	l->5	
 Med 	d->1	t->1	
 Mede	l->3	
 Mell	a->17	
 Men 	d->3	e->1	h->1	i->1	j->4	s->1	t->1	v->2	
 Men,	 ->1	
 Mexi	k->1	
 Mich	i->1	
 Midd	e->1	
 Midl	a->1	
 Min 	g->4	
 Mina	 ->1	
 Mini	s->1	
 Minu	c->1	
 Mist	e->1	
 Mitr	o->1	
 Mitt	 ->1	e->2	
 Mont	i->17	r->2	
 Mora	t->4	
 Morb	i->1	
 Morg	a->4	
 Mosk	v->1	
 Mour	a->8	
 Mous	k->1	
 Muld	e->1	
 Münc	h->1	
 Nana	 ->1	
 Napo	l->1	
 Nark	o->1	
 Nati	o->4	
 Nato	 ->1	a->1	b->1	s->2	
 Nede	r->9	
 Nej,	 ->1	
 New 	Y->1	
 Ni b	e->1	
 Ni h	a->3	
 Ni s	a->1	
 Ni v	i->1	
 Niel	s->5	
 Niki	t->2	
 Nogu	e->1	
 Noir	m->1	
 Nord	i->1	
 Norg	e->2	
 Nu f	å->1	
 Nya 	Z->2	
 Nytt	 ->1	
 När 	a->1	d->4	k->4	m->1	n->1	v->2	
 Näst	a->1	
 Någo	n->1	
 OCH 	B->1	
 OFSR	 ->1	
 OLAF	 ->5	,->5	.->4	:->1	
 OLFA	F->1	
 OM A	K->1	
 OSSE	 ->1	
 Ober	b->1	
 Och 	d->1	h->1	j->1	n->1	
 Och:	 ->1	
 Offe	n->1	
 Offi	c->1	
 Oil 	P->1	
 Oliv	i->1	
 Olje	t->1	
 Olym	p->1	
 Om E	U->1	
 Om i	n->1	
 Om m	a->1	
 Om n	å->1	
 Om o	m->1	
 Omag	h->1	
 Ones	t->1	
 Oran	i->1	
 Oslo	 ->1	,->2	
 Osma	n->1	
 Ouvr	i->1	
 Oz d	y->1	
 Oz, 	b->1	
 PPE 	h->1	ä->1	
 PPE-	D->5	g->5	
 PR-e	f->1	
 PSE)	J->1	
 PSE-	g->3	
 PVC,	 ->1	
 PVC-	l->1	
 PVC.	V->1	
 Pack	 ->2	s->1	
 Padd	i->2	
 Paki	s->5	
 Pala	c->15	
 Pale	r->1	s->10	
 Papa	y->2	
 Pari	s->3	
 Parl	a->4	
 Patt	e->23	
 Pays	 ->1	-->1	
 Peak	e->1	
 Peij	s->2	
 Peki	n->1	
 Pete	r->1	
 Petr	o->1	
 Plan	t->1	
 Plat	o->1	
 Ploo	i->1	
 Poet	t->5	
 Pohj	a->1	
 Pole	n->1	
 Poll	u->1	
 Pomé	s->1	
 Ponn	a->1	
 Poos	 ->1	
 Port	u->24	
 Powe	r->3	
 Preu	s->1	
 Prio	r->1	
 Proc	e->1	
 Prod	i->25	
 Prov	a->3	
 Prín	c->1	
 Purv	i->1	
 På d	e->2	
 På g	r->1	
 På s	a->1	
 Påst	å->1	
 Péta	i->1	
 Quec	e->1	
 REP 	(->1	r->1	
 RINA	 ->1	,->1	
 Rack	 ->1	,->1	
 Rafa	e->3	
 Rand	z->4	
 Rapk	a->11	
 Rasc	h->1	
 Read	i->1	
 Redi	n->8	
 Rege	r->1	
 Repu	b->1	
 Revi	d->1	s->1	
 Rhôn	e->1	
 Rich	a->1	t->2	
 Riis	-->2	
 Rikt	l->1	
 Riof	ö->1	
 Robe	r->1	
 Rois	s->1	
 Rojo	s->1	
 Rom-	 ->1	
 Roma	n->2	
 Romá	n->1	
 Roo 	f->1	
 Roth	-->5	
 Rott	e->2	
 Rove	r->2	
 Roya	l->1	
 Ruiz	 ->1	
 Rush	 ->1	
 Ryss	l->4	
 Råde	r->1	t->4	
 Råds	o->1	
 Réun	i->2	
 SEK 	(->1	
 SEK(	1->2	
 SEM-	2->1	
 SOLA	S->1	
 SPÖ 	o->1	
 SS o	c->1	
 Sage	s->1	
 Sain	t->1	
 Sala	f->1	
 Samm	a->15	
 San 	S->1	
 Sant	a->1	e->2	
 Save	 ->3	,->1	-->3	
 Sche	n->10	
 Schr	e->3	o->13	ö->1	
 Schu	l->2	
 Schw	a->1	e->1	
 Schö	r->1	
 Schü	s->3	
 Seat	t->4	
 Seba	s->1	
 Seda	n->4	
 Segn	i->1	
 Segu	r->1	
 Seix	a->5	
 Shar	m->5	
 Shel	l->2	
 Shep	h->3	
 Simp	s->1	
 Sjuk	h->1	
 Sjät	t->1	
 Sjös	t->4	
 Skog	s->1	
 Skot	t->4	
 Skul	l->1	
 Skäl	e->1	
 Slov	a->1	
 Soar	e->1	
 Soci	a->1	
 Sokr	a->1	
 Sola	n->4	
 Solb	e->2	
 Som 	T->1	e->2	j->1	n->3	t->1	v->1	
 Soul	a->1	
 Span	i->7	
 Spen	c->1	
 Sper	o->1	
 Sri 	L->3	
 St.V	a->1	
 Stad	g->1	
 Stat	e->1	
 Stoc	k->3	
 Stor	b->14	
 Stra	s->5	x->1	
 Stöd	 ->1	
 Suan	z->1	
 Sudr	e->2	
 Sver	i->7	
 Swob	o->3	
 Syda	f->2	
 Sydk	o->1	
 Sydo	s->2	
 Syri	e->22	
 Sánc	h->1	
 São 	T->2	
 Så l	å->1	
 Så r	i->1	
 Söde	r->2	
 TV a	n->1	
 TV-k	a->1	
 TV-p	r->1	
 TV-s	ä->1	
 Taci	s->2	
 Tack	 ->7	
 Tadz	j->4	
 Taiw	a->1	
 Talm	a->1	
 Tamm	e->22	
 Tang	 ->1	
 Tani	o->1	
 Taue	r->1	
 Terr	ó->3	
 Tesa	u->1	
 Texa	s->2	
 Thea	t->19	
 Thys	s->4	
 Tibe	t->19	
 Tidn	i->1	
 Till	 ->5	å->3	
 Todi	n->1	
 Tom 	S->1	
 Tomé	 ->2	
 Torr	e->3	
 Tota	l->6	
 Tran	s->1	
 Tred	j->1	
 Trit	t->1	
 Trot	s->1	
 Tsat	s->3	
 Turk	i->35	m->2	
 Tysk	l->20	
 Tågk	r->1	
 UCK 	n->1	
 UCLA	F->1	
 UEN-	g->1	
 UNIF	I->1	
 UNMI	K->3	
 USA 	-->1	a->1	e->1	h->1	p->1	
 USA,	 ->2	
 USA.	J->1	V->1	
 USA:	s->1	
 USD 	f->1	
 Ulst	e->1	
 Unde	r->6	
 Unio	n->3	
 Uppd	a->1	
 Urba	-->1	
 Urqu	i->1	
 Ursä	k->1	
 Utnä	m->1	
 Utsk	o->2	
 Utvä	r->1	
 Uzbe	k->2	
 V - 	R->1	
 VD b	ö->1	
 VI i	 ->1	
 VIII	 ->2	
 Vad 	b->3	g->1	j->2	v->1	ä->2	
 Vald	e->3	
 Vall	e->3	
 Van 	H->2	
 Vand	a->1	
 Vape	n->1	
 Vare	l->1	
 Varf	ö->1	
 Varj	e->2	
 Vark	e->1	
 Vata	n->3	
 Velz	e->1	
 Vem 	b->1	s->2	
 Vend	é->1	
 Vene	z->1	
 Vens	t->2	
 Verh	e->2	
 Vers	a->1	
 Vi b	e->1	
 Vi f	å->3	ö->3	
 Vi h	a->9	å->1	
 Vi k	a->1	o->2	ä->1	
 Vi m	i->1	å->2	
 Vi s	k->2	t->2	
 Vi u	t->1	
 Vi v	a->2	i->3	ä->2	
 Vi ä	r->3	
 Vi, 	d->1	
 Vich	y->1	
 Vid 	d->1	e->1	
 Vilk	a->1	
 Viss	a->1	
 Vito	r->7	
 Vivi	e->1	
 Vlaa	m->1	
 Voda	f->1	
 Volk	s->1	
 Värl	d->3	
 Väst	b->4	
 Vår 	d->1	u->1	
 Våra	 ->1	
 Vårt	 ->2	
 WTO?	E->1	
 Waff	e->2	
 Wale	s->11	
 Wall	s->4	
 Wash	i->3	
 Web,	 ->1	
 West	 ->1	
 Wide	 ->1	
 Wieb	e->1	
 Wiel	a->4	
 Wien	 ->3	,->1	
 Wilh	e->1	
 Woga	u->18	
 Wulf	-->2	
 Wurt	z->3	
 Wye 	P->1	
 Wye-	a->2	
 Wynn	,->1	
 X oc	h->1	
 XXVI	I->2	
 Yass	e->1	
 York	 ->1	
 Zeel	a->2	
 Zime	r->1	
 [KOM	(->2	
 [SEK	(->1	
 a pr	i->3	
 a) a	d->1	
 a) b	ä->1	
 abso	l->40	r->1	
 abst	r->1	
 absu	r->3	
 acce	p->57	
 acqu	i->1	
 ad h	o->2	
 ad i	n->1	
 addi	t->1	
 adek	v->5	
 adje	k->2	
 admi	n->23	
 adri	a->1	
 advo	k->5	
 affä	r->4	
 agen	d->1	
 ager	a->42	
 aggr	e->1	
 agit	a->1	
 agra	r->1	
 agro	t->1	
 aids	 ->2	-->1	p->2	
 ajou	r->1	
 akt 	a->2	o->2	p->2	u->1	
 akta	 ->3	t->1	
 akte	n->1	
 akti	e->3	o->2	v->22	
 aktu	a->1	e->30	
 aktö	r->10	
 akut	a->1	
 al-S	h->1	
 alba	n->9	
 aldr	i->29	
 alib	i->1	
 alke	m->1	
 alko	h->1	r->1	
 all 	E->1	a->1	d->3	e->1	f->2	g->1	h->1	k->3	m->2	o->2	p->3	r->6	s->4	t->3	u->1	v->2	
 alla	 ->347	!->1	,->5	.->4	s->5	
 alld	e->22	
 alle	g->1	h->3	n->1	s->5	u->2	
 alli	a->7	e->1	h->1	
 allm	o->1	ä->120	
 allo	k->1	
 allr	a->9	
 alls	 ->14	,->1	.->2	i->1	
 allt	 ->165	,->6	.->3	:->1	f->39	i->83	j->3	m->1	s->63	
 allv	a->74	
 alta	r->1	
 alte	r->11	
 amba	s->1	
 ambi	t->26	
 ambu	l->1	
 amer	i->11	
 an a	t->3	
 an d	e->2	
 an f	r->2	
 an p	å->1	
 an t	i->1	
 an å	t->1	
 ana 	a->1	d->1	e->1	g->1	
 anal	y->43	
 anam	m->4	
 anbl	i->1	
 anbu	d->4	
 and 	a->1	
 anda	 ->5	.->3	n->3	s->1	
 ande	l->7	m->5	
 andl	i->1	
 andr	a->313	e->1	
 anfö	r->16	
 anga	v->1	
 ange	 ->4	l->21	n->1	r->3	s->2	
 angi	v->2	
 angr	e->6	i->7	ä->1	
 angå	e->26	r->2	
 anhä	n->4	
 anin	g->5	
 ankl	a->3	
 ankn	y->1	
 anko	m->1	
 anle	d->48	
 anli	t->1	
 anlä	g->4	n->1	
 anlö	p->4	
 anmä	l->18	r->10	
 anna	n->43	r->15	t->69	
 anno	r->4	
 anon	y->4	
 anor	d->8	
 anpa	s->12	
 ansa	t->5	
 anse	 ->1	.->1	e->2	n->1	r->192	s->5	t->2	
 ansi	k->1	
 ansj	o->17	
 ansk	a->1	r->1	
 ansl	a->15	o->1	u->26	å->4	
 ansp	e->1	r->5	
 anst	r->44	ä->31	
 ansv	a->276	
 anså	g->12	
 ansö	k->10	
 anta	 ->23	g->35	l->58	r->9	s->10	
 ante	 ->2	,->2	
 anti	-->3	b->1	d->1	e->1	f->4	k->4	m->1	n->10	s->3	t->1	
 anto	g->23	
 anty	d->2	
 anvi	s->1	
 anvä	n->158	
 appa	r->1	
 appe	l->1	
 appl	å->6	
 apri	l->3	
 apro	p->1	
 arab	i->6	s->2	
 arbe	t->407	
 argu	m->16	
 arki	v->2	
 armo	d->1	
 armé	 ->1	n->2	
 arra	n->6	
 arre	s->2	
 arro	g->2	
 art 	o->1	
 art.	D->1	V->1	
 arte	n->1	r->1	
 arti	f->2	g->1	k->98	
 arto	n->1	
 arv.	"->1	B->1	
 arve	t->2	
 as".	J->1	
 aspe	k->30	
 assi	s->2	
 asso	c->1	
 astr	o->1	
 asyl	 ->4	,->2	-->1	.->3	b->1	f->2	r->2	s->6	
 atla	n->1	
 atom	e->3	f->1	
 att 	"->1	-->6	1->3	2->1	4->1	7->1	8->1	A->3	B->5	C->1	D->3	E->90	F->5	G->1	I->6	J->3	K->2	M->2	N->1	O->3	P->3	R->3	S->3	T->16	V->1	a->210	b->306	c->1	d->1067	e->146	f->468	g->296	h->173	i->196	j->91	k->318	l->147	m->349	n->102	o->76	p->141	r->150	s->460	t->243	u->258	v->567	y->6	z->1	ä->62	å->54	ö->68	
 att,	 ->8	
 att.	.->1	
 att:	 ->1	
 atta	c->1	
 atte	n->4	
 atti	t->5	
 attr	a->1	
 auct	o->1	
 aukt	o->6	
 auto	m->8	p->1	
 av "	p->1	r->2	
 av -	 ->5	
 av 1	4->1	9->3	
 av 2	0->1	
 av 5	 ->1	4->1	
 av A	h->2	m->2	r->1	
 av B	N->6	S->1	a->2	e->8	o->1	r->2	
 av C	a->1	
 av D	a->2	e->1	i->2	u->1	ü->1	
 av E	G->1	U->17	r->1	u->70	x->2	
 av F	N->1	P->2	l->1	ö->8	
 av G	a->1	e->2	r->3	
 av H	a->1	e->1	i->1	
 av I	s->2	
 av J	a->1	e->1	o->2	
 av K	i->2	o->10	u->1	
 av L	a->3	i->1	ö->1	
 av M	a->2	c->1	o->1	
 av O	L->3	s->1	z->1	
 av P	a->2	o->1	é->1	
 av R	a->1	i->1	
 av S	a->1	c->6	
 av T	a->1	e->1	h->4	i->1	o->1	
 av U	N->1	
 av V	a->2	ä->1	
 av W	a->1	i->1	y->1	
 av a	c->1	d->2	g->1	l->32	n->26	p->2	r->39	s->1	t->64	v->9	
 av b	a->2	e->37	i->14	l->3	o->3	r->10	u->8	y->2	å->2	ö->3	
 av c	e->2	i->6	o->1	
 av d	a->5	e->542	i->26	j->1	o->12	r->1	
 av e	f->3	g->2	k->10	n->109	r->18	t->51	u->7	v->1	x->8	
 av f	a->47	i->6	j->2	l->16	o->8	r->25	u->5	y->1	ä->1	å->2	ö->104	
 av g	a->3	e->31	i->3	l->1	o->1	r->11	
 av h	a->10	e->7	i->5	u->8	ä->1	ö->2	
 av i	 ->3	b->1	c->3	d->2	m->4	n->26	
 av j	o->5	u->4	ä->2	
 av k	a->10	l->4	n->1	o->109	r->5	u->5	v->5	ä->8	
 av l	a->19	e->10	i->13	o->5	ä->4	å->1	ö->1	
 av m	a->17	e->26	i->37	o->5	y->3	ä->7	å->7	ö->1	
 av n	a->14	i->1	o->1	y->11	ä->1	å->5	ö->2	
 av o	a->2	b->2	c->3	f->5	k->1	l->14	m->9	n->1	r->10	s->12	t->2	u->1	v->1	
 av p	a->22	e->12	i->1	o->8	r->36	
 av r	a->6	e->32	i->7	y->1	ä->12	å->12	ö->1	
 av s	a->12	c->1	e->7	i->23	j->3	k->18	l->2	m->2	o->8	p->2	t->72	u->4	v->2	y->20	ä->14	å->10	
 av t	a->2	e->8	i->12	j->28	o->2	r->11	u->6	v->1	y->2	ä->1	
 av u	n->27	p->4	t->33	
 av v	a->22	e->8	i->19	o->4	ä->18	å->24	
 av y	t->5	
 av Ö	s->2	
 av ä	l->1	m->1	n->5	r->1	
 av å	l->1	r->7	s->1	t->14	
 av ö	b->1	d->1	k->3	p->4	s->2	v->3	
 av, 	o->2	s->1	t->1	ä->1	
 av.D	e->2	ä->1	
 av.E	f->1	
 av.J	a->1	
 av.M	e->1	
 av.O	L->1	
 avan	c->1	t->1	
 avbr	o->2	y->3	ö->6	
 avde	l->8	
 avec	 ->1	
 aveu	r->1	
 avfa	l->22	
 avfo	l->1	
 avfö	r->3	
 avga	s->1	v->1	
 avge	 ->3	r->5	s->1	t->1	
 avgi	c->4	f->1	v->1	
 avgj	o->4	
 avgr	ä->3	
 avgå	.->1	e->1	n->1	r->1	t->1	
 avgö	r->55	
 avhj	ä->2	
 avhä	n->2	
 avhå	l->1	
 avis	e->4	
 avkl	a->1	
 avkr	ä->1	
 avku	n->1	
 avla	d->1	g->1	
 avle	d->2	
 avli	v->1	
 avlo	p->1	
 avlä	g->10	
 avma	t->1	
 avpr	i->1	
 avra	p->1	
 avre	g->2	
 avru	n->1	
 avrä	t->1	
 avsa	k->4	t->3	
 avse	 ->1	d->3	e->47	r->14	s->1	t->4	v->13	
 avsi	d->1	k->36	
 avsk	a->19	e->5	i->1	r->2	y->2	
 avsl	a->2	o->2	u->60	ä->1	å->3	ö->6	
 avsn	i->3	
 avsp	e->5	
 avst	a->1	o->2	ä->3	å->26	
 avsä	g->1	t->4	
 avta	l->54	r->1	
 avtv	i->1	
 avun	d->1	
 avva	k->6	
 avve	c->8	r->1	
 avvi	k->8	s->14	
 avvä	g->3	
 axel	r->1	
 axla	r->1	
 b) i	n->1	
 b) m	i->1	
 baci	l->1	
 back	-->1	
 bad 	F->1	e->1	k->1	o->1	
 bada	 ->1	
 baga	t->2	
 bain	"->1	
 bak 	i->1	
 bakd	ö->1	
 bakg	r->31	
 bako	m->21	
 bakå	t->3	
 bala	n->25	
 bana	l->3	n->1	t->1	
 banb	r->1	
 band	 ->2	e->2	
 bank	 ->1	e->1	f->1	i->1	s->1	
 bann	l->1	
 bano	r->2	
 bant	a->1	n->1	
 bar 	g->1	
 bara	 ->226	,->1	:->1	
 barb	a->2	
 bark	b->1	
 barn	 ->5	,->3	b->1	p->2	s->1	
 barr	i->2	
 bart	 ->1	
 bas 	f->1	i->1	
 bas,	 ->1	
 basa	r->2	
 base	b->1	n->2	r->7	
 basi	s->3	
 bask	i->4	r->1	
 bast	u->1	
 baxa	 ->1	
 be P	r->1	
 be e	r->5	
 be f	r->1	
 be h	e->1	o->1	
 be k	o->6	
 be o	m->2	
 be p	a->1	
 be s	t->1	
 beak	t->30	
 bear	b->2	
 beby	g->1	
 bebå	d->1	
 bedr	e->1	i->15	ä->32	
 bedö	m->44	
 befa	r->5	t->6	
 befi	n->41	
 befl	ä->1	
 befo	g->28	l->39	r->5	
 befr	a->9	i->3	ä->1	
 befä	l->1	n->1	s->10	
 bega	g->4	
 begr	a->1	e->12	i->5	u->2	ä->63	
 begä	r->60	
 begå	 ->2	r->3	s->3	t->3	
 beha	n->73	
 beho	v->65	
 behä	f->1	
 behå	l->12	
 behö	l->1	r->18	v->147	
 beiv	r->1	
 beka	n->3	
 bekl	a->42	
 beko	m->1	s->1	
 bekr	ä->30	
 bekv	ä->15	
 beky	m->16	
 bekä	m->33	n->1	
 bela	s->6	
 belg	i->8	
 belo	p->11	
 bely	s->4	
 belä	g->5	
 belö	n->2	
 bema	n->1	
 bemy	n->1	
 bemä	r->5	
 bemö	d->3	t->7	
 bene	n->1	
 benh	å->1	
 bens	i->1	
 benä	g->1	
 benå	d->1	
 beor	d->1	
 ber 	V->1	a->3	d->2	e->7	f->1	i->1	j->9	k->4	n->1	o->8	r->1	
 ber,	 ->1	
 bere	d->34	t->4	
 beri	k->8	
 bero	d->5	e->15	r->19	t->1	
 bery	k->1	
 berä	k->3	t->28	
 berö	m->2	r->42	v->1	
 bese	g->2	
 besi	k->2	t->2	
 besk	a->3	e->3	r->22	y->4	
 besl	u->196	ä->1	ö->1	
 besp	a->2	
 best	o->1	r->4	y->1	ä->127	å->39	ö->1	
 besv	a->14	i->8	ä->7	
 besy	n->1	
 besä	t->2	
 besö	k->8	
 beta	l->68	
 bete	c->4	e->3	r->1	
 betj	ä->1	
 beto	n->44	
 betr	a->23	y->1	ä->72	
 bett	 ->2	
 betu	n->1	
 betv	i->3	
 bety	d->122	
 betä	n->248	
 beun	d->3	
 beva	k->5	r->21	
 beve	k->1	
 bevi	l->48	s->37	t->1	
 bibe	h->11	
 bibl	i->2	
 bidr	a->106	o->3	
 bief	f->2	
 bifa	l->3	
 bigo	t->1	
 bil 	e->1	f->1	g->1	i->1	k->1	s->4	v->1	
 bil,	 ->2	
 bil-	 ->1	
 bil.	 ->1	D->1	T->1	
 bila	g->6	r->71	t->6	
 bilb	e->1	r->1	
 bild	 ->4	.->2	a->20	e->5	
 bile	n->6	
 bili	n->29	s->1	
 bilj	o->1	
 bilk	o->1	y->1	ö->2	
 bill	i->6	
 bilm	ä->1	
 bilp	a->6	r->1	
 bils	 ->2	e->1	k->2	
 bilt	i->15	
 bilv	r->6	
 bilä	g->1	
 bilå	t->1	
 bind	a->12	e->2	
 bio 	s->1	
 biol	o->4	
 biop	l->1	
 bios	f->1	ä->2	
 bist	å->20	
 bit 	p->1	
 bite	r->1	
 bitt	e->2	r->1	
 bjud	a->1	e->1	
 bl.a	.->27	
 blam	e->1	
 blan	d->54	k->2	
 blek	a->1	
 blev	 ->14	
 bli 	2->1	a->11	b->4	d->5	e->28	f->12	g->1	h->1	j->1	k->4	l->3	m->21	n->5	o->3	p->3	r->1	s->8	t->3	v->3	ä->1	ö->2	
 bli,	 ->1	
 bli.	U->1	
 blic	k->2	
 blin	d->1	t->1	
 blir	 ->106	,->2	:->1	
 bliv	a->1	i->26	
 blix	t->1	
 bloc	k->4	
 blom	m->3	s->3	
 blot	t->3	
 blun	d->4	
 bly 	å->1	
 bly,	 ->2	
 bly.	V->1	
 blyg	s->4	
 blå 	b->1	
 bo i	 ->1	
 bo k	v->1	
 boen	d->1	
 bogs	e->1	
 bojk	o->1	
 bok 	a->1	o->1	t->1	
 boks	l->1	t->1	
 bola	g->5	
 bomb	 ->1	.->1	a->2	e->4	n->1	
 bomu	l->1	
 bond	g->2	
 bor 	d->1	i->4	p->1	
 bord	 ->1	.->1	e->68	l->1	
 borg	a->1	m->2	
 bort	 ->20	,->5	.->6	a->1	f->6	o->2	p->1	s->6	
 bosa	t->3	
 bosn	i->2	
 bost	a->1	ä->4	
 bosä	t->4	
 bot 	p->2	
 bota	r->2	
 bott	e->5	n->4	
 bova	r->1	
 bove	n->1	
 bra 	a->11	b->5	d->5	e->2	f->3	i->3	j->1	m->5	n->2	o->9	s->9	t->1	u->4	v->1	ä->2	å->1	
 bra!	M->1	
 bra,	 ->8	
 bra.	D->1	E->1	J->1	P->1	S->1	V->1	
 bran	d->3	s->5	
 bred	 ->4	a->6	d->2	e->1	
 bret	a->1	t->6	
 brev	 ->4	.->1	l->1	
 brie	f->1	
 brin	g->3	
 bris	t->60	
 brit	t->16	
 bro 	m->1	
 broa	r->1	
 brod	e->2	
 brok	i->2	
 brom	e->4	s->6	
 bror	,->1	
 brot	h->1	t->40	u->1	
 bruk	 ->1	,->2	a->3	e->1	
 brun	a->1	
 brut	a->1	i->2	t->1	
 bryr	 ->2	
 bryt	a->7	e->3	n->2	
 brän	d->2	n->3	s->7	
 bräs	c->2	
 bråd	s->20	
 bråk	e->1	
 bröd	.->2	
 brös	t->1	
 bröt	 ->1	
 budd	h->1	
 budg	e->102	
 budo	r->1	
 buds	k->10	
 buri	t->1	
 buss	a->1	
 bygg	a->29	d->2	e->10	n->3	s->3	t->3	
 byrå	 ->2	e->1	k->29	n->2	
 byta	 ->1	
 byte	t->1	
 bytt	s->1	
 byxf	i->1	
 bär 	a->5	b->1	d->1	f->2	l->1	p->3	s->1	u->1	v->1	
 bära	 ->9	s->3	
 bärs	 ->2	
 bäst	 ->5	a->37	
 bätt	r->75	
 båda	 ->22	,->1	
 både	 ->46	
 båta	r->8	
 båte	n->1	
 bébé	 ->1	
 böck	e->3	
 böde	l->1	
 böje	l->1	
 böjt	 ->1	
 bör 	"->1	-->1	E->3	a->10	b->8	d->16	e->5	f->18	g->12	h->6	i->14	k->7	l->6	m->24	n->4	o->6	s->10	t->6	u->12	v->29	ä->4	å->4	ö->2	
 bör,	 ->1	
 bör.	F->1	
 börd	a->5	o->2	
 börj	a->104	
 börs	e->1	
 böte	r->1	
 c i 	E->1	
 c) l	i->1	
 ca 3	0->1	
 ca. 	1->1	
 calv	i->1	
 canc	e->2	
 cann	a->1	
 capi	t->10	
 case	.->1	
 ceme	n->2	
 cent	i->1	r->54	
 cert	i->5	
 chan	s->12	
 chap	e->1	
 char	a->1	t->1	
 chec	k->1	
 chef	 ->1	e->4	
 choc	k->4	
 chok	l->1	
 cirk	a->4	e->1	l->2	u->2	
 cita	t->1	
 cite	r->7	
 civi	l->19	
 comb	a->1	
 comm	o->1	
 comp	a->1	
 cond	i->1	
 cont	r->2	
 copy	r->1	
 corp	u->4	
 corr	e->1	
 cost	-->5	
 cric	k->1	
 d) i	 ->1	
 da C	o->5	
 da F	e->1	
 dag 	-->3	I->1	a->9	b->1	d->4	e->5	f->14	g->3	h->20	i->14	j->1	k->3	l->4	m->7	n->2	o->5	p->3	r->4	s->9	t->12	u->4	v->6	Ö->1	ä->16	
 dag,	 ->28	
 dag.	 ->1	(->1	A->1	D->7	E->1	F->2	G->1	H->3	I->2	J->6	K->1	O->1	V->1	
 dag:	 ->1	
 daga	r->17	
 dage	n->27	
 dagl	i->6	
 dago	r->52	
 dags	 ->14	l->2	t->2	
 dam 	s->1	
 dame	r->41	
 damm	 ->1	a->1	
 dans	k->24	
 data	 ->1	,->1	b->1	s->1	
 dato	 ->1	r->2	
 datu	m->13	
 de "	k->1	
 de 1	1->1	4->3	5->1	8->1	9->1	
 de 2	5->4	6->1	
 de 8	 ->1	
 de 9	 ->1	
 de C	e->2	
 de P	a->6	
 de a	d->2	f->1	k->5	l->21	m->3	n->33	r->9	t->5	v->8	
 de b	a->4	e->30	i->7	l->2	o->1	r->2	u->1	y->3	ä->5	å->6	ö->2	
 de c	e->3	h->1	
 de d	a->3	e->5	i->6	r->12	ä->3	
 de e	f->5	g->4	k->16	l->2	n->19	r->1	t->2	u->50	v->1	x->4	
 de f	a->22	e->7	i->6	j->3	l->24	o->8	r->36	u->2	y->7	å->7	ö->43	
 de g	a->10	e->9	j->1	o->4	r->26	ä->2	å->3	ö->1	
 de h	a->28	e->5	i->6	o->2	y->1	ä->11	å->3	ö->4	
 de i	 ->6	c->8	d->2	f->1	n->59	s->3	t->4	
 de j	o->1	u->3	
 de k	a->22	e->1	i->4	l->1	n->1	o->49	r->8	u->6	v->3	ä->1	
 de l	a->6	e->4	i->8	o->7	y->1	ä->11	å->4	ö->1	
 de m	a->4	e->35	i->18	o->1	u->3	y->9	ä->29	å->22	ö->2	
 de n	a->48	e->1	i->3	o->8	u->9	y->19	ä->11	ö->3	
 de o	b->3	c->5	f->9	l->45	m->19	p->1	r->8	v->2	
 de p	a->4	e->10	l->2	o->20	r->28	å->8	
 de r	a->3	e->34	i->12	u->1	ä->8	å->1	
 de s	a->4	e->35	i->3	j->4	k->28	l->2	m->21	n->1	o->48	p->2	t->53	u->2	v->8	y->5	ä->10	å->3	
 de t	a->6	e->3	i->17	j->1	o->3	r->12	u->3	v->19	y->3	
 de u	l->1	n->3	p->13	t->18	
 de v	a->9	e->18	i->26	ä->9	
 de y	r->2	t->11	
 de ä	l->1	m->1	n->10	r->18	v->1	
 de å	r->4	s->2	t->23	
 de ö	m->1	n->1	p->2	s->3	v->16	
 de, 	E->1	e->1	m->1	v->1	
 dead	l->1	
 deba	t->167	
 dece	m->19	n->22	
 defi	n->35	
 dege	n->1	
 degr	a->1	
 del 	-->1	a->70	b->1	d->1	f->1	h->3	i->11	k->3	l->1	m->5	o->2	p->5	s->3	t->1	v->1	ä->4	ö->1	
 del,	 ->4	
 del.	B->1	D->1	M->1	V->1	
 dela	 ->9	d->3	k->6	r->46	s->6	t->5	y->2	
 dele	g->20	n->30	
 delf	r->1	
 delg	i->1	
 dell	ö->1	
 deln	i->1	
 delr	a->1	
 dels	 ->13	t->4	
 delt	a->53	i->1	o->2	
 delu	t->2	
 delv	i->11	
 dem 	2->1	a->6	d->7	e->6	f->8	g->2	h->3	i->10	j->1	k->1	l->1	m->5	n->1	o->10	p->7	r->1	s->61	t->5	u->4	v->2	ä->1	
 dem,	 ->11	
 dem.	(->1	A->1	B->2	D->6	E->1	F->2	H->1	J->4	K->1	M->3	N->2	O->1	R->1	V->6	
 dem:	 ->2	
 dem?	D->1	
 dema	g->4	s->1	
 demo	g->3	k->106	n->13	
 den 	"->2	-->3	1->27	2->4	3->7	4->2	5->1	6->1	7->1	9->2	B->1	E->4	X->1	a->103	b->69	c->3	d->51	e->163	f->118	g->87	h->92	i->135	j->3	k->62	l->22	m->66	n->75	o->57	p->87	r->60	s->205	t->64	u->34	v->42	z->1	ä->25	å->11	ö->26	
 den)	,->1	
 den,	 ->10	
 den.	.->1	D->6	E->1	F->2	H->4	I->1	J->3	O->2	T->1	V->1	
 den;	 ->2	
 deni	e->2	
 denn	a->522	e->4	
 dens	a->4	
 depa	r->5	
 der 	E->1	L->7	
 dera	s->84	
 des 	f->1	
 desa	m->2	
 dess	 ->101	a->344	u->36	v->4	
 dest	o->2	r->1	
 det 	"->2	-->4	2->2	B->1	C->1	E->3	I->1	K->1	M->1	T->1	a->164	b->101	c->5	d->56	e->118	f->366	g->231	h->130	i->169	j->15	k->90	l->33	m->109	n->86	o->67	p->93	r->46	s->346	t->61	u->41	v->160	y->6	ä->321	å->11	ö->27	
 det!	.->2	
 det,	 ->44	
 det.	 ->2	(->1	A->4	D->8	E->6	H->8	I->3	J->5	K->1	M->7	O->1	P->1	S->1	V->13	
 det:	 ->2	
 det?	D->2	J->1	
 deta	l->34	
 dets	a->5	
 dett	a->828	
 dial	o->31	
 die 	a->1	
 diek	t->1	
 diff	e->5	
 dig 	f->1	s->1	
 dike	n->1	
 dikt	a->3	e->1	
 dile	m->3	
 dime	n->12	
 diox	i->2	
 dipl	o->11	
 dire	k->212	
 disc	i->14	
 disk	r->19	u->140	
 disp	e->1	o->3	
 dist	a->1	i->1	r->1	
 dit 	d->2	h->1	l->1	r->1	t->1	
 dith	ö->1	
 dive	r->4	
 djun	g->2	
 djup	 ->1	a->7	e->5	g->7	s->1	t->7	
 djur	 ->1	-->2	.->2	a->1	e->2	f->4	l->2	
 djär	v->7	
 djäv	u->2	
 dock	 ->59	,->2	
 dog 	i->1	
 dog.	D->1	S->1	
 dogm	 ->1	a->1	
 doku	m->39	
 doll	a->9	
 dom 	d->1	p->1	
 doma	r->16	
 dome	n->2	
 domi	n->7	
 doms	l->3	r->1	t->58	
 dra 	a->1	d->1	f->2	i->5	k->1	l->1	m->1	n->4	s->4	t->4	u->1	
 drab	b->45	
 drag	 ->3	,->1	.->1	a->1	i->2	n->1	
 dram	a->6	
 drar	 ->10	
 dras	 ->2	t->3	
 dric	k->3	
 drif	t->5	
 driv	a->13	e->4	k->3	
 drog	 ->1	b->1	e->1	k->1	s->2	
 drop	p->1	
 druc	k->2	
 drun	k->3	
 dryf	t->1	
 dryg	t->3	
 dråp	s->1	
 dröj	a->1	d->1	e->3	s->2	
 dröm	m->1	
 du b	a->1	e->1	
 du c	o->1	
 du m	i->1	
 du ä	r->2	
 dubb	e->6	l->9	
 duga	,->1	
 dukt	i->1	
 dumh	e->3	
 dump	a->1	n->3	
 dumt	 ->1	
 duna	n->1	
 duss	i->1	
 dvs.	 ->45	
 dyka	 ->2	
 dyke	r->5	
 dyli	k->3	
 dyna	m->5	
 dyr 	h->1	
 dyra	 ->2	r->2	
 dyrt	 ->1	.->1	
 dyst	r->1	
 däck	 ->1	
 dämp	a->2	
 där 	-->1	1->1	2->1	5->1	8->1	E->4	F->1	L->1	a->9	b->7	d->43	e->8	f->6	g->3	h->9	i->5	j->3	k->8	l->1	m->29	n->5	o->3	p->4	r->2	s->16	t->4	u->5	v->27	Ö->1	ä->4	å->1	
 där!	D->1	
 där,	 ->10	
 där.	 ->1	D->2	F->1	I->1	J->3	S->3	V->3	
 där?	J->1	
 dära	v->2	
 däre	f->7	m->13	
 därf	ö->184	
 därh	ä->1	
 däri	 ->1	b->6	f->2	g->15	
 därm	e->40	
 därp	å->2	
 därt	i->1	
 därv	i->4	
 då 2	4->1	
 då D	a->1	
 då E	G->1	r->1	u->1	
 då a	k->1	l->2	n->1	r->2	t->5	
 då b	a->1	e->5	l->1	ö->4	
 då d	e->16	
 då e	n->1	
 då f	a->1	i->1	o->1	r->3	å->1	ö->2	
 då g	e->2	
 då h	a->4	
 då i	 ->4	d->1	n->7	
 då j	a->2	u->1	
 då k	a->8	o->3	
 då m	a->2	e->3	y->1	å->2	ö->1	
 då o	c->6	l->1	m->2	
 då p	e->1	o->1	r->1	å->1	
 då r	i->1	ä->3	
 då s	e->1	j->1	k->5	n->1	o->2	ä->2	
 då t	a->2	i->3	r->1	y->1	ä->1	
 då u	n->1	
 då v	a->1	e->3	i->8	r->1	
 då ä	n->1	v->1	
 då ö	v->1	
 då, 	f->1	m->1	
 då.D	e->1	
 då?I	n->1	
 dåli	g->19	
 dåva	r->1	
 dö i	 ->1	
 död 	i->1	o->2	v->2	
 död.	A->1	J->1	M->1	
 döda	 ->1	,->1	d->3	n->1	s->2	t->1	
 dödf	ö->1	
 döds	d->1	f->1	
 döen	d->1	
 dölj	a->6	e->3	s->1	
 döma	 ->7	.->1	n->1	
 dömd	e->1	
 dömt	s->1	
 döpa	 ->1	
 döpe	r->2	
 döpt	e->1	
 dör 	e->1	f->1	m->1	u->1	
 dörr	 ->1	,->1	a->3	e->2	
 dött	.->2	r->1	
 e) i	 ->1	
 e-ma	i->1	
 e.d.	,->1	
 ecu 	m->1	
 ecu,	 ->1	
 ed g	e->1	
 eden	,->1	
 effe	k->129	
 efte	r->358	
 egen	 ->29	a->1	d->5	f->4	s->22	t->38	
 eget	 ->23	,->1	.->1	
 egna	 ->44	
 egoi	s->2	
 ej a	n->1	t->1	v->1	
 ej b	e->2	o->1	
 ej i	 ->1	
 ej k	o->1	
 ej l	ö->1	
 ej n	ä->1	
 ej ä	r->1	
 ej, 	m->1	
 ej.E	x->1	
 ej.R	å->1	
 ekol	o->13	
 ekon	 ->1	o->242	
 ekos	y->4	
 ekva	t->1	
 el- 	o->2	
 el-S	h->4	
 elef	a->1	
 elek	t->10	
 elem	e->9	
 elim	i->3	
 elle	r->323	
 elma	s->1	
 elog	e->2	
 elva	 ->2	
 emba	r->1	
 embl	e->1	
 embr	y->1	
 emed	a->1	
 emel	l->63	
 emig	r->2	
 emot	 ->50	.->4	i->1	
 en "	e->1	h->1	r->2	s->1	å->1	
 en P	R->1	
 en R	o->1	
 en S	c->1	
 en a	b->1	c->2	d->6	k->3	l->17	n->55	r->9	s->5	u->3	v->55	x->1	
 en b	a->6	e->38	i->10	l->2	o->5	r->24	u->4	y->2	ä->13	ö->3	
 en c	e->5	h->7	o->6	
 en d	a->5	e->68	i->18	j->5	o->4	r->2	u->1	y->1	ö->2	
 en e	f->17	g->7	k->17	l->8	n->33	r->2	u->55	v->2	x->11	
 en f	a->10	e->4	i->3	j->1	l->5	o->13	r->53	u->10	ä->1	ö->70	
 en g	a->14	e->45	i->3	l->1	n->2	o->8	r->24	u->1	å->48	
 en h	a->16	e->19	i->2	j->1	o->1	u->5	ä->6	å->13	ö->13	
 en i	 ->2	c->3	d->4	l->1	m->1	n->36	s->1	
 en j	a->2	u->2	ä->5	
 en k	a->14	e->1	l->10	o->76	r->14	u->8	v->5	ä->10	
 en l	a->5	e->4	i->15	o->2	u->1	y->1	ä->8	å->17	ö->13	
 en m	a->21	e->45	i->30	o->16	u->1	y->55	ä->13	å->3	ö->11	
 en n	a->8	e->6	i->2	o->3	y->30	ä->4	å->7	ö->8	
 en o	a->2	b->8	c->3	e->3	f->15	h->1	k->3	l->4	m->22	n->2	p->2	r->20	t->2	v->1	ä->1	ö->1	
 en p	a->9	e->11	l->3	o->40	r->14	u->8	y->1	å->1	
 en r	a->25	e->72	i->14	o->1	u->1	ä->16	å->2	é->1	ö->5	
 en s	a->29	c->2	e->7	i->14	j->6	k->15	l->6	m->4	n->7	o->20	p->8	t->110	u->4	v->2	y->8	ä->11	å->51	
 en t	a->3	e->7	i->32	j->4	o->4	r->10	u->5	v->1	y->15	
 en u	n->15	p->16	r->2	t->32	
 en v	a->6	e->13	i->66	ä->23	å->2	
 en y	t->3	
 en z	i->1	
 en ä	n->13	
 en å	k->2	l->1	s->2	t->11	
 en ö	d->1	k->19	m->1	n->1	p->3	r->1	s->2	v->27	
 en, 	N->1	s->1	
 en.E	f->1	
 ena 	e->5	f->1	g->4	h->1	i->1	l->1	m->1	o->1	p->1	r->1	s->14	y->1	ä->2	ö->1	
 enad	e->5	
 enas	 ->5	t->2	
 enat	.->1	s->1	
 enba	r->30	
 end 	o->1	
 enda	 ->48	.->1	s->71	
 ende	m->1	
 ener	g->98	
 enga	g->18	
 enge	l->10	
 enhe	t->53	
 enhä	l->32	
 enig	 ->1	a->4	h->5	
 enke	l->36	
 enkl	a->11	
 enli	g->122	
 enor	m->32	
 ens 	a->1	d->3	h->1	k->1	l->1	m->2	n->1	p->2	v->2	
 ensa	m->7	
 ense	 ->2	,->1	
 ensi	d->4	
 ensk	i->28	
 enst	a->5	
 entr	e->4	
 entu	s->3	
 enty	d->4	
 enve	t->1	
 envi	s->5	
 epok	 ->1	,->1	e->2	
 er -	 ->2	
 er a	l->1	n->2	t->22	
 er b	e->3	i->1	
 er d	e->3	
 er e	g->1	n->4	t->5	
 er f	r->3	ö->4	
 er g	r->1	
 er h	a->1	u->1	ä->1	
 er i	 ->1	g->1	n->2	
 er k	o->4	u->1	ä->1	
 er l	e->1	
 er m	e->1	y->1	
 er n	ä->1	
 er o	c->2	m->13	r->5	
 er p	o->1	r->1	å->2	
 er r	e->1	ö->1	
 er s	a->1	i->1	j->2	o->6	t->2	y->2	
 er t	a->3	i->5	o->1	
 er u	p->9	r->1	t->1	
 er v	a->2	i->3	
 er ä	r->1	
 er å	t->1	
 er, 	M->1	a->1	e->1	f->5	h->3	i->1	k->2	l->2	m->1	o->2	p->1	s->2	u->1	v->1	ä->1	
 er.B	e->1	
 er.J	a->3	
 er.K	o->1	
 er.N	ä->1	
 er.O	c->1	
 er.P	r->1	
 er: 	K->1	d->1	
 era 	d->1	e->3	f->5	i->2	k->3	l->1	m->1	o->2	p->4	r->6	t->7	u->1	ä->1	
 erbj	u->18	ö->1	
 erfa	r->26	
 erfo	r->5	
 erhå	l->7	
 erhö	l->3	
 erin	r->13	
 erkä	n->39	
 ersa	t->1	
 ersä	t->21	
 ert 	b->8	d->1	e->1	f->5	i->2	o->2	p->3	s->5	u->5	y->1	ä->3	
 ert,	 ->2	
 eröv	r->1	
 et o	r->1	
 etab	l->12	
 etap	p->4	
 etc.	 ->3	D->1	E->1	
 etc?	A->1	
 etik	 ->1	
 etis	k->1	
 etni	s->11	
 ett 	"->1	5->1	A->1	E->15	a->113	b->86	c->4	d->42	e->68	f->121	g->39	h->31	i->48	j->8	k->46	l->39	m->105	n->31	o->63	p->84	r->39	s->196	t->45	u->37	v->42	w->1	y->5	ä->14	å->23	ö->15	
 ett,	 ->2	
 ett.	.->1	F->1	
 ett:	 ->1	
 euro	 ->16	!->1	,->6	.->8	f->1	n->6	o->1	p->350	s->2	
 even	e->1	t->20	
 evig	 ->1	t->2	
 ex a	n->4	
 ex p	o->1	
 ex t	u->1	
 exak	t->18	
 exam	e->6	i->10	
 exce	p->5	
 exem	p->116	
 exil	r->1	t->1	
 exis	t->17	
 exkl	u->3	
 expa	n->6	
 expe	d->1	r->44	
 expl	i->1	o->1	
 expo	n->2	r->3	
 exte	r->7	
 extr	a->6	e->24	
 f.d.	 ->2	
 fabr	i->1	
 fack	f->4	
 fadd	e->1	
 fail	u->1	
 fakt	a->9	i->49	o->11	u->64	
 fall	 ->78	,->7	.->10	e->61	i->3	s->1	
 fals	k->3	
 fami	l->15	
 fann	 ->2	s->13	
 fant	a->11	
 far 	a->1	
 fara	 ->6	,->2	n->2	
 farh	å->2	
 farl	i->58	
 farm	a->1	
 faro	r->4	
 fars	o->1	
 fart	 ->1	y->60	
 farv	a->9	
 fas,	 ->1	
 fasc	i->7	
 faso	r->1	
 fast	 ->24	.->2	a->5	k->1	l->5	n->1	s->72	ä->1	
 fatt	a->49	i->30	
 faun	a->1	
 favo	r->1	
 faxa	 ->1	
 febr	u->16	
 fede	r->8	
 fel 	a->4	o->2	s->3	u->1	
 fel!	 ->1	
 fel,	 ->3	
 fel.	D->2	G->1	J->1	
 fela	k->12	n->1	
 felb	e->1	
 felk	v->1	
 felr	ä->1	
 fels	y->1	
 fem 	a->3	d->1	g->1	k->2	m->1	p->2	v->2	å->13	
 fem,	 ->1	
 fem:	 ->1	
 femp	u->1	
 femt	e->16	i->3	o->5	
 femå	r->3	
 feno	m->3	
 fick	 ->26	
 fien	d->1	t->2	
 film	e->1	
 filo	s->5	
 fin 	s->1	
 fina	 ->2	n->75	
 finl	ä->5	
 finn	a->56	e->10	s->315	
 fins	k->6	
 fira	 ->1	
 fisk	 ->1	a->6	b->4	e->29	
 fjol	 ->2	.->1	
 fjor	t->9	
 fjär	d->11	
 flag	g->12	r->1	
 flam	s->4	
 fler	 ->23	,->1	a->56	s->1	t->5	å->12	
 fles	t->25	
 flex	i->27	
 flic	k->1	
 flit	 ->1	e->1	
 flod	 ->2	e->2	
 flor	a->1	
 flot	t->2	
 flyg	,->1	a->2	b->1	e->2	k->1	p->4	t->2	
 flyk	t->14	
 flyr	 ->1	
 flyt	a->1	t->9	
 fläk	t->1	
 flöd	e->1	
 fode	r->6	
 fog 	f->1	
 foga	d->1	
 foku	s->5	
 folk	 ->11	,->1	.->8	e->20	g->2	h->9	o->6	p->10	r->3	s->5	v->2	
 fond	 ->6	e->16	m->3	u->1	
 fora	 ->1	
 forc	e->1	
 ford	o->60	r->8	
 form	 ->21	,->1	.->2	a->2	e->30	u->14	
 fors	k->36	
 fort	 ->3	b->1	f->89	g->5	l->1	s->93	
 foru	m->3	
 forê	t->1	
 foss	i->2	
 fotb	o->1	
 fotf	ä->1	
 fots	p->2	
 frak	t->1	
 fram	 ->205	,->8	.->7	f->143	g->50	h->24	k->11	l->20	m->1	s->48	t->114	å->21	ö->2	
 fran	c->1	s->35	
 fras	e->1	
 fred	 ->15	,->1	.->3	e->1	l->8	s->36	
 frek	v->1	
 fres	t->4	
 fri 	f->1	k->2	r->8	ö->1	
 fri,	 ->1	
 fri-	 ->8	
 fria	 ->21	,->2	t->1	
 frig	j->1	ö->5	
 frih	a->2	e->64	
 frik	t->1	
 fris	l->2	t->3	
 frit	t->3	
 friv	i->12	
 frod	a->4	
 fron	t->2	
 fru 	A->2	F->1	P->1	R->3	S->3	T->1	W->1	k->42	t->13	
 fru,	 ->1	
 fruk	t->16	
 frus	t->2	
 frys	a->2	
 fräc	k->1	
 främ	j->56	l->34	m->2	s->47	
 fråg	a->460	e->11	o->204	
 från	 ->565	,->1	g->1	t->3	v->8	
 full	 ->8	a->6	b->3	f->3	g->2	k->5	o->5	s->39	t->21	v->2	ä->2	
 fult	 ->1	
 fund	a->1	e->12	
 fung	e->54	
 funk	t->27	
 funn	i->9	
 fusi	o->7	
 fusk	.->1	
 futt	i->1	
 fyll	a->4	s->1	t->2	
 fyra	 ->23	,->1	:->1	
 fyrt	i->3	
 fysi	s->9	
 fäde	r->1	
 fäll	d->1	e->1	t->2	
 fält	 ->1	e->5	
 fäng	e->1	
 färd	 ->1	i->4	
 färg	,->1	
 färr	e->2	
 färs	k->1	
 fäst	 ->1	a->3	e->6	n->1	s->1	
 få 1	0->1	
 få E	u->1	
 få G	o->1	
 få a	l->1	n->1	r->1	v->2	
 få b	e->3	o->2	ä->2	ö->1	
 få d	e->14	i->1	o->1	
 få e	f->2	n->27	r->1	t->11	
 få f	a->1	i->1	l->1	o->1	r->4	u->1	ö->4	
 få g	a->1	e->1	
 få h	i->1	j->1	
 få i	 ->3	g->1	n->3	
 få k	o->4	v->2	
 få l	a->1	i->1	o->2	ä->3	
 få m	a->2	e->2	y->1	å->3	ö->1	
 få n	å->3	
 få o	b->1	m->1	r->2	s->2	
 få p	a->1	e->2	o->2	r->2	u->1	å->1	
 få r	e->3	y->1	ä->1	
 få s	a->2	e->6	i->2	l->1	t->9	ä->2	å->3	
 få t	a->6	i->16	
 få u	p->1	t->2	
 få v	a->1	e->6	i->3	å->1	
 få ä	r->1	
 få å	t->1	
 få ö	k->1	
 få, 	o->2	r->1	
 få.E	u->1	
 få.G	r->1	
 få.V	i->1	
 fåge	l->3	
 fågl	a->6	
 fång	a->2	s->3	
 får 	M->1	O->1	a->7	b->3	d->14	e->19	f->6	g->5	h->3	i->39	j->2	k->5	l->2	m->10	n->4	o->5	p->2	r->1	s->15	t->11	u->2	v->21	y->1	ä->2	å->1	
 får,	 ->2	
 får?	N->1	
 fårk	ö->1	
 fås 	f->1	
 fåta	l->1	
 fått	 ->56	.->1	
 född	e->1	
 föde	l->2	r->2	
 födo	ä->1	
 föds	 ->1	
 föga	 ->2	
 följ	a->63	d->39	e->12	s->4	t->3	
 föll	 ->3	.->1	
 föns	t->1	
 för 	"->4	-->2	1->15	2->5	3->1	5->2	7->1	A->4	B->4	C->1	D->2	E->62	F->5	G->2	H->1	I->4	K->3	L->2	O->1	P->3	S->2	T->8	V->1	W->1	a->804	b->59	c->7	d->501	e->211	f->103	g->35	h->69	i->37	j->22	k->128	l->52	m->126	n->73	o->69	p->64	r->95	s->163	t->76	u->86	v->89	y->2	Ö->1	ä->6	å->32	ö->44	
 för,	 ->16	
 för.	 ->1	(->1	D->2	H->1	J->1	M->3	V->4	
 för;	 ->1	
 för?	F->1	I->1	
 föra	 ->19	n->7	r->2	s->7	
 förb	a->3	e->31	i->32	j->14	l->15	r->4	u->28	ä->77	
 förd	a->3	e->32	j->11	o->2	r->110	u->3	ä->4	ö->20	
 före	 ->26	b->23	d->155	f->21	g->19	h->1	k->22	l->27	m->13	n->24	s->160	t->242	
 förf	a->53	i->1	j->1	l->18	o->18	r->5	ä->3	å->1	ö->4	
 förg	l->2	r->3	ä->1	
 förh	a->79	i->30	o->9	å->45	ö->1	
 föri	n->3	r->1	
 förk	a->8	l->60	n->3	o->2	r->1	u->2	
 förl	a->3	e->2	i->53	o->20	u->6	ä->6	å->2	
 förm	e->5	i->3	o->11	y->1	å->33	ö->1	
 förn	a->1	e->10	u->14	y->49	
 föro	l->2	r->67	
 förp	a->5	l->21	
 förr	 ->3	,->1	a->42	e->4	g->3	i->1	ä->5	
 förs	 ->6	a->10	e->31	i->63	k->8	l->257	o->5	t->381	u->9	v->81	ä->48	å->1	ö->60	
 fört	 ->6	e->1	i->6	j->19	r->59	s->2	v->1	y->3	ä->1	
 föru	n->1	t->75	
 förv	a->51	e->22	i->19	r->1	ä->51	å->6	
 förä	n->67	
 förå	l->3	
 förö	d->5	v->3	
 fött	e->3	
 gagn	 ->3	a->4	
 gale	n->1	
 gall	r->1	
 galn	a->1	
 gaml	a->28	
 gamm	a->4	
 gans	k->26	
 gara	n->90	
 gard	e->1	
 gask	a->1	
 gato	r->1	
 gav 	e->1	h->2	m->2	n->1	p->1	u->1	v->1	
 gav,	 ->1	
 gavs	 ->2	
 ge F	r->1	
 ge a	k->2	l->2	n->2	r->2	
 ge b	e->1	i->3	ä->1	å->1	
 ge d	e->13	
 ge e	n->9	r->6	t->12	
 ge f	e->1	ö->2	
 ge g	a->1	r->1	
 ge h	a->1	j->2	ö->1	
 ge i	n->3	
 ge j	o->1	
 ge k	l->2	o->2	
 ge m	a->1	e->1	i->2	
 ge n	ä->1	å->1	
 ge o	c->1	f->1	s->8	
 ge p	a->3	e->1	o->1	r->1	
 ge r	a->1	e->2	i->1	o->1	ä->1	å->3	
 ge s	i->4	t->2	å->1	
 ge t	i->2	y->1	
 ge u	n->1	p->2	t->9	
 ge v	a->1	i->1	ä->1	
 ge.J	a->1	
 gedi	g->2	
 geme	n->379	
 gena	n->1	s->10	
 gend	e->6	
 gene	r->37	t->1	
 geng	ä->1	
 geno	m->378	
 gens	v->1	
 gent	e->27	
 genu	s->1	
 geog	r->8	
 geos	t->2	
 ger 	E->1	b->1	d->4	e->5	f->3	g->2	i->6	k->3	m->8	n->2	o->5	p->1	r->2	s->7	t->2	u->10	v->1	
 ger,	 ->1	
 ges 	d->2	e->1	f->1	i->1	k->1	n->2	s->1	t->2	u->1	y->1	ö->1	
 gest	 ->1	?->1	
 gett	 ->21	
 gick	 ->8	
 gift	i->2	
 giga	n->5	
 gill	a->1	
 gilt	i->15	
 giss	l->1	
 giva	n->3	r->14	
 give	n->1	s->1	t->25	
 givi	t->4	
 gjor	d->29	t->83	
 glad	 ->19	a->3	d->2	
 glas	.->1	h->1	
 gles	a->1	
 glob	a->12	
 glup	s->1	
 gläd	e->19	j->15	s->6	
 glöm	m->14	s->1	t->4	
 gnut	t->2	
 gnäl	l->1	
 god 	a->2	b->1	f->6	i->3	j->1	l->1	m->1	t->6	u->1	v->1	
 god.	F->1	
 goda	 ->36	.->1	
 godk	ä->88	
 godo	.->3	
 gods	 ->29	,->1	.->4	;->1	N->1	e->2	
 godt	a->38	o->2	y->6	
 golv	e->1	
 gott	 ->17	.->1	g->1	
 grad	 ->12	.->2	e->6	v->3	
 gran	d->3	n->5	s->55	
 grat	i->4	u->36	
 grav	e->4	t->1	
 grek	e->1	i->6	
 grep	p->2	
 grip	a->4	e->2	i->2	
 grog	r->1	
 grou	p->1	
 grov	 ->1	
 grun	d->255	
 grup	p->138	
 gruv	a->1	
 grym	t->1	
 gräl	 ->2	
 gräm	e->1	
 grän	s->57	
 grå 	v->1	
 gråz	o->1	
 gröd	o->1	
 grön	 ->2	a->13	b->1	t->1	
 gröv	s->1	
 guds	 ->2	
 guld	e->1	
 gult	 ->1	
 gumm	i->1	
 guve	r->1	
 gynn	a->9	s->2	
 gäck	 ->1	
 gäll	a->29	d->11	e->362	t->2	
 gärn	a->32	i->1	
 gå a	n->1	t->1	
 gå b	e->2	
 gå e	t->1	
 gå f	r->4	ö->3	
 gå g	r->2	
 gå h	e->1	
 gå i	 ->1	g->4	n->15	
 gå l	ä->4	å->1	
 gå m	e->3	
 gå o	c->2	f->1	
 gå p	å->1	
 gå s	a->1	n->1	o->1	å->1	
 gå t	i->10	
 gå u	n->1	t->4	
 gå v	i->4	
 gå å	t->1	
 gå.O	m->1	
 gå.V	i->1	
 gång	 ->66	,->3	.->7	e->51	n->2	s->3	
 går 	a->6	b->2	d->7	f->5	g->2	h->2	i->13	k->1	l->2	m->6	o->2	p->2	s->3	t->12	u->12	v->3	å->2	ö->1	
 går,	 ->4	
 går.	J->1	V->1	
 gård	a->3	
 gått	 ->18	.->2	
 gömm	a->1	e->2	
 gömt	s->1	
 gör 	E->1	a->28	d->49	e->4	f->1	g->2	h->3	i->3	m->9	n->5	o->4	p->3	s->4	t->2	u->2	v->7	ä->4	
 gör,	 ->1	
 gör.	D->2	E->1	
 göra	 ->234	,->7	.->13	?->1	s->29	
 görs	 ->9	,->4	.->2	
 ha a	n->3	r->1	t->1	
 ha b	e->4	r->1	
 ha d	e->7	i->1	r->1	ö->1	
 ha e	g->1	n->36	r->1	t->17	
 ha f	r->3	u->1	ö->2	
 ha g	e->2	j->2	r->1	
 ha h	a->2	i->1	ö->4	
 ha i	 ->1	n->2	
 ha k	l->1	o->5	u->2	v->1	ä->1	
 ha l	y->3	ä->1	
 ha m	a->2	e->2	i->1	o->2	y->2	ö->3	
 ha n	e->1	y->1	å->8	
 ha o	c->1	f->1	
 ha p	r->2	
 ha r	ä->2	å->1	
 ha s	a->4	e->1	j->1	k->3	t->3	u->1	y->1	
 ha t	a->1	i->4	r->1	v->3	y->2	
 ha u	n->2	p->1	t->2	
 ha v	a->7	e->1	i->3	ä->3	
 ha y	t->1	
 ha ä	g->1	n->1	
 ha å	s->1	
 ha ö	n->2	v->1	
 ha, 	e->1	
 ha.A	l->1	
 hade	 ->84	?->1	
 haft	 ->34	,->2	.->1	
 haka	t->1	
 halt	 ->1	
 halv	 ->3	a->4	h->1	m->1	t->5	v->2	å->5	ö->3	
 hamb	u->1	
 hamm	a->1	
 hamn	 ->3	.->1	a->28	b->1	e->2	i->1	k->2	
 han 	a->6	b->3	d->2	e->1	f->5	g->3	h->22	i->14	j->2	k->7	l->5	m->2	n->3	o->3	p->3	s->12	t->5	u->3	v->6	ä->9	ö->1	
 han,	 ->2	
 hand	 ->39	,->3	.->2	?->1	e->21	f->1	i->4	l->177	s->8	u->2	
 hank	a->1	
 hans	 ->76	
 hant	e->32	v->2	
 happ	y->1	
 har 	-->2	1->2	4->1	A->1	B->1	E->7	G->1	L->2	P->1	S->1	a->85	b->78	c->1	d->97	e->96	f->171	g->92	h->61	i->102	j->39	k->55	l->91	m->67	n->63	o->30	p->37	r->53	s->131	t->72	u->54	v->139	ä->21	å->4	ö->12	
 har,	 ->14	
 har.	D->1	T->1	
 har:	 ->1	
 har?	N->1	
 harm	o->18	
 hast	i->1	
 hat 	o->1	
 hate	t->1	
 hati	s->1	
 hatt	e->1	
 hav 	f->1	o->1	
 hav,	 ->1	
 have	n->2	r->6	t->15	
 havs	 ->4	,->4	.->4	?->1	f->2	m->2	v->1	
 hebr	e->1	
 hede	r->3	
 hedr	a->3	
 hejd	a->2	
 hekt	a->2	
 hel 	b->1	d->6	k->1	p->1	r->2	
 hela	 ->105	
 helg	e->1	
 helh	e->21	j->8	
 heli	g->1	
 hell	e->47	r->5	
 hels	i->1	t->46	
 helt	 ->135	,->1	.->3	ä->4	
 hem 	e->1	f->1	o->2	t->1	
 hem.	 ->1	N->1	
 hemb	y->1	
 hemf	ö->1	
 heml	a->3	i->5	ä->2	ö->5	
 hemm	a->9	e->1	
 hems	k->3	
 hemv	i->1	
 henn	e->27	
 herr	 ->165	a->44	
 hes 	i->1	
 heta	 ->1	
 hete	r->2	
 hets	 ->1	e->1	
 hett	 ->1	a->1	e->1	
 hier	a->4	
 high	 ->1	
 hind	e->23	r->20	
 hinn	a->2	
 hist	o->33	
 hit 	m->2	o->1	s->1	
 hit,	 ->1	
 hitt	a->17	i->41	
 hjäl	p->99	
 hjär	t->18	
 hobb	y->2	
 hoc-	d->1	t->1	
 homo	f->1	g->2	s->1	
 hon 	a->1	f->4	h->4	i->4	j->1	k->2	l->1	p->2	s->4	t->2	u->1	v->1	ä->2	
 hono	m->28	
 hopp	 ->1	a->97	e->1	l->1	
 hord	 ->1	e->1	
 hori	s->3	
 horm	o->1	
 hos 	D->1	E->2	F->1	R->1	a->3	b->2	d->12	e->2	f->3	k->6	m->4	o->4	p->2	r->1	s->2	t->1	v->2	
 hosp	i->1	
 hot 	-->1	f->1	m->6	o->1	p->1	s->1	
 hota	 ->1	d->5	n->1	r->6	s->4	t->1	
 hotb	i->1	
 hote	l->1	t->7	
 hotf	u->1	
 hugg	 ->3	
 huma	n->6	
 huml	e->1	
 humö	r->2	
 hund	.->1	r->10	
 hur 	E->2	a->5	b->7	d->42	e->3	f->5	g->2	h->4	i->1	k->11	l->9	m->24	n->5	o->2	p->6	r->1	s->26	t->3	u->7	v->31	
 hur.	K->1	R->1	
 huru	v->14	
 hus 	h->1	o->1	s->1	
 hus,	 ->2	
 hus.	H->1	
 husö	v->1	
 huvu	d->47	
 hyck	l->5	
 hygi	e->2	
 hyll	a->1	n->1	
 hypo	t->2	
 hyrd	 ->1	
 hysa	 ->3	
 hyse	r->5	
 hyst	e->1	
 häft	i->1	
 häle	r->1	
 hälf	t->3	
 häls	a->15	n->1	o->7	
 hämm	a->1	
 hämn	a->1	i->1	
 händ	a->12	e->60	
 hänf	ö->1	
 häng	a->1	b->1	e->12	
 häns	e->8	y->71	
 hänt	 ->5	.->1	:->1	
 hänv	i->35	
 här 	-->6	D->1	a->6	b->9	c->1	d->9	e->3	f->41	g->4	h->6	i->59	k->8	l->5	m->3	n->2	o->14	p->16	r->5	s->18	t->15	u->5	v->11	y->2	ä->8	å->2	ö->2	
 här,	 ->14	
 här.	 ->1	D->3	E->1	F->1	K->1	V->2	
 här;	 ->1	
 här?	D->1	
 häre	f->1	
 häri	g->2	
 härj	a->2	
 härl	e->1	
 härm	e->3	
 härr	ö->4	
 härt	i->1	
 härv	i->1	
 häst	e->1	
 häva	 ->1	
 hävd	a->27	v->1	
 hävt	s->1	
 hål 	i->1	
 hål,	 ->1	
 håll	 ->8	,->3	.->1	:->1	a->34	b->25	e->53	i->8	n->11	s->3	
 hån 	m->1	
 håna	r->1	
 hård	 ->3	,->1	a->11	n->2	
 håre	t->1	
 hårk	l->1	
 hårt	 ->7	,->1	.->1	
 håva	r->1	
 hög 	a->1	b->1	f->1	g->6	i->1	k->1	n->2	p->2	s->6	
 hög,	 ->1	
 höga	 ->13	,->1	.->1	k->1	
 höge	 ->2	r->16	
 högl	j->1	
 högn	i->3	
 högr	a->1	e->19	
 högs	k->1	t->28	
 högt	 ->9	,->1	.->1	e->2	i->4	
 höja	 ->4	s->1	
 höjd	 ->5	e->1	p->2	
 höje	r->1	
 höjn	i->2	
 höjt	s->1	
 höll	 ->4	s->2	
 höna	 ->1	
 hör 	a->4	b->1	d->1	e->1	f->1	h->6	i->3	j->1	n->2	s->2	t->7	v->2	
 hör.	 ->1	
 höra	 ->19	,->1	s->2	
 hörd	.->1	e->4	
 hörn	 ->2	s->1	
 hört	 ->15	,->1	s->1	
 höst	 ->1	
 i "g	e->1	
 i - 	a->1	
 i 15	 ->1	
 i 20	 ->1	0->2	
 i AB	B->1	
 i Ad	a->1	r->1	
 i Af	r->3	
 i Ak	k->2	
 i Al	s->1	
 i Am	s->17	
 i As	i->1	
 i Au	v->1	
 i Av	i->1	
 i BN	I->1	
 i Be	l->2	r->9	
 i Bi	s->5	
 i Bo	r->1	
 i Br	a->2	e->2	y->7	
 i Bu	d->1	
 i CE	N->1	
 i Ca	v->1	
 i Ce	n->5	r->1	
 i Cu	s->1	
 i DD	R->1	
 i Da	n->9	
 i Du	b->4	
 i EC	H->1	
 i EG	-->8	
 i EK	S->3	
 i EM	U->1	
 i EU	 ->2	,->1	-->5	:->7	
 i Ek	o->1	
 i Et	i->1	
 i Eu	r->171	
 i Fa	c->1	
 i Fe	i->1	
 i Fi	n->2	
 i Fo	l->1	
 i Fr	a->11	
 i Fö	r->14	
 i GU	E->1	
 i Ga	z->2	
 i Ge	n->2	
 i Go	l->2	
 i Gr	e->2	u->2	
 i Gu	a->1	l->1	
 i Ha	i->1	
 i He	l->14	
 i IC	E->2	
 i In	d->1	
 i Ir	l->10	
 i Is	r->1	t->1	
 i It	a->6	
 i Jo	n->1	
 i Ka	r->1	u->2	
 i Kf	o->1	
 i Ki	n->3	
 i Ko	s->34	u->1	
 i Ky	o->1	
 i Kä	r->1	
 i Kö	l->1	
 i La	n->1	p->2	
 i Le	a->1	
 i Li	l->1	s->5	
 i Lo	m->1	n->4	r->1	
 i Lu	t->1	x->4	
 i Ma	a->2	c->1	d->2	
 i Mc	N->1	
 i Me	d->1	l->14	x->1	
 i Mi	t->1	
 i Mo	n->2	s->1	
 i Ne	d->4	w->1	
 i No	r->1	
 i OL	A->1	
 i Om	a->1	
 i PP	E->3	
 i Pa	d->1	r->1	y->1	
 i Pe	k->1	
 i Po	r->5	
 i Ra	p->1	
 i Ro	m->1	
 i Ry	s->2	
 i Sa	i->1	n->2	
 i Sc	h->4	
 i Se	a->3	
 i Sh	a->1	e->3	
 i Sk	o->2	
 i Sr	i->3	
 i St	o->11	r->4	
 i Sv	e->2	
 i Sy	d->2	r->2	
 i TV	-->1	
 i Ta	d->2	m->14	u->1	
 i Te	x->1	
 i Th	e->4	y->1	
 i Ti	b->5	
 i Tu	r->7	
 i Ty	s->5	
 i UE	N->1	
 i US	A->3	
 i Ur	b->1	
 i Va	n->1	
 i Ve	n->1	
 i Vä	r->1	
 i Wa	l->3	s->1	
 i Wi	e->1	
 i Ya	s->1	
 i ab	s->1	
 i ai	d->1	
 i ak	t->4	
 i al	l->52	
 i an	a->1	d->15	n->4	p->1	s->7	v->1	
 i ar	b->21	t->15	
 i at	t->12	
 i av	s->3	t->2	v->2	
 i ba	l->1	
 i be	g->1	h->5	r->3	s->12	t->15	
 i bi	l->12	o->2	
 i br	i->1	o->1	u->1	ä->1	
 i bu	d->9	
 i bå	d->3	
 i bö	c->1	r->5	
 i ce	n->2	
 i ci	r->1	
 i da	g->165	n->1	t->1	
 i de	 ->80	b->10	c->7	m->3	n->200	r->1	s->25	t->197	
 i di	a->2	r->14	s->3	
 i do	k->1	m->2	
 i dr	i->1	
 i ef	t->8	
 i eg	e->12	
 i ek	o->5	
 i en	 ->98	k->1	l->27	s->1	
 i er	 ->3	a->4	t->7	
 i et	t->61	
 i eu	r->3	
 i ex	a->1	p->1	
 i f.	d->1	
 i fa	l->3	r->2	t->2	
 i fe	b->7	m->3	
 i fi	n->1	
 i fj	o->2	
 i fl	e->5	
 i fo	l->4	r->27	
 i fr	a->56	e->8	i->1	o->1	ä->1	å->74	
 i fu	l->2	n->1	
 i fy	r->2	
 i fä	r->2	
 i fö	l->2	r->139	
 i ga	r->1	
 i ge	m->14	n->9	
 i gl	a->1	
 i go	d->7	t->1	
 i gr	u->8	
 i gä	l->1	
 i gå	n->6	r->17	
 i ha	m->6	n->13	r->1	v->7	
 i he	l->21	m->1	n->1	
 i hi	e->1	s->1	
 i hj	ä->2	
 i hu	v->7	
 i hä	n->9	
 i hå	r->1	
 i hö	g->8	s->1	
 i ic	k->2	
 i in	d->1	f->2	i->1	k->2	l->2	s->2	
 i it	a->1	
 i ja	n->1	
 i jo	r->1	
 i ju	l->5	n->6	
 i jä	m->3	
 i ka	b->1	l->1	m->21	n->1	p->3	t->1	
 i ke	d->1	
 i kl	a->3	
 i kn	i->1	
 i ko	a->1	m->27	n->17	
 i kr	a->24	i->2	
 i ku	l->2	r->2	
 i kv	ä->4	
 i la	g->10	n->6	
 i le	d->2	
 i li	k->9	n->5	v->1	
 i lj	u->5	
 i ly	s->1	
 i lä	n->1	
 i lå	t->1	
 i ma	j->5	k->1	n->2	r->3	s->1	
 i me	d->33	l->1	r->1	
 i mi	g->1	l->6	n->20	t->18	
 i mj	u->1	
 i mo	r->32	t->9	
 i my	c->2	
 i mä	n->1	
 i må	l->6	n->15	
 i mö	b->1	
 i na	t->3	
 i ni	v->4	
 i no	r->2	v->5	
 i nu	l->1	
 i ny	a->1	h->1	
 i nä	r->7	s->1	
 i nå	g->10	
 i nö	d->1	
 i oc	h->16	
 i of	f->3	ö->1	
 i ok	t->2	
 i ol	i->4	j->1	y->1	
 i om	f->1	r->17	
 i on	s->1	
 i or	d->7	o->1	
 i ou	n->1	
 i oö	v->1	
 i pa	r->38	
 i pe	n->1	r->3	
 i pl	a->3	e->4	å->1	
 i po	l->6	r->2	s->2	
 i pr	a->10	e->4	i->12	o->14	
 i pu	n->2	
 i ra	d->1	m->1	p->8	
 i re	a->5	f->2	g->21	l->2	s->6	t->1	
 i ri	k->4	n->1	
 i ru	l->1	
 i rä	t->11	
 i rå	d->34	
 i sa	k->1	m->54	
 i se	n->1	p->12	x->1	
 i si	d->1	g->19	k->2	n->56	s->2	t->24	
 i sj	u->1	ä->23	
 i sk	a->2	e->1	o->2	u->1	y->2	
 i sl	u->19	
 i sm	å->2	
 i sn	a->2	
 i so	c->2	m->1	r->1	
 i sp	ä->1	
 i st	a->5	i->2	o->11	r->13	y->1	ä->47	å->4	ö->12	
 i sv	a->1	
 i sy	d->1	f->8	n->45	s->4	
 i sä	k->2	m->1	n->1	
 i så	 ->5	d->6	v->1	
 i sö	d->1	
 i t.	e->1	
 i ta	k->3	l->2	n->2	
 i te	x->1	
 i ti	d->12	l->9	
 i tj	ä->1	
 i to	l->1	p->3	r->1	
 i tr	a->4	e->4	ä->1	å->1	
 i tv	e->1	å->5	
 i tä	t->2	
 i un	d->3	g->1	i->31	
 i up	p->4	
 i ur	s->1	v->1	
 i ut	b->2	f->3	k->1	l->2	n->1	o->1	s->24	t->1	v->5	ö->1	
 i va	c->1	d->2	l->1	n->6	r->17	
 i ve	c->1	r->8	t->1	
 i vi	k->1	l->18	n->1	s->23	t->13	
 i vä	g->3	l->1	n->3	r->12	s->1	
 i vå	r->60	
 i yr	k->2	
 i yt	t->2	
 i zo	n->2	
 i ÖV	P->1	
 i Ös	t->37	
 i äg	a->1	
 i äk	t->1	
 i äm	n->2	
 i än	d->8	n->1	
 i är	e->1	
 i år	 ->3	,->3	.->4	a->1	t->1	
 i åt	a->1	e->3	g->1	
 i ör	e->1	
 i ös	t->3	
 i öv	e->12	r->5	
 i, s	å->1	
 i, u	t->1	
 i.An	l->1	
 i.De	t->2	
 i.Nä	r->1	
 i.Se	d->1	
 i.Så	 ->1	
 iakt	t->8	
 ians	p->1	
 iber	i->1	
 ibla	n->19	
 icke	 ->15	-->19	
 idag	,->1	
 idea	l->5	
 idee	l->2	
 iden	t->18	
 ideo	l->5	
 idro	t->4	
 idé 	-->1	a->2	j->1	k->1	o->1	s->3	ä->1	
 idé,	 ->1	
 idée	r->8	
 idén	 ->13	,->1	
 ifal	l->2	
 ifrå	g->21	n->14	
 igen	 ->10	"->1	,->7	.->9	:->1	o->18	
 igno	r->4	
 igån	g->7	
 ihjä	l->1	
 ihop	 ->8	.->2	
 ihär	d->1	
 ihåg	 ->15	.->1	
 ikap	p->1	
 ikra	f->4	
 illa	 ->3	,->2	v->1	
 ille	g->8	
 illo	j->2	
 illv	i->1	
 ilsk	a->2	
 imag	e->1	i->1	
 imma	t->1	
 immi	g->6	
 immu	n->1	
 impl	e->1	
 impo	n->3	p->1	r->5	
 impu	l->6	
 in 2	6->1	
 in F	r->1	
 in a	n->1	
 in b	i->2	l->1	
 in d	e->6	
 in e	t->1	
 in f	y->1	ö->2	
 in h	ä->1	
 in i	 ->25	,->1	
 in k	o->2	
 in l	i->1	
 in m	å->2	
 in n	a->1	
 in o	c->2	s->1	
 in p	a->1	å->23	
 in r	a->1	e->1	
 in s	i->3	k->1	y->1	
 in u	n->2	t->1	
 in v	a->1	e->1	å->2	
 in y	t->1	
 in, 	o->2	p->1	s->1	
 inbe	g->12	
 inbj	u->6	ö->1	
 inbl	a->14	
 inby	g->1	
 inci	d->1	t->7	
 inde	l->2	
 indi	k->5	r->7	s->1	v->14	
 indu	s->43	
 inef	f->3	
 infe	k->2	
 infi	l->1	n->2	
 infl	y->11	
 info	r->89	
 infr	a->14	i->1	
 infö	r->159	
 inga	 ->23	l->3	
 inge	n->80	r->2	t->31	
 ingi	v->6	
 ingr	e->7	i->9	
 ingå	 ->8	.->1	e->5	r->13	t->6	
 inhe	m->2	
 inhä	m->6	
 inif	r->1	
 init	i->68	
 inkl	u->21	
 inko	m->13	n->1	
 inkr	ä->1	
 inkö	p->2	r->1	
 inle	d->59	t->13	
 inlä	g->18	m->5	
 inlå	s->1	t->1	
 inlö	p->1	
 inna	n->39	
 inne	 ->5	,->1	b->116	f->6	h->81	r->4	v->2	
 inno	v->5	
 inom	 ->282	e->1	
 inpr	ä->1	
 inre	 ->81	s->3	
 inri	k->46	
 inry	m->1	
 inrä	t->54	
 insa	m->5	t->37	
 inse	 ->13	;->1	r->24	
 insi	k->4	s->6	
 insk	r->11	
 insl	a->6	
 insp	e->8	i->3	
 inst	a->7	i->122	r->45	ä->47	
 insy	n->13	
 inta	 ->4	g->4	r->4	
 inte	 ->1566	!->2	,->13	.->14	:->1	?->2	g->42	l->8	n->11	r->108	t->2	
 inti	m->1	
 into	g->2	l->4	
 intr	e->113	o->6	y->15	ä->28	å->1	
 inty	g->4	
 intä	k->2	
 inva	l->1	n->18	
 inve	c->2	n->1	r->7	s->14	
 invi	t->1	
 invo	l->9	
 invä	n->13	
 invå	n->8	
 inöv	a->1	
 irak	i->1	
 irlä	n->8	
 iron	i->2	
 irra	t->2	
 irrg	å->1	
 irri	t->4	
 is j	u->2	
 isce	n->1	
 isol	e->7	
 isra	e->19	
 istä	l->1	
 isär	 ->2	
 ital	i->17	
 itu 	m->20	
 iver	 ->2	
 iväg	 ->2	,->1	
 ja -	 ->1	
 ja e	l->1	
 ja i	 ->1	
 ja n	ä->1	
 ja t	.->1	i->2	
 ja, 	d->1	l->1	m->1	t->1	v->1	
 jag 	-->5	1->1	G->1	a->111	b->36	c->2	d->14	e->24	f->75	g->25	h->78	i->73	j->1	k->57	l->15	m->46	n->23	o->29	p->18	r->23	s->119	t->102	u->30	v->116	ä->40	å->4	ö->1	
 jag,	 ->15	
 jag.	 ->1	S->1	
 jaga	r->2	
 jakt	 ->3	
 janu	a->16	
 japa	n->1	
 jett	o->1	
 jobb	 ->2	,->2	
 joni	s->1	
 jord	 ->1	.->2	b->61	e->3	m->1	s->1	
 jour	n->2	
 ju E	g->1	
 ju M	o->1	
 ju a	b->1	l->5	n->1	t->3	v->1	
 ju b	a->2	
 ju d	e->2	i->1	ä->1	å->1	
 ju e	m->1	n->1	
 ju f	ö->2	
 ju h	ä->1	
 ju i	n->10	s->1	
 ju l	ä->1	
 ju m	e->4	å->1	
 ju o	c->7	f->1	
 ju p	a->1	o->1	å->1	
 ju r	e->2	
 ju s	a->2	i->1	t->3	
 ju t	i->1	
 ju u	t->1	
 ju v	i->1	
 ju ä	n->1	r->5	
 ju, 	o->1	p->1	
 jubl	a->1	
 juda	r->1	
 jude	u->1	
 judi	s->1	
 jul 	o->1	
 julf	e->1	
 juli	 ->8	,->2	
 julk	l->1	
 jung	f->1	
 juni	 ->12	
 juri	d->30	s->15	
 just	 ->87	:->1	e->6	i->10	
 juve	l->1	
 jämf	ö->16	
 jämk	a->1	
 jäml	i->8	
 jämn	 ->1	,->1	a->1	v->1	
 jäms	i->1	t->23	
 jämv	i->2	
 järn	-->2	v->15	
 jätt	e->1	
 kaba	r->1	
 kabi	n->3	
 kadm	i->3	
 kall	a->29	e->2	t->2	
 kam,	 ->1	
 kamm	a->58	
 kamp	 ->7	a->5	e->16	
 kamr	a->1	
 kan 	A->1	E->3	a->32	b->46	d->36	e->19	f->75	g->61	h->23	i->73	j->33	k->29	l->28	m->36	n->13	o->19	p->9	r->15	s->52	t->44	u->41	v->71	ä->5	å->12	ö->5	
 kan,	 ->3	
 kana	d->2	l->5	
 kand	i->13	
 kani	n->1	
 kano	n->1	
 kans	k->56	l->1	
 kaos	 ->2	
 kapa	c->4	d->1	
 kapi	t->20	
 kapp	 ->1	
 kapt	e->2	
 kara	k->11	
 karg	a->1	
 karr	i->1	
 kart	e->13	l->1	
 kask	a->1	
 kast	a->3	
 kata	l->4	s->61	
 kate	g->5	
 kato	l->7	
 kedj	a->3	o->1	
 kelt	i->1	
 kemi	k->5	s->1	
 kidn	a->1	
 kilo	 ->3	,->1	m->1	
 kine	s->9	
 kl. 	1->17	2->3	
 kl.1	2->1	
 klag	a->1	o->4	
 klap	p->1	
 klar	 ->12	a->24	g->17	h->7	l->5	t->78	
 klas	s->19	
 klau	s->4	
 klav	e->1	
 klib	b->1	
 klie	n->1	
 klim	a->12	
 kloa	k->1	
 kloc	k->2	
 klok	a->2	t->5	
 klyf	t->5	
 km l	å->1	
 km m	i->1	
 km, 	t->1	
 km.T	r->1	
 knap	p->16	
 knip	a->1	
 know	-->1	
 knus	s->1	
 knut	e->4	n->2	p->1	
 knyt	a->5	e->2	s->1	
 knäc	k->2	
 koal	i->12	
 kod 	h->1	k->1	
 kode	n->2	r->1	
 koff	e->1	
 kohe	r->1	
 koko	r->1	
 kol-	 ->1	
 kold	i->5	
 koll	e->199	i->3	
 kolo	s->1	
 kom 	a->1	d->2	f->6	h->1	i->3	m->2	n->1	r->1	s->1	t->2	u->1	v->1	ö->3	
 komb	i->1	
 komm	a->134	e->724	i->1082	u->25	
 komp	e->17	l->43	o->4	r->21	
 konc	e->35	i->2	
 konf	e->24	i->4	l->15	r->1	
 kong	r->1	
 konj	u->1	
 konk	r->57	u->270	
 kons	e->61	o->3	t->97	u->63	
 kont	a->20	e->1	i->7	o->7	r->145	
 konv	e->19	
 koop	e->1	
 kopi	a->1	e->1	
 kopp	l->5	
 kor,	 ->1	
 korn	a->1	
 korr	e->28	i->2	u->9	
 kort	 ->43	,->1	.->5	:->1	?->1	a->5	e->11	f->2	s->4	
 kost	a->9	h->1	n->89	s->2	
 kraf	t->71	
 kras	s->1	
 krav	 ->33	,->3	.->5	?->1	a->1	e->27	
 krea	t->3	
 kret	s->6	
 krig	 ->5	"->1	,->1	.->1	e->4	s->2	
 krim	i->7	
 krin	g->16	
 kris	 ->3	?->1	e->4	m->2	o->1	s->2	t->11	
 krit	a->1	e->15	i->46	
 kroa	t->1	
 krom	 ->1	,->1	
 krop	p->1	
 kros	s->1	
 kryp	h->3	
 krys	s->1	
 krän	k->17	
 kräv	a->31	d->4	e->42	s->55	t->2	
 krån	g->2	
 krön	a->1	
 kubi	k->1	
 kula	 ->1	.->1	
 kuli	s->1	
 kull	k->1	
 kulo	r->1	
 kult	u->107	
 kumu	l->2	
 kund	,->1	e->28	v->1	
 kung	a->15	
 kunn	a->252	i->2	
 kuns	k->15	
 kurs	 ->2	.->1	e->4	ä->1	
 kust	 ->1	b->1	e->16	l->2	m->3	o->2	r->1	v->1	
 kval	i->42	
 kvan	t->7	
 kvar	 ->19	,->2	.->2	;->1	h->3	s->8	
 kves	t->3	
 kvic	k->3	
 kvin	n->59	
 kvot	 ->3	!->1	,->1	e->6	
 kväl	l->9	
 kväv	a->2	
 kyla	.->1	n->1	
 kyli	g->1	
 käll	a->5	o->4	
 kämp	a->5	
 känd	,->1	.->1	a->4	e->1	
 känn	a->5	e->52	s->1	
 käns	l->35	
 känt	 ->7	,->1	
 kära	 ->53	
 käre	 ->1	
 kärl	 ->1	e->2	
 kärn	a->4	e->8	f->2	k->21	p->4	s->4	t->2	v->8	
 köks	b->1	
 köl 	n->1	
 köl,	 ->1	
 köla	r->1	
 köld	b->1	g->1	
 köne	n->3	
 köns	g->1	
 köp 	a->1	
 köpa	r->1	
 köpe	r->1	
 köpk	r->1	
 köps	l->1	
 köpt	 ->1	
 kör 	ö->1	
 köra	 ->1	s->1	
 körn	i->1	
 körs	 ->2	
 kört	 ->2	
 kött	 ->1	k->1	
 l'ea	u->1	
 la L	o->1	
 labo	r->3	
 lade	 ->11	s->6	
 lag 	i->1	s->1	v->1	ä->1	
 lag,	 ->4	
 lag.	D->2	F->1	
 laga	r->13	
 lagd	 ->1	
 lage	n->6	r->1	t->1	
 lagf	ö->5	
 lagl	i->6	
 lago	m->1	
 lagr	a->1	
 lags	t->115	
 lagt	 ->38	e->2	s->18	
 land	 ->67	,->8	.->13	e->23	s->52	v->2	
 lans	e->4	
 lant	l->1	
 lapp	a->1	v->2	
 larm	r->2	s->2	
 larv	e->1	
 last	 ->1	.->1	e->4	n->1	
 law,	 ->1	
 law.	M->1	
 le b	é->1	
 le p	a->1	
 led 	i->1	
 leda	 ->36	m->114	n->4	r->12	s->1	
 ledd	a->1	e->10	
 lede	r->32	
 ledn	i->15	
 leds	e->2	t->2	
 lega	l->13	t->2	
 legi	t->18	
 lejd	a->1	
 leke	r->1	
 lekt	i->1	
 lem.	M->1	
 leml	ä->1	
 leta	r->1	
 lett	 ->10	
 leva	 ->10	n->3	
 levd	e->1	
 leve	b->1	l->1	r->13	
 levn	a->6	
 levt	 ->1	
 liba	n->1	
 libe	r->25	
 lice	n->1	
 lida	 ->1	
 lide	r->7	
 lidi	t->3	
 liga	?->1	
 ligg	a->12	e->63	
 lika	 ->47	.->2	b->1	d->2	l->1	r->4	s->2	
 likg	i->2	
 likh	e->16	
 likn	a->20	
 likr	i->3	
 liks	o->47	t->2	
 likt	 ->2	
 likv	ä->8	
 lill	a->4	f->1	
 linb	a->1	
 lind	a->2	r->4	
 linj	e->12	
 lino	r->1	
 list	a->10	i->2	
 lita	 ->2	d->1	r->5	
 lite	 ->5	n->21	t->30	
 litt	e->8	
 liv 	f->2	i->1	o->2	s->2	
 liv,	 ->3	
 liv.	A->1	D->1	M->1	
 live	t->10	
 livs	c->3	d->2	k->6	m->88	u->1	v->1	
 ljud	e->1	l->1	
 ljug	e->1	
 ljus	 ->1	.->1	e->8	
 lobb	y->5	
 lock	a->2	
 logi	k->6	s->7	
 loja	l->5	
 loka	l->42	
 lopp	 ->2	
 loss	 ->1	n->1	
 lott	 ->1	a->3	
 lov 	a->1	i->1	
 lova	 ->2	d->3	r->1	t->5	
 lovo	r->2	
 lovv	ä->2	
 lovy	t->1	
 luck	a->3	o->2	
 ludd	i->2	
 luft	b->1	o->1	
 lugn	 ->1	a->5	
 lukt	a->1	
 lunc	h->1	
 lura	s->1	t->1	
 luta	 ->1	
 luth	e->1	
 lyck	a->48	l->5	o->1	ö->5	
 lyda	 ->2	
 lyde	r->3	
 lyft	 ->2	a->4	e->2	
 lykt	a->1	
 lysa	 ->2	n->4	
 lyss	n->29	
 läck	o->1	t->3	
 läge	 ->8	,->1	.->1	r->1	s->3	t->7	
 lägg	a->82	e->33	n->1	s->14	
 lägl	i->1	
 lägr	e->10	
 lägs	t->1	
 läka	r->4	
 läke	m->1	
 lämn	a->56	
 lämp	l->46	
 länd	e->114	
 läng	d->1	e->35	r->62	s->2	t->1	
 länk	a->1	
 lär 	e->1	
 lära	 ->5	r->2	
 lärd	e->1	o->7	
 läro	a->1	s->1	
 lärt	 ->2	
 läs 	y->1	
 läsa	 ->3	
 läsb	a->2	
 läse	r->6	
 läsf	r->1	
 läsk	u->1	
 läst	 ->4	e->1	
 lät 	d->1	m->1	s->3	
 lätt	 ->9	.->2	a->21	f->1	i->2	v->2	
 läxa	n->1	t->1	
 låg 	a->1	d->1	h->1	i->1	n->2	t->1	
 låga	 ->5	
 lågt	 ->2	
 lång	 ->30	,->1	.->1	a->9	d->1	f->2	r->1	s->13	t->52	v->6	
 låse	r->1	
 låst	 ->1	a->1	
 låt 	e->1	m->5	o->8	
 låta	 ->27	
 låte	r->6	
 låti	t->1	
 låts	a->2	
 löft	e->11	
 löje	v->3	
 lökm	o->1	
 lön 	f->1	
 löne	-->1	a->1	
 löns	a->5	
 lönt	 ->1	a->3	
 löpa	 ->1	n->5	
 löpe	r->7	
 löpt	 ->5	e->2	
 lörd	a->1	
 lös 	e->1	
 lösa	 ->28	.->1	s->5	
 löse	r->1	
 lösg	ö->1	
 lösn	i->48	
 lösr	y->1	
 löst	 ->2	a->3	e->1	s->1	
 lövs	k->1	
 m.m.	O->1	
 mage	r->1	
 magn	i->1	
 main	s->5	
 maj 	1->3	2->1	f->1	
 maj,	 ->1	
 maj.	J->1	T->1	
 majo	r->38	
 makr	o->6	
 makt	 ->13	,->2	.->4	b->4	d->2	e->5	f->1	h->1	k->1	l->3	m->3	
 malt	e->3	
 man 	"->1	E->1	a->35	b->31	d->22	e->13	f->28	g->20	h->39	i->86	j->5	k->40	l->16	m->26	n->14	o->19	p->14	r->13	s->86	t->30	u->17	v->37	y->1	ä->14	å->6	ö->7	
 man,	 ->13	
 man.	D->1	
 mana	r->1	t->1	
 mand	a->23	
 mani	f->1	
 manl	i->1	
 mann	e->1	
 mant	r->2	
 marg	i->5	
 mari	t->3	
 mark	 ->5	a->3	e->9	n->171	
 mars	 ->5	,->3	.->2	c->1	
 mask	e->1	i->3	
 maso	c->1	
 mass	a->5	i->3	m->3	
 mast	o->1	
 matc	h->1	
 mate	m->1	r->25	
 matn	y->1	
 matp	e->1	
 matt	a->2	
 maxb	e->1	
 maxi	m->7	
 med 	"->3	-->1	1->6	2->8	3->2	5->1	8->1	A->3	B->2	D->2	E->19	F->4	G->1	H->4	I->3	J->1	K->2	L->3	M->4	O->2	P->1	R->1	S->5	T->3	U->4	V->2	a->193	b->21	d->250	e->133	f->83	g->19	h->52	i->36	j->3	k->50	l->13	m->66	n->38	o->44	p->48	r->37	s->118	t->73	u->29	v->51	y->5	Ö->2	ä->8	å->6	ö->12	
 med,	 ->12	
 med.	D->3	F->1	V->2	
 meda	n->22	r->2	
 medb	e->15	o->155	r->1	
 medd	e->57	
 mede	l->96	
 medf	i->2	ö->20	
 medg	e->18	i->2	
 medh	j->1	
 medi	a->5	c->1	e->5	n->1	
 medk	ä->5	
 medl	e->339	i->4	
 medv	e->57	
 mega	p->1	
 meka	.->1	n->8	
 mell	a->199	
 men 	A->1	E->1	F->1	I->1	a->16	b->6	d->97	e->11	f->11	g->2	h->3	i->27	j->40	k->2	l->1	m->14	n->11	o->35	r->2	s->29	t->11	u->3	v->44	ä->13	ö->1	
 men,	 ->4	
 mena	d->2	r->27	s->2	
 meni	n->47	
 mer 	B->1	a->10	b->4	d->14	e->12	f->9	g->2	h->2	i->5	k->12	l->7	m->8	n->1	o->8	p->11	r->4	s->11	t->6	u->3	v->5	ä->34	ö->4	
 mer!	"->2	
 mer,	 ->2	
 mer.	 ->1	B->1	D->2	K->1	V->2	
 mera	 ->11	
 merg	e->1	
 meri	t->1	
 merp	a->1	
 merv	ä->5	
 mest	 ->39	a->5	
 meta	l->4	
 meto	d->23	
 midd	a->1	
 mig 	a->39	b->9	d->8	e->6	f->13	g->4	h->5	i->15	k->3	l->2	m->10	n->5	o->25	p->11	r->1	s->12	t->8	u->5	v->12	y->1	ä->8	å->6	ö->2	
 mig!	"->1	
 mig,	 ->15	
 mig.	D->1	E->1	J->3	
 mig:	 ->1	
 mig?	V->1	
 migr	a->2	
 mikr	o->4	
 mild	a->1	r->3	
 mili	s->1	t->8	
 milj	a->15	o->62	ö->184	
 mill	e->7	
 mils	t->1	
 min 	a->2	b->5	d->5	e->5	f->14	g->23	i->1	k->25	m->19	o->3	p->5	r->8	s->3	t->5	u->15	v->2	å->9	ö->2	
 min,	 ->1	
 mina	 ->72	
 mind	r->52	
 mini	m->26	r->1	s->39	
 minn	a->2	e->12	s->6	
 mino	r->22	
 mins	k->62	t->31	
 minu	s->5	t->16	
 mira	k->1	
 miss	a->1	b->9	f->5	g->7	h->1	i->1	k->6	l->18	n->3	t->23	u->2	
 mist	e->2	
 misä	r->2	
 mitt	 ->68	e->2	
 mix.	D->1	
 mjuk	a->1	
 mobi	l->7	
 mod 	a->1	f->1	i->1	s->1	
 mode	l->9	r->40	t->6	
 modi	f->3	g->3	
 moge	n->1	t->1	
 moms	p->1	
 mone	t->7	
 moni	t->1	
 mono	k->3	p->16	
 mons	t->1	
 mont	e->1	
 mora	l->6	
 mord	 ->3	,->1	.->1	b->1	e->1	i->1	
 morg	o->36	
 mors	e->6	
 mot 	1->1	5->1	A->1	D->1	E->8	F->3	G->1	H->3	M->1	S->1	a->19	b->18	d->40	e->18	f->8	g->2	h->3	i->2	k->5	l->1	m->7	n->4	o->6	p->5	r->9	s->15	t->2	u->3	v->9	Ö->2	å->1	ö->4	
 mot,	 ->1	
 mota	r->1	
 motg	å->1	
 moti	v->21	
 moto	r->8	
 motp	a->4	
 mots	a->23	t->16	v->17	ä->17	
 mott	a->16	
 motv	e->4	i->2	
 motå	t->3	
 mult	i->9	
 munt	l->8	
 mura	r->1	
 musi	k->4	
 muss	e->2	
 muto	r->1	
 myck	e->452	
 mygg	o->1	
 myll	r->1	
 mynd	i->109	
 mynn	a->1	
 myti	s->1	
 mäkt	a->1	i->2	
 män 	i->1	o->6	p->1	s->1	
 män.	J->1	T->1	
 mäng	d->18	
 männ	e->1	i->93	
 mäns	 ->1	k->42	
 märk	a->3	b->3	e->9	l->4	n->3	t->1	
 mäta	 ->2	r->1	
 mätt	e->1	
 må h	a->1	e->1	
 må v	a->1	
 måhä	n->5	
 mål 	1->16	2->10	5->2	a->3	b->2	e->1	f->6	h->1	i->4	j->1	l->1	n->1	o->4	p->2	r->1	s->11	u->2	ä->3	
 mål,	 ->12	
 mål-	2->1	
 mål.	D->3	E->1	F->1	H->2	I->1	J->1	K->1	M->1	N->2	
 mål:	 ->1	
 måla	r->1	
 måle	n->14	t->19	
 måli	n->4	
 målm	e->1	
 måls	ä->15	
 mån 	b->1	d->4	h->1	l->1	o->1	s->2	
 mån,	 ->1	
 måna	 ->3	d->69	
 månd	a->3	e->1	
 mång	a->141	f->17	s->3	
 mår.	H->1	
 måst	e->696	
 mått	 ->1	.->1	f->1	o->2	
 möbl	e->1	
 mödo	s->1	
 mödr	a->1	
 möjl	i->281	
 mörd	a->5	
 mörk	 ->1	l->1	
 möta	 ->6	
 möte	 ->10	n->3	r->2	s->2	t->7	
 mött	e->1	
 nack	d->6	
 naiv	a->1	i->1	
 nakn	a->1	
 namn	 ->7	,->1	.->2	e->2	u->4	
 nark	o->6	
 nati	o->177	
 natt	 ->1	e->2	
 natu	r->120	
 nazi	s->8	
 ned 	a->2	d->1	e->3	f->1	i->5	m->3	n->1	o->1	p->2	t->1	v->1	
 ned.	E->1	J->1	
 nede	r->9	
 nedg	å->2	
 nedl	a->1	ä->3	
 nedm	o->3	
 nedr	u->1	
 neds	k->4	t->3	
 nedv	ä->1	
 nega	t->26	
 nej 	l->1	t->1	
 nej,	 ->2	
 nej.	(->1	
 neka	 ->2	d->1	n->1	s->1	
 neon	a->1	l->1	
 nepo	t->5	
 ner 	f->1	o->1	s->2	v->1	
 nere	 ->2	.->1	
 neut	r->2	
 ni a	l->4	n->1	r->1	t->18	v->1	
 ni b	e->7	l->1	r->1	ä->1	
 ni d	e->2	i->1	ä->1	å->3	
 ni e	f->1	n->1	r->2	
 ni f	i->1	r->3	å->1	ö->7	
 ni g	e->2	ö->3	
 ni h	a->19	e->1	ä->2	å->2	
 ni i	 ->2	n->12	
 ni j	u->3	
 ni k	a->3	o->8	u->1	ä->5	
 ni l	e->1	ä->1	ö->1	
 ni m	e->2	å->1	
 ni n	u->2	ä->6	
 ni o	c->3	m->2	s->1	
 ni p	a->1	e->1	å->1	
 ni r	a->2	e->2	ä->1	
 ni s	a->9	e->4	j->2	k->6	l->1	o->2	t->2	ä->4	
 ni t	a->5	i->1	o->1	
 ni u	n->1	p->3	t->1	
 ni v	a->3	e->8	i->9	ä->2	å->1	
 ni ä	r->6	v->1	
 ni ö	n->1	
 ni, 	b->1	f->3	h->4	m->1	o->2	
 ni.D	ä->1	
 nimb	u->1	
 nio 	b->2	f->1	l->1	m->7	p->1	t->1	
 nion	d->1	
 nivå	 ->29	,->7	.->14	;->1	e->9	n->7	
 njut	n->1	
 nog 	a->3	b->1	d->2	h->2	i->1	k->1	n->1	o->1	p->1	ö->1	
 nog,	 ->1	
 nog.	M->2	
 noga	 ->9	,->1	.->2	
 nogg	r->12	
 noll	,->1	n->1	r->1	
 nomi	n->3	
 non 	f->2	
 nord	a->4	e->1	i->3	k->1	l->4	t->1	v->1	
 norm	a->12	e->21	
 norr	?->1	a->4	
 nota	n->1	
 note	r->28	
 nove	m->11	
 nr 1	 ->1	2->2	7->2	
 nr 2	8->1	9->1	
 nr 3	0->1	1->1	2->1	3->2	5->1	6->1	7->1	8->1	9->1	
 nr 4	0->1	1->1	2->1	3->1	4->1	5->1	6->1	
 nr 5	 ->1	
 nr 6	 ->1	
 nr 7	.->1	
 nr 8	 ->1	
 nr 9	 ->1	
 nu -	 ->1	
 nu 3	4->1	
 nu E	r->1	
 nu a	n->1	t->5	v->1	
 nu b	e->4	l->4	
 nu d	e->4	i->2	ö->1	
 nu e	f->1	g->1	n->3	t->5	u->1	
 nu f	a->2	i->3	r->2	å->3	ö->10	
 nu g	e->5	ä->3	å->3	ö->3	
 nu h	a->13	å->1	ö->1	
 nu i	 ->3	g->1	n->6	
 nu k	a->5	o->6	
 nu l	i->1	y->1	ä->3	
 nu m	e->1	ä->1	å->8	
 nu n	u->1	ä->8	
 nu o	c->4	f->2	m->1	
 nu p	l->1	r->2	å->3	
 nu r	u->1	å->2	ö->1	
 nu s	e->2	i->1	k->6	l->1	o->1	p->1	t->5	ä->2	å->1	
 nu t	a->5	i->3	y->3	
 nu u	n->1	p->3	
 nu v	a->1	e->2	i->4	
 nu ä	n->6	r->10	
 nu å	t->1	
 nu, 	e->1	i->1	m->2	u->1	ö->1	
 nu..	T->1	
 nu.J	a->1	
 nu.L	å->1	
 nu.V	i->1	
 nu: 	g->1	
 nu?J	a->1	
 null	i->1	
 nulä	g->1	
 nume	r->5	
 numm	e->2	
 nunn	o->1	
 nuva	r->45	
 ny b	i->1	
 ny e	u->1	
 ny f	a->1	o->1	ö->2	
 ny g	r->1	
 ny h	ä->1	
 ny i	n->2	
 ny k	e->1	o->3	u->3	v->1	
 ny l	a->1	e->1	i->1	
 ny m	y->1	
 ny o	c->1	l->1	
 ny p	e->2	
 ny r	ö->2	
 ny s	e->1	i->1	p->1	t->1	y->2	
 ny t	y->1	
 ny u	p->1	
 ny v	e->1	i->2	
 nya 	"->1	8->1	E->3	a->12	b->14	d->5	e->2	f->10	g->3	i->4	j->1	k->17	l->7	m->16	n->2	o->6	p->13	r->16	s->7	t->8	u->3	v->4	ä->2	å->6	
 nya,	 ->1	
 nya;	 ->1	
 nyan	s->3	
 nyas	t->1	
 nybi	l->2	
 nyck	e->7	
 nyda	n->1	
 nye 	o->1	
 nyet	a->1	
 nyfa	s->1	
 nyfö	r->1	
 nyhe	t->12	
 nykt	e->2	r->1	
 nyli	b->1	g->29	
 nyna	z->6	
 nypl	a->1	
 nysk	a->1	
 nyss	 ->10	,->2	.->1	
 nytt	 ->40	,->3	.->3	a->20	i->10	o->1	
 nyva	l->1	
 nyår	s->1	
 näml	i->43	
 nämn	a->27	d->22	e->5	s->9	t->19	v->1	
 när 	C->1	E->1	M->1	P->1	a->8	b->3	c->1	d->199	e->8	f->5	g->2	h->12	j->14	k->7	l->1	m->21	n->10	p->1	r->3	s->2	t->1	v->43	ä->2	ö->2	
 när,	 ->1	
 nära	 ->19	,->1	
 närh	e->5	
 näri	n->12	
 närm	a->36	
 närs	y->1	
 närv	a->46	
 näsd	u->1	
 näst	a->47	
 nät 	o->1	s->1	
 nät.	 ->1	
 näte	n->1	
 näts	t->1	
 nätt	e->1	
 nätv	e->11	
 nå a	n->1	
 nå d	e->2	
 nå e	n->6	t->1	
 nå f	r->4	
 nå h	ö->1	
 nå v	å->1	
 nå ä	n->1	
 nå å	t->1	
 nåba	r->2	
 nåd 	a->1	
 någo	n->165	r->1	t->191	
 någr	a->147	
 når 	d->1	e->1	
 nått	 ->7	
 nödb	e->1	
 nöde	n->1	
 nödi	n->1	
 nöds	i->1	
 nödv	ä->123	
 nöja	 ->8	k->2	
 nöjd	 ->1	a->8	
 nöje	 ->3	r->1	t->2	
 nöjt	 ->1	
 nöt.	D->1	
 nötk	ö->3	
 nöts	k->1	
 nött	e->1	
 oacc	e->31	
 oakt	a->1	
 oans	v->5	
 oanv	ä->1	
 oavb	r->2	
 oavs	e->8	i->2	
 obal	a->6	
 obeb	o->1	
 obef	o->1	
 obeg	r->5	
 obeh	a->2	
 ober	o->49	ä->1	
 obes	t->2	v->3	
 obje	k->1	
 obli	g->14	
 obse	r->2	
 och 	"->3	(->1	-->6	0->1	1->21	2->13	3->7	4->10	5->3	6->2	7->6	8->11	9->4	A->4	B->6	C->4	D->4	E->35	F->15	G->7	H->3	I->14	J->2	K->9	L->8	M->5	N->2	O->2	P->15	R->3	S->25	T->8	U->1	V->2	W->1	X->1	a->290	b->119	c->10	d->588	e->210	f->317	g->91	h->160	i->231	j->152	k->197	l->93	m->278	n->79	o->95	p->114	r->188	s->440	t->150	u->106	v->229	y->7	Ö->7	ä->54	å->37	ö->43	
 och,	 ->9	
 och/	e->1	
 ocks	å->585	
 ocku	p->5	
 odds	 ->1	
 odel	b->1	
 odis	k->1	
 odju	r->2	
 odug	l->1	
 oeft	e->1	
 oege	n->5	
 oeko	n->1	
 oeni	g->4	
 oens	e->4	
 oerh	ö->12	
 oers	ä->1	
 oeti	s->1	
 of t	h->1	
 ofan	t->2	
 ofel	b->1	
 offe	n->79	r->10	
 offi	c->5	
 offr	a->2	e->14	
 ofre	d->1	
 ofrå	n->3	
 ofta	 ->49	.->1	r->3	s->1	
 oful	l->2	
 oför	d->2	e->5	l->2	m->5	s->3	t->2	ä->2	
 ogen	o->2	
 ogru	n->2	
 ogyn	n->1	
 ohjä	l->1	
 ohäm	m->1	
 ohöv	l->1	
 oige	n->1	
 oins	k->2	
 oint	r->4	
 ojäm	l->5	n->2	
 okla	n->2	r->12	
 okon	t->2	
 okri	t->1	
 okrä	n->1	
 okto	b->8	
 okun	n->2	s->1	
 okän	d->1	s->1	
 olag	l->4	
 olik	 ->1	a->114	h->5	
 olja	 ->3	,->1	.->1	n->3	
 olje	b->13	f->1	i->3	k->2	s->1	t->10	u->2	
 olog	i->1	
 olyc	k->45	
 olym	p->1	
 oläm	p->3	
 olös	t->2	
 om "	K->1	o->1	ö->1	
 om -	 ->5	
 om 1	 ->1	5->1	6->1	9->1	
 om 2	0->1	
 om 3	-->1	1->1	5->3	
 om 4	0->2	
 om 6	,->1	
 om A	l->1	m->1	t->1	
 om B	e->1	r->1	
 om C	E->1	
 om D	u->1	
 om E	G->1	U->2	r->1	t->1	u->13	
 om F	l->1	ö->1	
 om G	U->1	e->1	o->1	r->1	
 om H	a->3	i->1	
 om I	N->1	s->1	t->1	
 om J	ö->1	
 om K	a->1	o->5	
 om L	a->3	
 om M	a->1	c->1	
 om P	o->1	
 om S	c->1	j->1	
 om T	a->1	h->1	i->2	u->3	
 om a	g->1	l->15	n->16	r->9	s->2	t->206	v->10	
 om b	a->2	e->26	i->2	o->1	r->7	u->1	ä->1	å->3	ö->1	
 om c	o->1	
 om d	a->3	e->327	i->4	o->1	r->2	ö->1	
 om e	f->2	g->1	k->2	l->1	n->72	r->8	t->38	u->3	x->4	
 om f	a->1	i->5	l->1	o->3	r->20	u->1	ö->52	
 om g	a->2	e->11	o->1	r->6	
 om h	a->19	e->1	j->3	o->6	u->32	ä->4	å->2	
 om i	 ->7	c->4	d->1	f->1	g->1	n->38	s->1	
 om j	a->23	o->2	u->1	ä->2	
 om k	a->5	e->1	o->61	r->3	u->5	ä->7	
 om l	a->3	e->2	i->17	o->1	ä->3	å->1	ö->1	
 om m	a->45	e->9	i->11	o->5	y->4	ä->12	å->1	ö->3	
 om n	a->4	e->2	i->16	y->3	ä->2	å->12	ö->1	
 om o	c->11	g->1	l->4	m->3	r->3	s->1	
 om p	a->5	e->2	o->2	r->9	å->2	
 om r	a->2	e->31	i->6	o->1	u->1	ä->9	å->11	
 om s	.->1	a->17	e->2	i->4	j->2	k->8	l->2	m->1	o->3	p->3	t->25	u->3	v->1	y->2	ä->7	å->10	
 om t	.->1	a->1	i->16	j->2	o->3	r->11	v->1	y->2	
 om u	n->4	p->5	r->5	t->30	
 om v	a->23	e->7	i->78	o->1	ä->1	å->5	
 om y	r->1	t->1	
 om Ö	s->3	
 om ä	n->11	r->1	v->1	
 om å	r->3	t->9	
 om ö	a->1	k->1	m->1	p->4	v->2	
 om".	D->1	
 om);	 ->1	
 om, 	a->3	d->4	h->2	l->1	m->2	o->3	s->2	u->1	v->1	ä->2	
 om. 	D->1	
 om.A	v->1	
 om.D	e->6	ä->1	
 om.E	K->1	x->1	
 om.I	n->1	
 om.J	a->6	
 om.M	e->3	
 om.N	ä->1	
 om.O	c->1	
 om.S	t->1	å->1	
 om.V	i->1	
 omI.	 ->1	
 omba	d->1	
 ombe	d->1	s->2	t->2	
 ombo	r->1	
 ombu	d->12	
 omde	f->1	
 omdi	r->1	
 omdö	m->2	
 omed	e->18	g->2	v->1	
 omfa	t->83	
 omfl	y->1	
 omfo	r->3	
 omfå	n->2	
 omfö	r->1	
 omge	r->1	
 omgi	v->1	
 omgå	e->1	n->2	
 omhu	l->1	
 omis	t->1	
 omkr	i->15	
 omla	s->1	
 omlo	k->2	
 ommö	b->1	
 omor	a->1	g->2	
 ompl	a->1	
 ompr	ö->8	
 omri	n->1	
 områ	d->222	
 omrö	s->35	
 omso	r->9	
 omst	r->12	ä->35	
 omsv	e->1	
 omsä	t->8	
 omta	l->1	
 omva	n->5	
 omvä	g->2	l->4	n->5	x->1	
 omöj	l->16	
 ond 	c->1	
 onda	 ->3	
 ondo	.->1	
 onds	k->1	
 one-	s->1	
 onsd	a->5	
 ont 	o->1	
 ont.	S->1	
 onöd	i->11	
 opar	t->2	
 oper	a->11	e->1	
 opin	i->4	
 oppo	n->3	r->2	s->2	
 opra	k->1	
 opro	p->2	
 opti	m->7	o->1	
 ord 	a->4	e->1	f->6	i->4	j->1	k->2	m->1	n->1	o->8	s->5	t->4	v->3	
 ord,	 ->2	
 ord.	V->1	
 ord:	 ->2	
 orda	l->6	
 orde	n->20	t->17	
 ordf	ö->193	
 ordl	i->1	
 ordn	a->1	i->21	
 ordr	e->1	i->2	
 ordv	r->1	ä->1	
 orea	l->2	
 ored	l->1	
 oreg	l->1	
 orga	n->69	
 orie	n->5	
 orig	i->2	
 orik	t->3	
 orim	l->5	
 orka	n->3	
 orm 	s->1	
 orme	n->1	
 oro 	-->1	E->1	b->1	d->1	f->5	i->3	l->1	n->2	o->4	p->1	s->12	ä->3	ö->1	
 oro,	 ->4	
 oro.	A->1	B->1	F->2	J->2	O->1	T->1	V->1	
 oroa	 ->3	d->5	n->9	r->4	
 orol	i->6	
 oron	 ->5	
 oros	m->4	
 orov	ä->2	
 orsa	k->29	
 ort,	 ->1	
 ort.	D->1	
 orwe	l->1	
 oräk	n->1	
 orät	t->10	
 osan	n->1	
 oss 	-->1	a->39	b->1	d->18	e->16	f->16	g->4	h->6	i->29	k->3	l->3	m->12	n->6	o->29	p->13	r->2	s->29	t->16	u->8	v->13	y->1	ä->10	å->10	ö->3	
 oss,	 ->15	
 oss.	D->3	E->2	F->2	H->1	J->4	N->1	V->3	Ä->2	
 oss:	 ->1	
 oss?	.->1	V->1	
 ostr	o->3	
 osv.	 ->3	,->1	?->1	S->1	
 osyn	l->1	
 osäk	e->8	
 osår	b->1	
 otac	k->1	
 otil	l->17	
 otjä	n->1	
 otro	l->2	
 otry	g->1	
 otve	t->2	
 otvi	v->1	
 otyd	l->4	
 otän	k->1	
 otål	i->1	
 oumb	ä->4	
 ound	g->2	v->4	
 outh	ä->2	
 outn	y->1	
 ovan	a->1	i->1	l->1	n->2	p->1	s->1	
 over	h->1	
 ovil	j->2	l->1	
 ovis	s->1	
 oväd	e->1	r->1	
 oväl	k->1	
 oväs	e->1	
 oänd	l->4	
 oöns	k->1	
 oöve	r->6	
 p.g.	a->1	
 pake	t->2	
 pakt	e->1	
 pale	s->12	
 papp	e->5	
 par 	a->3	b->1	g->1	m->2	o->1	p->4	s->2	å->2	
 para	d->6	g->1	l->5	m->2	
 parc	o->1	
 park	e->3	
 parl	a->389	
 part	e->19	i->67	n->25	
 pas 	l->1	
 pass	 ->4	a->7	e->3	i->2	u->1	
 pate	t->1	
 pati	e->2	
 pean	u->1	
 peda	g->1	
 pedo	f->1	
 peka	 ->6	d->3	r->6	t->4	
 pela	r->8	
 peng	a->55	
 penn	d->1	i->10	
 pens	i->6	
 per 	b->2	c->10	d->1	i->1	j->1	k->2	l->1	m->2	s->1	å->3	
 perf	e->7	
 peri	f->5	o->55	
 perm	a->8	
 perr	o->1	
 pers	o->103	p->15	
 pess	i->2	
 pest	e->4	
 peti	t->1	
 phar	m->1	
 phta	l->1	
 pilo	t->3	
 pion	j->1	
 pira	t->1	
 plac	e->14	
 plan	 ->7	,->1	:->1	e->71	t->1	
 plas	t->5	
 plat	s->31	
 plen	a->4	u->5	
 plik	t->5	
 plim	s->1	
 plun	d->1	
 plur	a->1	
 plus	 ->2	
 pläd	e->2	
 plån	b->1	
 plöt	s->4	
 poet	 ->1	
 pole	 ->1	m->1	
 poli	c->2	s->14	t->323	
 pool	,->1	
 popu	l->5	
 pors	l->1	
 port	-->2	m->1	u->70	v->1	
 posi	t->80	
 post	 ->1	v->1	
 pote	n->5	
 poän	g->12	
 prac	k->1	
 prag	m->1	
 prak	t->32	
 prat	a->4	
 prax	i->7	
 prec	i->43	
 pref	e->3	
 prej	u->4	
 prel	i->3	
 prem	i->10	
 prer	o->1	
 pres	e->28	i->8	s->18	t->4	
 pric	k->2	
 prim	i->1	
 prin	c->113	
 prio	r->36	
 pris	 ->4	.->1	a->1	e->13	n->1	s->1	u->1	
 priv	a->21	i->7	
 prob	l->156	
 proc	e->134	
 prod	u->62	
 prof	e->7	i->3	
 prog	r->153	
 proj	e->54	
 prok	l->1	
 pron	a->1	
 prop	a->4	o->7	
 pros	t->1	
 prot	e->13	o->18	
 prov	 ->9	i->5	k->1	
 präg	l->4	
 pröv	a->3	n->3	o->1	
 psyk	o->1	
 publ	i->7	
 pump	a->2	
 pund	 ->2	.->1	
 punk	t->168	
 puri	t->1	
 pyra	m->1	
 på -	 ->5	
 på 1	0->1	3->2	4->1	
 på 2	0->3	2->1	
 på 3	3->1	4->1	7->1	
 på 4	0->1	
 på 5	 ->1	0->2	
 på 7	,->1	5->1	
 på 8	0->2	6->1	
 på 9	0->1	5->1	
 på A	l->2	t->1	
 på B	S->1	a->5	e->1	
 på C	E->1	S->1	
 på E	G->3	U->4	r->1	u->10	
 på F	ö->1	
 på G	e->1	o->1	
 på H	o->1	
 på I	S->1	n->6	r->1	s->1	
 på M	a->1	
 på O	l->1	
 på P	a->1	
 på R	i->2	o->1	
 på T	y->1	
 på V	ä->2	
 på a	c->1	k->1	l->29	n->16	r->11	s->1	t->145	v->1	
 på b	a->3	e->8	i->5	l->1	o->3	r->7	ä->9	å->3	
 på c	e->1	i->1	r->1	
 på d	a->8	e->291	i->2	j->7	u->4	y->1	
 på e	f->2	g->3	k->2	l->1	m->1	n->55	r->5	t->142	u->12	x->1	
 på f	a->3	e->4	i->2	l->3	r->12	y->2	ä->6	ö->64	
 på g	a->1	e->16	l->1	o->2	r->79	ä->1	å->5	ö->1	
 på h	a->5	e->1	j->1	u->14	ä->1	ö->1	
 på i	 ->4	c->1	l->1	n->19	t->1	
 på j	a->1	o->1	u->2	ä->3	
 på k	a->5	l->2	n->1	o->36	r->1	u->1	v->1	ä->1	ö->1	
 på l	a->12	i->3	o->3	ä->6	å->9	ö->1	
 på m	a->12	e->19	i->28	o->6	y->2	ä->1	å->5	ö->4	
 på n	a->4	e->1	o->4	y->26	ä->8	å->21	
 på o	b->2	c->4	l->4	m->19	n->2	r->2	s->5	
 på p	a->1	e->3	l->9	o->1	r->9	
 på r	a->2	e->26	i->2	y->1	ä->11	å->7	
 på s	a->22	e->11	i->31	j->1	k->6	l->1	m->1	n->1	o->1	p->10	t->13	u->2	v->1	y->4	ä->5	å->16	
 på t	a->7	e->4	i->9	j->1	o->10	r->10	v->7	ä->1	
 på u	n->8	p->3	t->5	
 på v	a->16	e->8	i->16	ä->34	å->16	
 på y	t->1	
 på z	i->1	
 på Ö	s->2	
 på ä	n->6	r->3	
 på å	h->1	r->1	t->5	
 på ö	k->1	n->1	p->5	v->1	
 på, 	e->2	f->1	h->1	l->1	m->3	n->1	o->5	v->1	ä->1	
 på.B	e->1	
 på.D	e->3	o->1	
 på.E	n->1	u->1	
 på.J	a->3	
 på.N	o->1	
 på.O	r->1	
 på.U	n->1	
 på.V	i->1	
 på.Ä	r->2	
 på: 	f->2	Ö->1	
 på?.	 ->1	
 på?J	a->1	
 påbj	u->1	
 påbö	r->11	
 pådr	a->1	
 påfr	e->1	
 påfö	l->3	
 pågi	c->3	
 pågå	 ->1	e->6	r->10	t->1	
 påla	g->1	
 påli	t->1	
 pålä	g->1	
 påmi	n->30	
 påpe	k->49	
 påsk	y->7	
 påst	r->1	å->20	
 påta	g->4	l->5	
 påtr	y->3	
 påtv	i->4	
 påve	r->36	
 påvi	s->3	
 qua 	n->2	
 quo 	s->1	
 quo,	 ->1	
 rad 	a->1	b->2	d->2	f->3	g->1	i->2	k->1	m->1	n->1	o->2	p->2	r->1	s->1	
 rade	n->1	r->3	
 radi	k->16	o->2	
 rak 	k->1	
 raka	 ->2	
 rakr	y->1	
 rakt	 ->3	
 ram 	-->1	f->2	p->1	s->4	v->1	
 ram,	 ->2	
 ram.	D->1	T->1	
 rama	r->3	v->3	
 rame	n->58	
 ramp	r->11	
 ramv	i->3	
 rand	o->14	
 rann	s->1	
 rapp	o->98	
 rasa	d->2	t->1	
 rash	a->1	
 rasi	s->25	
 rati	f->13	o->7	
 reag	e->16	
 reak	t->20	
 real	i->14	
 reci	r->1	
 recy	c->1	
 reda	 ->5	k->1	n->155	r->4	s->1	
 rede	r->2	
 redl	i->1	
 redo	 ->3	g->10	v->4	
 reds	k->1	
 redu	c->4	
 reel	l->4	
 refe	r->4	
 refl	e->7	
 refo	r->127	
 rege	l->46	r->267	
 regi	,->1	m->1	o->234	s->17	
 regl	e->89	
 reha	b->1	
 rejä	l->3	
 rekl	a->2	
 reko	m->39	n->3	r->2	
 rekr	y->1	
 rela	t->23	
 rele	v->9	
 reli	g->4	k->1	
 remi	s->1	
 ren 	b->1	d->1	n->1	o->1	
 rena	 ->2	
 reng	ö->1	
 reno	v->3	
 rens	a->3	n->5	
 rent	 ->21	a->1	
 repa	r->5	
 repr	e->16	
 repu	b->10	
 resa	 ->5	,->1	.->1	
 rese	r->9	
 resi	d->1	
 reso	l->93	n->4	r->1	
 resp	.->2	e->80	o->1	
 rest	 ->2	a->1	e->3	r->4	s->1	
 resu	l->103	r->44	
 reto	r->3	
 retr	o->11	ä->1	
 revi	d->17	s->18	
 revo	l->1	
 rida	 ->1	
 righ	t->1	
 rigo	r->4	
 rika	 ->5	,->1	r->2	s->3	
 rike	d->8	t->2	
 rikl	i->2	
 rikt	 ->1	a->25	i->35	l->69	n->24	p->2	
 riml	i->18	
 rimm	a->1	
 ring	a->6	
 ris,	 ->1	
 ris:	 ->1	
 risk	 ->9	,->1	a->3	b->4	e->49	f->4	h->6	k->3	n->1	u->1	v->3	
 ro i	 ->1	
 ro, 	o->1	s->1	
 rock	s->1	
 roli	g->1	
 roll	 ->42	,->11	.->8	e->3	
 rome	r->5	
 ropa	r->2	
 rope	t->1	
 ros 	f->1	o->1	
 rose	n->1	
 rost	b->1	
 rota	t->1	
 rots	y->1	
 rubb	a->3	
 rubr	i->1	
 ruin	e->1	
 rull	a->3	s->3	
 rum 	e->1	f->1	h->1	i->15	o->3	p->3	u->2	y->1	
 rum,	 ->1	
 rum.	 ->1	D->1	M->1	O->1	
 rund	a->2	r->2	
 runt	 ->4	.->1	o->1	
 rusa	 ->1	r->2	
 rust	a->1	n->1	
 ruti	n->7	
 rutt	n->2	
 ryck	t->1	
 rygg	e->3	r->1	
 rykt	b->1	e->7	
 rymm	a->1	
 rysk	 ->1	a->1	
 ryss	a->1	
 räck	a->9	e->20	s->1	t->1	v->3	
 rädd	 ->4	,->1	a->11	n->4	
 räds	l->8	
 räke	n->8	
 räkn	a->37	e->1	i->10	
 räta	s->1	
 rätt	 ->82	,->6	.->4	?->1	a->17	e->23	f->8	i->100	m->1	s->184	v->63	ä->1	
 råd 	a->1	b->1	f->2	n->1	o->4	s->2	
 råd,	 ->1	
 råd.	J->1	M->1	
 råd?	Ä->1	
 råda	 ->7	n->3	
 rådd	e->1	
 råde	n->1	r->24	t->283	
 rådf	r->6	
 rådg	i->12	ö->1	
 råds	b->1	l->3	m->3	o->19	t->1	
 råga	t->1	
 råka	r->1	
 råol	j->1	
 rått	o->1	
 réfé	r->1	
 röda	 ->2	
 rödg	r->1	
 rör 	E->1	a->2	b->1	d->5	f->5	i->1	j->1	p->3	s->14	t->1	u->2	v->1	
 röra	 ->2	n->23	s->1	
 rörd	e->1	
 röre	l->5	
 röri	g->2	
 rörl	i->24	
 rört	 ->1	
 röst	 ->9	,->2	.->2	a->89	e->5	f->7	r->3	v->3	
 rött	 ->1	e->4	
 röva	t->1	
 s.k.	 ->4	
 sa a	t->1	
 sade	 ->55	,->14	.->5	:->1	
 safe	t->1	
 sagt	 ->28	,->8	.->1	s->12	
 sak 	a->4	g->3	h->2	j->1	k->1	m->3	n->1	s->9	t->2	v->5	ä->1	
 sak,	 ->2	
 sak.	A->1	D->1	T->1	
 sak:	 ->1	
 sake	n->11	r->31	
 sakf	ö->1	
 sakk	u->2	
 sakl	i->1	
 sakn	a->35	
 sako	m->2	
 sakp	r->1	
 sali	n->1	
 salu	f->1	
 sama	r->80	
 samb	a->47	
 same	x->2	
 samf	i->1	u->5	ö->7	
 samh	ä->42	
 saml	a->19	e->1	i->1	
 samm	a->275	
 samo	r->37	
 samr	å->9	
 sams	t->4	y->3	
 samt	 ->53	a->11	i->53	l->25	y->6	
 samv	e->5	
 sank	t->7	
 sann	 ->1	a->1	e->4	i->3	o->7	
 sans	a->2	
 sant	 ->10	!->1	,->2	.->1	:->1	
 sate	l->1	
 sats	a->13	n->4	
 satt	 ->6	,->1	a->1	e->6	
 scen	 ->1	a->4	e->1	
 scha	b->1	
 scie	n->1	
 scor	e->1	
 se a	t->12	
 se b	a->1	
 se d	e->8	
 se e	n->1	t->3	
 se f	r->4	ö->1	
 se h	o->2	u->3	ä->1	
 se i	 ->5	
 se k	o->1	
 se m	e->2	
 se n	ä->1	
 se o	m->6	
 se p	e->1	å->7	
 se r	e->1	i->1	
 se s	i->1	k->1	n->2	p->1	
 se t	i->68	
 se u	p->2	t->3	
 se v	a->1	e->1	i->7	
 se ä	n->1	
 se ö	v->10	
 seda	n->101	
 sede	r->1	
 seg 	t->1	
 segd	r->1	
 sege	r->4	
 segl	a->13	
 segr	a->1	
 seis	m->2	
 seke	l->4	
 sekl	e->2	
 sekr	e->12	
 sekt	o->47	
 seku	n->3	
 sele	k->1	
 seme	s->4	
 semi	n->1	
 sen 	a->1	
 sena	r->29	s->67	t->1	
 senf	ä->1	
 sens	i->1	
 sent	 ->2	,->1	.->3	
 sepa	r->1	
 sept	e->15	
 ser 	a->2	d->10	e->3	f->12	h->3	i->3	j->4	m->5	o->3	p->2	r->2	s->3	t->8	u->4	v->5	ä->1	ö->1	
 serb	,->1	e->7	i->6	
 seri	ö->7	
 serv	a->1	i->6	
 ses 	m->1	s->4	ö->5	
 sess	i->6	
 sett	 ->40	,->2	.->5	:->1	s->1	
 sex 	a->2	e->1	m->11	p->1	t->1	ö->1	
 sex,	 ->1	
 sexi	s->1	
 sexm	å->1	
 sext	o->1	
 sexu	e->2	
 sexv	ä->1	
 sida	 ->13	,->9	.->8	?->1	n->43	
 sido	e->1	r->6	
 siff	r->17	
 sig 	E->1	O->1	a->43	b->11	d->14	e->18	f->36	g->4	h->4	i->39	j->1	k->2	l->2	m->27	n->7	o->34	p->27	r->2	s->25	t->26	u->9	v->11	ä->5	å->13	ö->4	
 sig,	 ->8	
 sig.	A->1	B->1	D->2	E->2	H->2	J->2	K->1	M->1	S->1	T->1	V->3	Ä->1	
 sig;	 ->1	
 sign	a->12	e->1	
 sikt	 ->15	,->4	.->3	a->2	e->3	
 simm	a->1	
 simu	l->2	
 sin 	a->5	b->10	d->6	e->14	f->12	g->2	h->16	i->3	k->2	l->3	m->5	n->8	o->6	p->8	r->17	s->17	t->4	u->9	v->5	w->1	å->2	ö->1	
 sina	 ->138	
 sine	 ->3	
 sinn	a->1	e->4	
 sino	m->1	
 sins	e->3	
 sist	 ->8	,->4	a->43	n->2	
 sitt	 ->94	,->1	a->1	e->6	n->2	
 situ	a->116	
 sju 	g->1	m->1	p->1	r->1	
 sju,	 ->1	
 sjuk	.->1	d->1	f->1	h->6	v->3	
 sjun	d->4	k->9	
 sjut	t->2	
 själ	,->1	.->2	e->2	v->168	
 sjät	t->19	
 sjöf	a->7	
 sjöm	ä->2	
 sjön	.->1	k->4	
 sjös	s->4	
 sjöt	r->1	
 sjöv	ä->1	
 ska 	g->1	v->1	
 skad	a->25	e->3	l->7	o->21	
 skaf	f->5	
 skak	a->2	
 skal	a->1	d->1	l->670	
 skam	 ->2	!->1	l->2	m->1	p->1	
 skan	d->7	
 skap	a->175	
 skar	 ->1	a->1	p->2	
 skat	t->33	
 ske 	-->1	e->3	g->2	i->2	m->1	p->5	s->1	u->2	
 ske!	Ä->1	
 ske,	 ->1	
 sked	e->4	
 skep	p->8	s->1	t->5	
 sker	 ->27	.->4	
 sket	t->15	
 skic	k->16	
 skil	d->5	j->14	l->42	
 skin	g->1	
 skip	a->2	
 skis	s->4	
 skju	t->25	
 skog	 ->3	a->8	e->5	r->1	s->19	
 skol	a->6	o->2	
 skon	a->1	
 skra	t->2	
 skre	v->5	
 skri	d->1	f->8	k->1	v->20	
 skro	t->24	v->5	
 skrä	c->3	d->1	m->4	
 skug	g->3	
 skul	d->2	l->496	
 skur	a->1	
 skut	a->3	
 skyd	d->74	
 skyf	a->1	
 skyh	ö->1	
 skyl	d->26	l->3	
 skym	t->1	
 skyn	d->7	
 skäl	 ->29	,->1	.->2	e->10	i->1	
 skäm	m->2	t->1	
 skän	k->2	
 skär	 ->2	p->11	s->1	
 skåd	a->2	
 skön	h->1	
 skör	.->1	a->2	d->3	
 sköt	 ->2	a->7	e->1	s->3	t->4	
 sköv	l->1	
 slag	 ->14	.->2	e->2	i->1	s->15	
 slak	t->1	
 slam	 ->1	
 slap	p->3	
 slav	a->1	
 slip	p->2	
 slir	a->1	
 slit	a->1	
 slog	 ->2	
 slot	t->1	
 slov	e->1	
 sluk	a->3	
 slum	p->4	r->1	
 slus	s->2	
 slut	 ->19	,->4	.->3	a->11	e->26	f->9	g->8	h->1	i->2	k->1	l->38	n->1	p->1	r->2	s->40	v->1	ä->5	
 släc	k->3	
 släk	t->1	
 släp	a->1	p->9	
 slå 	f->6	i->1	s->1	v->2	
 slåe	n->1	
 slår	 ->2	.->1	
 slås	s->1	
 slös	a->2	e->2	
 smak	ä->1	
 smid	i->3	
 smit	a->1	n->1	
 smul	a->1	
 smus	s->1	
 smut	s->3	
 smäd	e->1	
 smär	r->1	t->2	
 små 	E->1	a->1	b->1	e->1	f->4	l->2	m->4	o->32	p->1	s->5	å->1	
 små,	 ->2	
 små.	D->1	
 småf	ö->5	
 småg	r->1	
 smån	i->4	
 smås	k->1	
 snab	b->71	
 snar	 ->2	a->36	l->1	t->27	
 sned	v->12	
 snäl	l->1	
 snäv	a->1	
 snår	i->1	
 snöv	i->1	
 so f	a->1	
 soci	a->199	e->1	o->3	
 soft	 ->1	
 sola	 ->1	
 sold	a->2	
 soli	d->30	
 sols	k->1	
 som 	"->3	-->3	1->1	2->1	4->2	A->3	B->9	C->2	D->3	E->38	F->3	G->3	H->3	I->2	J->3	L->4	M->2	N->1	P->3	R->3	S->3	T->2	W->1	a->112	b->149	c->4	d->158	e->149	f->262	g->126	h->283	i->211	j->100	k->178	l->97	m->168	n->88	o->63	p->60	r->100	s->259	t->95	u->87	v->290	y->1	Ö->1	ä->196	å->17	ö->13	
 som,	 ->21	
 soml	i->3	
 somm	a->3	
 sopa	 ->1	
 sorg	 ->1	l->3	
 sort	e->1	s->7	
 sovj	e->1	
 span	j->1	s->10	
 spar	a->5	k->3	s->1	
 spec	i->84	
 speg	l->3	
 spek	t->5	u->2	
 spel	 ->5	,->2	.->2	;->1	a->34	e->2	p->1	r->5	
 spen	d->5	
 spet	s->2	
 spil	l->1	
 spli	t->3	
 spon	s->1	t->4	
 spor	t->1	
 spot	s->1	
 spri	d->15	
 språ	k->8	n->1	
 spän	n->10	
 spär	r->3	
 spår	 ->3	,->1	a->3	e->1	
 spök	e->3	s->1	
 sril	a->1	
 stab	 ->1	i->22	
 stac	k->1	
 stad	 ->1	.->1	g->26	i->5	s->3	
 stag	n->2	
 stal	i->2	
 stan	d->21	n->7	
 star	k->60	t->15	
 stat	 ->11	,->2	.->3	e->73	i->9	l->79	s->33	u->7	
 stee	r->1	
 steg	 ->33	,->1	e->1	
 stel	a->2	t->1	
 sten	 ->1	d->1	k->1	
 ster	i->1	
 stic	k->5	
 stif	t->1	
 stig	a->2	e->1	i->2	m->1	
 stil	 ->1	l->3	
 stim	u->11	
 stod	 ->5	
 stol	t->11	
 stop	p->18	
 stor	 ->102	.->1	a->117	d->2	e->1	f->2	h->1	k->1	m->27	s->4	t->40	
 stra	f->38	m->1	n->1	t->48	x->2	
 stri	d->18	k->20	n->1	
 stru	k->120	n->4	
 stry	k->7	p->1	
 strä	c->3	n->19	v->15	
 strå	e->1	l->3	
 strö	k->1	m->8	
 stud	e->5	i->8	
 stug	o->1	
 stum	 ->1	
 stun	d->10	
 styc	k->2	
 stym	p->2	
 styr	 ->1	a->7	e->12	k->10	n->2	s->2	
 städ	a->2	e->10	
 stäl	l->172	
 stäm	d->1	m->14	n->1	p->1	
 stän	d->18	g->2	
 stär	k->22	
 stäv	 ->1	j->1	
 stå 	a->1	e->1	f->11	i->5	k->4	t->1	u->2	
 ståe	n->3	
 stål	f->5	g->1	i->25	s->4	v->5	
 stån	d->117	
 står	 ->94	,->1	
 ståt	t->4	
 stöd	 ->142	,->8	.->32	?->1	d->2	e->105	j->67	m->2	n->1	p->1	r->2	s->11	å->5	
 stöl	d->1	
 stör	 ->1	n->4	r->73	s->36	
 stöt	a->2	e->2	f->1	t->12	
 subj	e->1	
 subs	i->23	t->4	
 subv	e->10	
 succ	e->5	
 sudd	a->1	
 summ	a->3	o->7	
 sund	 ->1	a->4	
 supr	a->1	
 susp	e->1	
 sutt	i->1	
 suve	r->17	
 svag	 ->2	a->7	h->12	
 svan	s->1	
 svar	 ->27	,->2	.->6	a->23	e->12	s->2	t->2	
 svek	 ->2	
 sven	s->2	
 svep	s->1	t->1	
 sväl	t->2	
 svåg	e->1	
 svån	g->1	
 svår	 ->5	a->23	b->2	i->30	l->2	t->28	ö->1	
 syde	u->1	
 sydk	u->1	
 sydv	ä->1	
 sydö	s->1	
 syft	a->31	e->37	
 symb	o->9	
 symp	a->8	t->1	
 syn 	a->1	i->1	p->4	
 syna	 ->1	s->3	
 synd	 ->4	a->2	e->1	r->1	
 syne	n->1	r->2	s->1	
 synl	i->7	
 synn	e->51	
 syno	n->1	
 synp	u->21	
 syns	 ->1	ä->4	
 synt	e->1	
 synv	i->12	
 syri	e->4	s->4	
 syss	e->102	l->6	
 syst	e->114	
 säg:	 ->1	
 säga	 ->147	,->15	.->2	:->4	s->5	
 säge	r->73	
 sägs	 ->5	
 säke	r->224	
 säkr	a->19	
 sälj	a->3	
 säll	a->2	s->3	
 sämr	e->5	
 säms	t->5	
 sänd	a->4	e->9	n->1	
 sänk	a->5	n->1	
 sära	r->1	
 särb	e->1	
 särk	i->1	
 särs	k->156	
 säso	n->1	
 säte	.->1	
 sätt	 ->169	,->24	.->45	:->1	?->2	a->28	e->36	s->3	
 så a	l->3	m->1	n->1	t->127	v->1	
 så b	a->1	e->3	l->4	o->1	r->3	y->1	
 så d	e->6	r->2	
 så e	f->3	n->1	
 så f	a->3	i->4	o->3	r->1	å->3	ö->4	
 så g	r->3	ö->1	
 så h	a->2	e->2	j->4	o->2	ä->3	ö->1	
 så i	l->1	m->1	n->5	
 så j	a->1	
 så k	a->15	o->7	r->3	u->1	ä->1	
 så l	i->4	ä->15	å->12	
 så m	a->1	y->33	å->18	
 så n	o->1	ä->2	ö->2	
 så o	f->4	g->1	m->1	
 så p	a->2	å->1	
 så r	i->2	ä->1	
 så s	a->1	e->1	k->8	m->6	n->27	o->19	t->10	v->3	ä->18	
 så t	i->3	r->3	
 så u	p->3	t->2	
 så v	e->1	i->24	ä->3	
 så ä	r->16	
 så ö	p->1	
 så, 	a->2	i->1	n->1	s->1	t->1	
 så. 	D->1	
 så.D	e->1	
 så.I	 ->1	
 så.O	c->1	
 så: 	a->1	
 såda	n->163	
 såg 	i->1	n->1	s->1	u->2	Ö->1	
 sågv	e->1	
 såhä	r->1	
 såle	d->40	
 sålu	n->4	
 sång	 ->1	e->2	
 sårb	a->2	
 såso	m->31	
 såti	l->1	
 såvi	d->3	
 såvä	l->40	
 södr	a->6	
 söka	 ->3	s->1	
 söke	r->5	
 sönd	e->7	
 söne	r->1	
 sörj	a->7	d->1	e->2	
 t.ex	.->19	
 t.o.	m->7	
 ta A	m->1	
 ta a	n->3	t->1	v->2	
 ta b	o->2	
 ta d	e->21	
 ta e	m->4	n->4	t->5	
 ta f	o->1	r->7	u->1	
 ta g	e->1	
 ta h	a->7	e->1	j->1	ä->27	
 ta i	 ->1	n->2	s->1	t->14	
 ta l	ä->3	å->1	
 ta m	e->3	i->3	å->1	
 ta n	y->1	
 ta o	c->1	m->1	s->3	
 ta p	å->2	
 ta r	e->2	
 ta s	i->9	k->1	t->8	
 ta t	i->8	v->1	
 ta u	p->58	t->1	
 ta v	e->1	ä->1	å->1	
 ta ö	v->3	
 ta.J	a->1	
 ta?D	e->1	
 tabu	 ->1	
 tack	 ->27	,->1	.->2	a->104	l->1	o->1	s->8	
 tag 	i->2	s->2	
 tage	t->14	
 tagi	t->58	
 tagn	a->1	
 tak 	f->1	
 tak,	 ->1	
 take	t->1	
 takt	 ->4	i->3	
 tal 	h->1	i->2	o->3	
 tal,	 ->1	
 tal.	H->1	K->1	V->1	
 tala	 ->48	d->17	n->3	r->80	s->5	t->15	
 tale	n->1	s->4	t->2	
 talm	a->418	
 talr	i->4	
 tals	.->1	
 tank	-->1	a->11	e->62	f->6	r->2	
 tapp	a->3	
 tar 	a->3	d->3	e->4	f->5	g->1	h->3	i->10	k->1	l->1	m->2	n->2	p->4	r->1	s->3	t->4	u->10	v->5	ö->2	
 tarv	l->1	
 tas 	b->3	d->1	f->2	i->5	k->1	m->2	n->1	o->3	p->1	u->13	
 task	 ->1	
 tax-	f->3	
 taxe	r->1	
 teat	e->1	
 teck	e->9	n->2	
 tekn	i->45	
 tele	f->1	k->3	n->1	v->1	
 tema	,->1	t->1	
 temp	e->4	o->2	
 tend	e->12	
 teor	e->2	
 tera	t->2	
 term	e->3	
 terr	i->17	o->10	
 text	 ->9	,->5	.->1	e->20	
 the 	R->1	c->1	i->1	
 tibe	t->9	
 tid 	a->6	b->1	c->1	d->6	e->1	f->5	g->1	h->3	i->1	k->2	l->1	o->1	p->3	s->6	t->2	v->2	ä->2	å->2	
 tid,	 ->7	
 tid.	D->3	F->1	K->1	S->1	T->1	
 tide	n->48	r->3	
 tidi	g->85	
 tidn	i->4	
 tidp	u->10	
 tids	b->1	f->10	g->1	i->1	m->2	p->9	r->7	s->1	å->3	ö->1	
 tidt	a->6	
 tige	r->2	
 tigg	e->1	
 till	 ->1735	!->1	,->17	.->14	:->1	?->3	b->55	d->12	e->3	f->107	g->47	h->50	k->15	m->5	n->6	r->65	s->69	t->11	v->89	ä->192	å->42	
 timm	a->6	e->3	
 ting	 ->3	
 tio 	f->1	g->2	m->2	ä->1	å->4	
 tiot	a->5	u->1	
 tisd	a->2	
 tite	l->1	
 titt	 ->2	a->20	
 tjat	a->1	
 tjoc	k->2	
 tjug	o->4	
 tjän	a->8	s->110	
 tjär	a->1	
 toba	k->2	
 tog 	d->2	e->1	h->2	i->1	l->1	m->1	n->1	o->1	r->1	s->1	u->9	
 togs	 ->8	
 tole	r->14	
 tolk	a->10	n->14	
 tolv	 ->1	
 tom 	r->1	
 tomm	a->1	
 tomr	u->2	
 ton 	5->1	a->2	f->3	i->2	k->1	o->2	s->1	t->1	å->1	
 ton,	 ->1	
 ton/	å->2	
 tong	i->1	
 tonv	i->4	
 tonå	r->1	
 topp	e->3	m->9	
 tord	e->1	
 tork	a->1	
 torn	e->1	
 torp	e->2	
 tors	d->8	
 tort	e->1	y->1	
 torv	e->4	
 tota	l->34	
 toxi	s->1	
 trad	i->18	
 traf	i->7	
 trag	e->4	i->6	
 trak	a->1	
 tram	p->1	
 tran	s->107	
 tras	a->1	m->1	s->1	
 trau	m->1	
 trav	a->1	e->1	
 tre 	a->4	b->1	d->1	f->7	g->3	i->1	k->4	m->15	o->6	p->2	r->1	s->8	t->1	v->5	å->3	ö->1	
 tre,	 ->2	
 tre:	 ->1	
 tred	j->72	
 trek	l->1	
 trem	å->1	
 tren	d->1	
 tret	t->5	
 trev	l->3	
 tril	j->1	
 trio	 ->1	
 tro 	a->4	d->1	m->1	n->2	p->2	ä->1	
 tro.	V->1	
 trod	d->3	
 trog	e->1	
 troj	k->1	
 trol	i->9	
 tron	 ->1	
 tror	 ->150	,->1	
 trot	s->46	t->2	
 trov	ä->14	
 trup	p->2	
 trus	t->3	
 tryc	k->6	
 tryg	g->6	
 trä 	u->1	ö->1	
 träd	 ->4	,->1	.->1	a->6	d->6	e->5	
 träf	f->9	
 trän	g->2	i->1	
 träp	r->1	
 träs	k->1	
 trät	o->1	t->6	
 tråd	a->3	e->1	
 tråk	i->3	
 trån	g->1	
 trög	h->1	
 trös	k->3	t->1	
 tröt	t->1	
 tuff	 ->1	a->1	
 tull	f->1	g->1	
 tumm	a->3	
 tunc	 ->1	
 tung	 ->6	a->2	m->6	r->1	t->2	
 tunn	e->2	l->2	
 tur 	b->1	d->2	k->1	v->1	ä->1	
 tur,	 ->1	
 tur.	N->1	
 ture	r->1	
 turi	s->22	
 turk	a->2	i->6	
 tuse	n->9	
 tvek	a->23	l->1	s->5	
 tvet	y->5	
 tvin	g->25	
 tvis	t->6	
 tviv	e->32	l->6	
 tvun	g->11	
 tvär	p->2	s->1	t->14	
 tvät	t->1	
 två 	a->10	b->3	d->2	e->7	f->23	g->2	h->2	i->3	j->1	k->4	l->2	m->8	n->2	o->2	p->12	r->2	s->12	t->8	u->3	v->5	y->1	å->8	
 två.	B->1	
 två:	 ->2	
 tvåh	u->1	
 tvån	g->6	
 ty E	u->1	
 ty d	e->4	
 ty i	 ->1	
 ty n	a->1	ä->1	
 ty p	å->2	
 ty v	i->2	
 tyck	a->3	e->59	s->8	t->7	
 tyde	r->6	
 tydl	i->104	
 tyge	l->1	
 tyna	n->1	
 tyng	a->1	d->6	e->1	s->2	
 typ 	C->1	a->18	f->1	
 typ,	 ->1	
 typ.	D->1	E->1	
 type	n->12	r->4	
 typf	a->1	
 typg	o->1	
 tysk	a->20	t->2	
 tyst	 ->3	
 tyvä	r->29	
 täck	a->2	e->8	s->4	
 täml	i->3	
 tänd	a->1	
 tänk	 ->1	a->28	b->2	e->34	t->8	
 täpp	a->3	e->1	
 tärt	 ->1	
 täta	,->1	r->1	
 täte	n->2	
 tävl	a->2	i->1	
 tåg 	e->1	
 tåg,	 ->1	
 tåge	t->1	
 tågk	r->1	
 tågo	l->1	
 tål 	a->1	
 tåla	m->2	
 tömm	e->1	
 u-lä	n->1	
 ulti	m->1	
 ultr	a->2	
 umgä	n->1	
 unda	n->52	
 unde	r->473	
 undg	å->1	
 undr	a->11	
 undv	i->35	
 ung 	m->1	
 unga	 ->5	,->1	
 ungd	o->14	
 unge	f->8	
 unik	a->1	t->1	
 unil	a->2	
 unio	n->432	
 univ	e->4	
 upp 	-->1	E->1	T->1	a->11	b->2	d->41	e->20	f->14	g->3	h->5	i->22	k->2	l->3	m->8	n->4	o->7	p->9	r->4	s->10	t->13	u->5	v->3	ä->7	
 upp,	 ->11	
 upp.	A->1	D->4	J->7	P->1	V->2	Ä->2	
 uppb	a->1	r->3	y->7	ä->1	å->1	
 uppd	a->2	e->3	r->21	
 uppe	h->12	n->35	
 uppf	a->50	y->54	ö->22	
 uppg	i->75	r->1	å->8	ö->1	
 upph	e->1	o->13	ä->5	ö->10	
 uppk	o->6	
 uppl	e->17	y->4	ö->3	
 uppm	a->58	j->2	u->21	ä->55	
 uppn	å->93	
 uppr	e->53	i->6	o->1	u->1	y->1	ä->30	ö->5	
 upps	a->7	k->28	p->2	t->36	ä->3	
 uppt	a->2	r->10	ä->10	
 uppv	i->5	ä->2	
 ur E	U->1	u->1	
 ur U	C->1	
 ur b	i->1	r->1	u->1	y->1	
 ur d	e->4	
 ur e	k->2	n->6	r->1	t->3	
 ur i	n->1	
 ur j	o->1	
 ur k	o->1	u->1	
 ur m	a->1	i->5	y->1	å->1	
 ur p	e->1	o->1	
 ur s	i->1	t->1	ö->1	
 ur t	e->1	
 ur v	i->1	
 uran	 ->3	.->1	?->1	i->2	v->4	
 urba	n->1	
 urho	l->4	
 urmi	n->1	
 ursk	i->3	u->1	
 ursp	r->19	å->1	
 ursä	k->14	
 urva	l->5	t->8	
 ut 1	0->1	
 ut T	o->1	
 ut a	c->1	m->1	n->1	t->3	v->1	
 ut b	e->1	
 ut d	e->7	
 ut e	n->3	t->2	x->1	
 ut f	r->4	ö->4	
 ut g	e->1	
 ut h	a->2	ö->1	
 ut i	 ->3	n->1	
 ut k	o->1	u->1	
 ut m	e->3	i->2	o->2	y->1	
 ut n	a->1	å->1	
 ut o	c->4	s->1	
 ut p	e->2	o->1	r->2	å->14	
 ut r	e->2	
 ut s	i->2	o->2	t->1	y->1	å->2	
 ut t	i->3	
 ut u	n->1	p->1	
 ut ö	v->5	
 ut, 	a->3	b->1	e->1	f->1	h->1	m->4	n->1	o->2	s->2	t->1	u->2	å->1	
 ut. 	D->1	
 ut.D	e->4	å->1	
 ut.F	i->1	ö->2	
 ut.G	r->1	
 ut.J	a->4	
 ut.K	r->1	
 ut.S	t->1	
 ut.V	i->1	
 ut.Ä	v->1	
 ut: 	f->1	
 ut?.	 ->1	
 ut?E	t->1	
 utan	 ->286	,->1	f->32	
 utar	b->31	m->10	
 utba	s->1	
 utbe	t->5	
 utbi	l->45	
 utbr	e->4	
 utbu	d->4	
 utby	g->3	t->11	
 utde	l->1	
 ute 	e->1	p->1	t->1	u->1	
 utel	ä->3	
 utes	l->19	t->4	
 utfa	l->1	s->3	
 utfl	a->1	y->1	
 utfo	r->39	
 utfr	å->7	
 utfä	r->12	s->1	
 utfö	r->37	
 utga	v->1	
 utgi	c->1	f->13	v->2	
 utgj	o->4	
 utgå	 ->4	n->16	r->8	v->1	
 utgö	r->59	
 uthä	r->2	
 utif	r->16	
 utjä	m->5	
 utka	n->1	s->15	
 utko	m->2	n->1	
 utkr	ä->3	
 utla	n->5	
 utlo	v->3	
 utlä	g->1	m->2	n->4	
 utlå	t->2	
 utlö	s->2	
 utma	n->20	
 utmy	n->1	
 utmä	r->32	
 utny	t->40	
 utnä	m->4	
 utom	 ->4	e->3	o->7	s->2	
 utpe	k->1	
 utpl	å->2	
 utpr	e->1	ä->1	
 utre	d->8	
 utri	k->19	
 utro	p->2	t->3	
 utru	s->3	
 utry	m->7	
 uträ	t->2	
 utsa	t->6	
 utse	 ->3	d->1	e->1	r->1	s->2	t->1	
 utsi	k->1	
 utsk	o->126	
 utsl	a->14	ä->6	
 utst	a->10	r->28	ä->2	å->1	ö->1	
 utsu	g->1	
 utsä	t->7	
 utså	g->3	
 utta	l->98	
 uttj	ä->24	
 utto	l->1	r->1	
 uttr	y->71	ä->1	
 uttö	m->5	
 utva	l->1	
 utve	c->225	r->3	
 utvi	d->103	s->1	
 utvä	r->31	
 utök	a->11	n->1	
 utöv	a->15	e->13	
 vack	e->2	l->1	r->6	
 vad 	B->1	E->1	G->1	K->2	S->1	a->1	b->14	d->30	e->3	f->3	g->47	h->4	i->1	j->7	k->8	m->9	n->5	o->3	p->1	r->2	s->60	t->1	v->27	ä->6	
 vad?	D->1	
 vaga	 ->2	
 vagn	e->1	
 vagt	.->1	
 vaka	 ->1	r->1	
 vaks	a->9	
 vakt	 ->1	
 vaku	u->2	
 val 	a->4	d->1	g->1	i->1	s->2	u->1	ä->1	å->1	
 val,	 ->2	
 val.	D->1	I->1	M->1	V->1	
 val;	 ->1	
 valb	a->1	
 vald	 ->3	a->11	e->8	i->1	
 vale	n->3	t->4	
 valf	r->5	
 valk	r->4	
 vall	f->1	
 valr	e->1	
 valt	 ->5	,->1	a->1	i->1	s->4	
 valu	t->22	
 van 	D->2	H->20	V->1	d->9	
 vana	 ->1	
 vanh	e->2	
 vanl	i->11	
 vano	r->1	
 vans	k->1	
 vape	n->13	
 vapn	e->2	
 var 	1->5	9->1	K->1	W->1	a->18	b->12	d->33	e->28	f->12	g->1	h->4	i->13	j->3	k->4	l->6	m->15	n->9	o->9	p->2	r->3	s->13	t->6	u->3	v->9	ä->2	ö->4	
 var,	 ->1	
 var.	D->1	
 vara	 ->342	"->1	,->1	.->2	:->1	d->1	k->4	n->12	v->4	
 vard	a->4	e->1	
 vare	 ->18	f->1	n->2	
 varf	ö->39	
 varg	a->1	
 vari	 ->1	e->2	t->71	
 varj	e->83	
 vark	e->14	
 varm	a->3	t->12	
 varn	a->7	i->5	
 varo	r->1	
 vars	 ->28	a->1	
 vart	 ->4	a->3	e->1	
 varv	i->3	s->3	
 vatt	e->23	n->3	
 veck	a->23	o->17	
 vede	r->13	
 vekh	e->4	
 vela	t->7	
 vem 	b->1	f->1	i->1	s->13	ä->1	
 vems	 ->1	
 vent	i->1	
 verb	a->1	
 veri	f->1	
 verk	.->1	a->51	e->31	l->183	n->1	s->62	t->8	
 vers	i->11	
 vert	i->3	
 vet 	a->36	b->1	f->3	g->1	h->3	i->9	j->3	k->3	m->2	n->4	o->3	r->1	s->2	t->1	v->10	ä->3	
 vet,	 ->11	
 veta	 ->27	,->1	
 vete	n->69	r->12	
 vett	i->3	v->1	
 vi -	 ->3	
 vi 1	9->1	
 vi 5	5->1	
 vi E	u->2	
 vi L	i->1	
 vi P	r->1	
 vi a	)->1	b->3	c->1	g->2	l->37	n->30	r->6	t->41	v->7	
 vi b	a->5	e->54	i->3	l->6	o->10	r->2	y->1	ö->27	
 vi d	a->1	e->26	i->15	o->1	r->1	ä->6	å->6	
 vi e	f->5	g->3	k->1	m->5	n->14	r->3	t->9	u->2	v->1	x->1	
 vi f	a->14	i->2	o->13	r->6	u->3	å->18	ö->41	
 vi g	a->1	e->15	i->1	j->4	l->4	o->4	r->2	ä->2	ö->19	
 vi h	a->135	e->7	i->5	j->1	o->4	ä->14	å->7	ö->2	
 vi i	 ->56	a->1	b->2	g->1	n->134	
 vi j	u->11	
 vi k	a->65	l->2	n->1	o->41	r->4	u->7	v->1	ä->2	
 vi l	a->3	i->7	o->1	y->5	ä->9	å->2	
 vi m	e->20	i->3	o->3	y->1	å->63	
 vi n	a->4	u->21	y->2	ä->6	å->2	
 vi o	b->1	c->31	f->2	m->1	s->9	
 vi p	l->2	r->1	å->12	
 vi r	e->13	i->2	o->1	u->2	ä->2	å->1	ö->7	
 vi s	a->6	e->17	j->4	k->68	l->3	n->8	o->16	p->2	t->24	v->1	y->2	ä->6	å->4	
 vi t	.->1	a->24	e->1	i->15	o->1	r->8	v->1	y->7	ä->4	
 vi u	n->7	p->17	r->1	t->13	
 vi v	a->9	e->22	i->34	ä->6	å->3	
 vi y	t->1	
 vi ä	g->4	n->10	r->28	v->5	
 vi å	l->1	r->1	s->1	t->4	
 vi ö	n->5	v->3	
 vi, 	g->1	j->3	k->1	l->1	m->1	n->1	s->5	t->1	ä->2	
 vi.V	i->1	
 vi?.	H->1	
 via 	B->1	E->1	R->1	a->1	b->1	d->1	e->1	k->1	o->1	s->1	t->1	u->1	
 vice	 ->13	
 vid 	1->1	7->1	B->1	E->6	G->1	H->1	K->1	M->1	P->1	a->13	b->7	d->34	e->15	f->21	g->3	h->5	i->1	j->2	k->7	l->1	m->3	n->5	o->7	p->8	r->5	s->15	t->12	u->14	v->8	å->2	ö->2	
 vid,	 ->2	
 vid.	H->1	J->1	
 vida	 ->2	r->37	
 vidd	 ->1	e->1	
 vidg	a->2	
 vidh	å->4	ö->1	
 vidm	a->1	
 vids	t->1	
 vidt	a->62	o->2	
 vift	a->1	
 vigv	a->1	
 vigö	r->1	
 vikt	 ->11	,->2	.->2	e->9	i->328	
 vila	r->2	
 vild	a->1	
 vilj	a->175	e->2	
 vilk	a->90	e->227	
 vill	 ->529	,->8	.->2	e->10	i->4	k->38	o->1	
 vils	e->3	
 vilt	,->1	
 vin 	E->1	
 vind	 ->1	f->4	
 vinn	a->4	e->2	
 vins	t->11	
 virk	e->3	
 virr	v->1	
 vis 	a->1	d->2	f->1	h->1	i->1	m->1	o->2	s->1	u->1	
 vis,	 ->2	
 vis.	D->1	
 visa	 ->29	d->7	r->55	s->2	t->29	v->1	
 visd	o->1	
 vise	r->2	t->5	
 visi	o->2	
 visk	a->1	
 viss	 ->35	a->128	e->11	h->3	t->10	
 vist	a->4	e->1	
 visu	a->1	e->1	m->1	
 vitb	o->50	
 vitt	 ->1	n->4	
 volu	n->4	
 voly	m->3	
 von 	B->1	E->1	W->16	
 vore	 ->29	
 vote	r->3	
 votu	m->1	
 vrak	 ->3	,->1	
 vred	g->1	
 vrid	e->1	
 vräk	t->1	
 vunn	e->1	i->2	
 vuxi	t->1	
 vuxn	a->2	
 väck	a->4	e->5	s->1	t->7	
 väde	r->1	
 vädj	a->9	
 väg 	[->1	a->6	b->1	g->2	h->1	i->1	m->2	t->1	ä->1	å->1	
 väg,	 ->9	
 väg.	B->1	D->1	E->1	J->1	M->1	
 vägN	ä->1	
 väga	 ->1	r->11	
 vägb	y->1	
 väge	n->16	r->3	
 vägl	e->5	
 vägm	ä->1	
 vägn	a->16	
 vägr	a->19	ö->1	
 vägs	k->2	
 väkt	a->2	
 väl 	a->6	b->2	d->2	e->1	f->5	g->2	h->3	i->3	k->4	l->1	m->5	o->2	p->1	r->3	s->2	t->3	u->4	v->2	ä->3	ö->1	
 väl,	 ->2	
 väl.	J->1	M->1	S->1	
 välb	e->1	
 väld	i->20	
 välf	u->1	ä->8	
 välg	r->2	ö->1	
 välj	a->17	e->5	
 välk	l->1	o->49	ä->3	
 väll	e->1	
 välm	e->2	å->2	
 väls	i->1	t->7	
 vält	a->2	
 välu	t->3	
 vän 	o->1	
 vänd	a->6	e->9	p->5	
 vänl	i->4	
 vänn	e->2	
 väns	k->1	t->15	
 vänt	 ->1	a->44	
 väpn	a->2	
 värd	 ->4	a->2	e->60	i->4	
 värl	d->50	
 värn	a->3	
 värr	e->2	
 värs	t->8	
 värt	 ->4	
 väse	n->29	
 väst	k->1	v->1	
 vävn	a->3	
 vävt	 ->1	
 växa	 ->1	.->2	n->6	
 växe	l->3	r->7	
 växl	a->1	i->2	
 växt	e->2	h->7	s->3	
 våg 	a->1	
 våga	r->5	t->1	
 våge	n->1	
 vågl	ä->1	
 våld	 ->2	e->2	s->6	t->2	
 våll	a->1	
 våni	n->2	
 vår 	a->1	b->8	d->12	e->3	f->12	g->15	i->4	k->7	l->6	m->10	n->1	o->2	p->8	r->10	s->17	t->4	u->9	v->5	å->4	ö->1	
 vår,	 ->1	
 våra	 ->150	
 vård	s->2	
 vårt	 ->105	,->1	
 vörd	n->1	
 wale	s->1	
 webb	p->1	
 wors	t->1	
 yngr	e->1	
 yngs	t->1	
 yppa	s->1	
 yppe	r->1	
 yrka	 ->1	r->1	
 yrke	n->3	s->15	
 yta.	I->1	
 ytli	g->2	
 ytte	r->89	
 yttr	a->39	e->3	
 zige	n->4	
 zon 	3->1	V->1	
 zone	r->1	
 zoni	n->1	
 º C.	 ->1	
 Ämna	r->1	
 Ändå	 ->1	
 Ännu	 ->2	
 Är k	o->1	
 Ärad	e->2	
 Även	 ->11	
 Å PS	E->1	
 Å ko	m->1	
 Å so	c->1	
 Årli	g->1	
 Åtgä	r->3	
 Île-	d->1	
 ÖVP 	(->1	a->2	m->1	
 Öppe	n->1	
 Öste	r->75	u->5	
 Östt	y->2	
 äckl	a->1	
 äga 	r->18	
 ägan	d->3	
 ägar	a->1	e->12	n->2	
 ägde	 ->1	
 äger	 ->5	
 ägg"	 ->1	
 ägna	 ->9	r->13	s->2	t->4	
 ägt 	r->9	
 äkte	n->1	
 äldr	e->7	
 älsk	a->2	
 ämbe	t->7	
 ämna	d->2	r->2	
 ämne	 ->3	.->2	:->1	n->15	t->4	
 än 1	 ->2	0->3	6->1	
 än 2	0->1	1->1	
 än 3	0->2	
 än E	u->1	
 än F	o->1	
 än W	a->1	
 än a	l->2	t->12	v->1	
 än b	a->2	
 än d	e->18	i->2	
 än e	j->1	n->29	t->3	
 än f	a->2	e->2	ö->5	
 än g	e->1	
 än h	a->2	i->1	
 än i	 ->10	n->2	
 än j	a->1	
 än k	a->2	o->4	
 än l	i->1	o->1	ä->1	
 än m	a->4	e->2	i->5	å->1	
 än n	ä->1	å->6	
 än o	c->1	m->1	
 än p	.->1	e->1	å->2	
 än r	e->4	
 än s	a->1	o->1	t->2	ä->1	å->5	
 än t	i->3	r->2	v->2	
 än v	a->7	i->7	ä->3	å->1	
 än ä	r->4	
 än, 	m->1	
 än.J	a->1	
 ända	 ->7	,->1	m->12	
 ändl	ö->1	
 ändp	u->1	
 ändr	a->48	i->240	
 ändå	 ->51	,->1	.->1	
 ängs	l->1	
 ännu	 ->72	.->4	;->1	
 äntl	i->20	
 är "	k->1	
 är -	 ->4	
 är 1	0->1	
 är 2	5->1	
 är 3	0->1	
 är E	U->3	g->1	u->8	
 är F	N->1	
 är P	o->2	
 är W	a->1	
 är a	b->10	c->2	k->4	l->30	m->1	n->29	r->1	t->117	v->37	
 är b	a->11	e->65	o->3	r->20	y->1	ä->6	å->4	
 är c	e->2	
 är d	a->7	e->290	i->2	j->4	o->17	r->1	ä->29	å->5	ö->1	
 är e	f->4	g->6	k->1	m->11	n->216	t->116	u->1	v->1	x->4	
 är f	a->20	e->6	i->2	l->3	o->15	r->26	u->11	y->1	å->1	ö->76	
 är g	a->7	e->7	i->1	j->2	l->13	o->8	r->7	
 är h	a->1	e->32	i->1	j->1	o->4	u->6	ä->4	å->1	ö->1	
 är i	 ->39	b->2	d->1	l->1	n->132	s->1	
 är j	a->26	u->18	ä->1	
 är k	a->4	l->14	n->5	o->35	r->2	v->1	ä->7	
 är l	a->4	e->5	i->19	o->1	y->1	ä->15	å->4	ö->4	
 är m	a->1	e->44	i->12	o->2	u->1	y->55	å->4	ö->21	
 är n	a->16	e->2	i->2	o->2	u->11	y->4	ä->10	å->25	ö->33	
 är o	a->5	b->4	c->38	e->8	f->10	j->1	k->2	l->2	m->8	n->1	r->6	s->2	t->3	u->3	
 är p	a->4	e->1	l->2	o->8	r->15	å->11	
 är r	e->21	i->10	o->2	u->2	ä->12	å->2	
 är s	a->10	e->2	i->1	j->8	k->15	l->1	o->7	p->5	t->16	u->2	v->10	y->7	ä->44	å->25	
 är t	a->1	e->3	i->34	o->2	r->5	v->7	y->10	ä->2	
 är u	n->7	p->20	r->1	t->21	
 är v	a->12	e->9	i->72	u->1	ä->27	å->10	
 är y	r->1	t->9	
 är ä	l->2	n->11	r->1	v->2	
 är å	t->2	
 är ö	d->1	n->2	p->3	v->25	
 är, 	a->1	f->2	h->1	i->1	k->1	m->3	o->2	s->1	t->1	
 är..	 ->1	
 är.D	e->2	
 är.E	n->1	
 är.F	ö->1	
 är.H	e->1	
 är.J	a->2	
 är.k	o->1	
 är: 	F->1	h->1	n->1	v->1	Ä->1	
 är?H	a->1	
 ärad	e->22	
 äran	 ->4	
 ären	d->18	
 ärli	g->8	
 äro 	t->1	
 äter	 ->1	
 även	 ->266	t->9	
 å PP	E->1	
 å an	d->7	
 å de	n->3	
 å en	a->11	
 å mi	n->2	
 å re	g->1	
 å ut	s->1	
 åber	o->1	
 åhör	a->1	
 åkla	g->37	
 åkte	 ->1	
 ålag	d->1	t->2	
 ålde	r->9	
 ålig	g->5	
 åläg	g->5	
 ånyo	 ->1	
 år -	 ->1	
 år 1	9->19	
 år 2	0->33	
 år a	n->2	t->4	v->1	
 år b	o->1	
 år d	ä->1	å->1	
 år e	f->4	l->2	
 år f	r->4	ö->4	
 år h	a->2	
 år i	 ->3	n->1	
 år k	o->2	r->1	
 år l	e->1	
 år n	u->1	
 år o	c->6	m->1	
 år p	å->2	
 år s	e->15	k->3	o->8	
 år t	i->3	
 år u	n->1	t->1	
 år v	i->1	
 år ä	g->1	r->1	
 år å	t->1	
 år, 	d->1	e->1	f->1	k->1	m->4	n->1	o->3	t->1	u->3	v->1	ä->1	
 år.D	e->9	
 år.E	n->1	
 år.F	ö->2	
 år.H	u->1	ä->1	
 år.I	 ->1	
 år.J	a->2	
 år.K	ä->1	
 år.L	y->1	
 år.O	m->1	
 år.R	e->1	
 år.S	a->1	
 år.T	y->1	
 år.V	e->1	i->2	
 år.Ä	n->1	
 årat	a->1	
 åren	 ->26	,->5	.->6	s->2	
 året	 ->18	,->6	.->3	s->4	
 århu	n->7	
 årli	g->8	
 års 	E->1	b->3	e->1	p->1	s->1	t->3	ö->1	
 årsb	e->2	
 årsr	a->2	
 årst	i->1	
 årta	l->1	
 årti	o->1	
 årtu	s->3	
 åsam	k->3	
 åsat	t->1	
 åsik	t->50	
 åskå	d->2	
 åsta	d->25	
 åsyf	t->5	
 åt E	u->1	
 åt F	ö->1	
 åt a	n->1	t->7	
 åt b	e->1	
 åt d	e->27	
 åt e	g->1	n->3	t->2	
 åt f	o->1	r->1	
 åt g	e->1	
 åt h	u->1	
 åt i	 ->1	m->1	n->1	
 åt j	ä->1	
 åt k	o->3	v->1	
 åt l	i->1	
 åt m	a->1	
 åt n	u->1	y->1	
 åt p	a->1	
 åt r	e->1	ä->3	
 åt s	a->1	i->4	y->1	
 åt t	i->1	v->1	ä->1	
 åt u	n->1	
 åt Ö	s->1	
 åt ä	m->1	r->2	
 åt å	t->1	
 åt, 	k->1	u->1	
 åt.K	o->1	
 åt.N	ä->1	
 åta 	s->3	
 åtag	a->28	i->2	
 åtal	 ->5	.->1	a->5	s->7	
 åtan	k->1	
 åtar	 ->2	
 åter	 ->21	a->18	b->1	e->1	f->12	g->7	h->4	i->25	k->8	l->2	n->10	s->33	t->9	u->32	v->67	
 åtfö	l->12	
 åtgä	r->218	
 åtmi	n->27	
 åtnj	u->1	
 åtsk	i->3	
 åtst	r->2	
 åtta	 ->4	,->1	
 åtto	n->1	
 åvil	a->1	
 öar 	s->1	
 öarn	a->5	
 öbo 	v->1	
 öde 	i->1	
 öde,	 ->4	
 öde.	D->1	
 öde?	H->1	
 ödel	a->1	
 ödem	a->1	
 ödes	b->1	d->2	g->1	
 ögat	.->1	
 ögon	 ->5	,->1	b->13	
 öka 	a->6	b->1	d->2	f->2	i->1	j->1	k->7	m->2	s->6	v->1	
 öka.	O->1	R->1	T->1	
 ökad	 ->27	e->9	
 ökan	d->3	
 ökar	 ->12	,->3	.->1	
 ökas	 ->2	,->1	
 ökat	 ->15	.->1	
 ökni	n->18	
 öl o	c->1	
 öm t	a->1	
 ömma	 ->1	
 ömse	s->5	
 ömtå	l->1	
 ön N	o->1	
 önsk	a->48	e->3	n->2	v->10	
 öppe	n->64	t->14	
 öppn	a->16	i->4	
 öre 	m->1	
 öreg	i->7	
 öron	,->1	m->2	
 öst 	o->1	
 östb	l->1	
 öste	r->49	u->3	
 östl	ä->1	
 östr	a->2	
 östu	t->2	
 övat	 ->1	
 över	 ->200	,->3	.->8	a->9	b->9	c->1	d->14	e->71	f->23	g->40	h->4	i->1	k->6	l->34	m->1	n->4	o->1	p->1	r->4	s->46	t->53	v->69	
 övni	n->5	
 övri	g->65	
! 199	9->1	
! All	a->1	t->1	
! Att	 ->1	
! Av 	o->1	
! Avf	a->1	
! Avs	e->1	
! Ber	e->1	
! Bes	l->1	
! Bet	r->1	
! Bla	n->1	
! Cen	t->1	
! Dag	e->1	
! De 	k->1	o->1	s->1	
! Den	 ->6	n->4	
! Det	 ->36	t->3	
! Dir	e->1	
! Där	 ->1	
! Díe	z->1	
! EU 	u->1	
! Eft	e->4	
! End	a->1	
! Era	 ->1	
! Ert	 ->1	
! Ett	 ->1	
! Eur	o->7	
! Fra	m->1	
! Fru	 ->1	
! Frå	g->1	
! Får	 ->1	
! För	 ->6	s->10	
! Gen	e->1	
! Got	t->1	
! Gru	p->3	
! Her	r->1	
! Hit	t->1	
! I b	e->1	u->1	ö->1	
! I d	a->5	e->4	
! I e	g->3	
! I l	i->1	
! I m	o->1	
! I u	t->1	
! Ing	e->1	
! Int	e->1	
! Ja,	 ->1	
! Jag	 ->109	
! Jon	c->1	
! Jäm	f->1	
! Kar	t->1	
! Kom	m->4	
! Kon	k->1	
! Lik	s->2	
! Låt	 ->9	
! Man	 ->1	
! Med	 ->1	
! Min	 ->4	a->1	
! Ni 	b->1	h->2	s->1	v->1	
! Nu 	f->1	
! När	 ->7	
! Någ	o->1	
! Olj	e->1	
! Om 	n->1	o->1	
! PPE	-->1	
! Par	l->1	
! Pri	o->1	
! På 	d->2	
! Pås	t->1	
! Reg	e->1	
! Rot	h->1	
! Råd	e->2	
! Sch	r->1	
! Sed	a->3	
! Sku	l->1	
! Som	 ->7	
! Str	a->1	
! Tac	k->3	
! The	a->1	
! Til	l->7	
! Tor	r->1	
! Tro	t->1	
! Und	e->4	
! Upp	d->1	
! Urs	ä->1	
! Uts	k->2	
! Vad	 ->4	
! Var	j->1	
! Vi 	f->4	h->6	k->2	m->1	s->2	v->3	ä->2	
! Vid	 ->2	
! Vis	s->1	
! Vår	 ->2	t->1	
! Änn	u->1	
! Äve	n->9	
! Å P	S->1	
! Å k	o->1	
! Å s	o->1	
! Årl	i->1	
! Öst	e->1	
!".De	t->1	
!"Det	 ->1	
!"Jag	 ->1	
!"Om 	e->1	
!(Par	l->1	
!. (F	R->1	
!.(NL	)->1	
!.Her	r->1	
!Allt	s->2	
!Amst	e->1	
!Andr	a->1	
!Av d	e->1	
!De a	n->1	
!De f	ö->1	
!De s	e->1	
!Den 	a->1	r->1	
!Denn	a->1	
!Det 	d->1	f->3	s->2	ä->7	
!Dett	a->1	
!Därf	ö->1	
!Efte	r->2	
!En v	i->1	
!Erik	a->1	
!Euro	p->1	
!Fru 	k->1	t->2	
!För 	m->1	
!Före	d->1	
!Geno	m->1	
!Han 	n->1	
!Herr	 ->9	
!Här 	r->1	
!I de	t->1	
!Jag 	f->3	h->3	k->1	n->1	r->1	s->3	t->2	u->1	v->2	ä->1	
!Kult	u->1	
!Leda	m->1	
!Låt 	o->1	
!Med 	d->1	
!Men 	F->1	e->1	j->1	v->1	
!Min 	d->1	
!Mina	 ->1	
!Myck	e->1	
!Männ	i->1	
!Ni h	a->1	
!När 	j->1	v->2	
!Om n	i->1	
!Om v	i->1	
!Prec	i->1	
!Röst	a->1	
!Sann	i->1	
!Skal	l->1	
!Tack	 ->1	
!Till	 ->2	å->1	
!Tror	 ->1	
!Tvär	t->1	
!Unde	r->1	
!Vi b	e->1	
!Vi f	å->1	
!Vi h	a->1	
!Vi s	k->1	
!Vi ä	r->1	
!Även	 ->2	
" (se	 ->1	
" - e	n->1	
" ald	r->1	
" att	 ->1	
" av 	k->1	
" bil	e->1	
" etc	.->1	
" fra	m->1	
" för	 ->1	
" gem	e->1	
" gör	 ->1	
" har	 ->1	
" i A	m->1	
" med	 ->2	
" mås	t->2	
" och	 ->6	
" på 	r->1	
" ska	l->1	
" som	 ->8	
" til	l->2	
" var	 ->1	
" Ära	d->1	
" är 	m->1	
"!I d	e->1	
"), v	i->1	
", "s	e->1	
", al	l->1	
", be	s->1	
", de	 ->1	t->1	
", dv	s->1	
", dä	r->1	
", ef	t->1	
", fö	r->1	
", i 	d->1	
", me	n->1	
", oc	h->4	
", so	m->5	
", vi	l->3	
".. (	F->1	
".Bar	a->1	
".Båd	a->1	
".De 	f->1	s->1	
".Den	n->1	
".Des	s->1	
".Det	 ->4	t->2	
".En 	s->1	
".Eur	o->1	
".His	t->1	
".I n	ä->1	
".Jag	 ->4	
".Jus	t->1	
".Kan	 ->1	
".Kin	n->1	
".När	 ->1	
".Om 	m->1	
".Ord	 ->1	
".Råd	e->1	
".Vi 	f->1	
"; öv	e->1	
"Amst	e->1	
"Att 	i->1	
"Big 	b->1	
"Det 	b->1	s->2	ä->3	
"EU-k	o->1	
"Equa	l->1	
"Euro	d->1	p->1	
"I de	n->1	
"Ja E	r->1	
"Ja, 	d->1	
"Jag 	a->1	s->1	
"Kult	u->4	
"Kvin	n->3	
"Loth	a->1	
"Med 	d->1	
"Mind	r->1	
"Mist	e->1	
"Olje	b->1	
"Om d	u->1	
"Om e	n->1	
"Port	u->1	
"Tibe	t->2	
"Ty h	a->1	
"Urba	n->1	
"affä	r->1	
"aldr	i->2	
"allm	ä->1	
"angi	v->3	
"avgö	r->1	
"bank	"->1	
"coup	 ->1	
"den 	b->1	s->2	
"dett	a->1	
"die 	R->1	
"döda	"->1	
"egen	f->1	
"ekol	o->1	
"en e	n->1	
"en l	ö->1	
"en w	a->1	
"entr	e->1	
"euro	p->3	
"fort	s->1	
"för"	.->1	
"geme	n->1	
"gend	e->1	
"hell	r->1	
"hero	i->1	
"in s	o->1	
"indi	k->1	
"inle	d->1	
"irre	p->1	
"ja t	i->1	
"koll	e->2	
"kron	j->1	
"kult	u->1	
"länd	e->1	
"läs 	t->1	u->1	
"mell	a->1	
"natu	r->1	
"ne j	e->1	
"norm	a->1	
"någo	t->1	
"ober	o->1	
"orme	n->1	
"ovil	l->1	
"part	i->1	
"påpe	k->1	
"refu	s->1	
"rest	e->1	
"resu	l->3	
"rikt	l->1	
"se p	å->1	
"shal	l->1	
"skad	e->1	
"spec	i->1	
"svag	a->1	
"till	b->1	
"utve	c->1	
"utåt	"->1	
"valu	t->1	
"varj	e->1	
"åter	n->1	
"öppe	n->1	
"över	m->1	
'Vad 	ä->1	
'eau 	d->1	
("die	 ->1	
(1409	4->2	
(1997	)->1	
(1998	)->3	-->2	
(1999	)->7	
(5713	/->1	
(8095	/->2	
(9614	/->1	
(98)0	6->1	
(99)0	0->1	5->1	
(A5-0	0->27	1->9	
(Appl	å->5	
(Arbe	t->1	
(B5-0	0->4	
(Bene	l->1	
(Brys	s->2	
(C5-0	2->2	3->5	
(CEN)	 ->2	
(CERN	)->1	
(CNS)	)->9	
(COD)	)->12	]->1	
(COS)	]->2	
(DA) 	D->1	V->1	
(DE) 	H->1	J->1	Ä->1	
(EG, 	E->1	
(EIF)	,->1	
(EL) 	F->1	H->1	J->1	
(EN) 	D->2	F->6	H->4	I->3	J->7	K->1	L->2	M->1	S->1	T->4	U->1	V->2	
(ES) 	-->1	
(EU-f	ö->1	
(EUGF	J->2	
(FI) 	J->1	
(FIPO	L->1	
(FPÖ)	.->1	
(FR) 	"->1	D->4	E->1	F->1	H->1	I->2	J->4	N->3	T->1	
(FUF)	 ->1	
(Geno	m->1	
(H-00	0->1	
(H-07	7->1	8->6	9->5	
(H-08	0->4	1->3	2->1	
(Howi	t->1	
(ICES	)->1	
(IFOP	)->1	
(IMO)	.->1	
(IT) 	D->1	H->1	O->1	
(Ihål	l->1	
(Inte	r->1	
(KOM(	1->6	9->2	
(Kult	u->2	
(Livl	i->2	
(NL) 	A->1	H->3	
(PPE-	D->1	
(PT) 	E->1	F->1	H->9	J->2	L->1	N->1	V->1	
(Parl	a->16	
(Prot	o->1	
(SEK(	1->1	
(SPÖ)	 ->1	
(SYN)	)->1	
(Samm	a->4	
(Talm	a->8	
(Utsk	o->2	
(art.	 ->1	
(arti	k->6	
(att 	s->1	
(avsn	i->1	
(de n	y->1	
(det 	e->1	
(efte	r->1	
(elle	r->1	
(en i	n->1	
(en m	i->1	
(fisk	e->4	
(fort	s->1	
(före	d->3	
(häls	o->1	
(i de	t->1	
(i så	d->1	
(infö	r->1	
(inre	 ->1	
(kodi	f->2	
(komm	i->1	
(kons	u->1	
(kris	t->2	
(main	s->2	
(mer 	k->1	
(och 	p->1	
(reco	v->1	
(råde	t->1	
(se a	r->1	
(såso	m->1	
(t.ex	.->1	
(tyvä	r->1	
(ung.	 ->1	
(ÖVP)	 ->1	
(Öste	r->4	
(åter	v->1	
) "Ty	 ->1	
) (C5	-->1	
) (KO	M->2	
) (SE	K->1	
) (Ut	s->2	
) (fö	r->1	
) - A	l->1	
) - H	e->1	
) - S	a->1	
) 011	3->1	
) 055	0->1	
) 065	2->1	
) 158	 ->1	
) 344	 ->1	
) 519	 ->1	
) 520	 ->1	
) 522	 ->1	
) Att	 ->1	
) Bor	t->1	
) C5-	0->1	
) De 	d->1	
) Den	 ->5	
) Det	 ->2	
) Eft	e->2	
) FPÖ	:->1	
) Fru	 ->5	
) Frå	g->1	
) Får	 ->1	
) För	 ->1	
) Her	r->23	
) I S	c->1	
) I d	e->2	
) I g	å->1	
) I s	i->1	
) Ja,	 ->1	
) Jag	 ->14	
) Jör	g->1	
) Kom	m->1	
) Led	a->1	
) Låt	 ->2	
) Mit	t->1	
) Nej	,->1	
) När	 ->3	
) Om 	i->1	
) Sed	a->1	
) Tac	k->3	
) Tal	m->1	
) Thy	s->1	
) Tid	n->1	
) Und	e->1	
) Vad	 ->2	
) Ven	s->1	
) Vi 	s->1	u->1	
) ad 	h->1	
) av 	A->2	B->8	D->2	F->1	G->2	J->1	K->3	L->3	M->2	R->1	S->2	T->1	V->1	v->3	
) bät	t->1	
) eft	e->1	
) fin	a->1	
) frå	n->3	
) för	 ->3	e->1	r->1	
) had	e->1	
) har	 ->2	
) i G	e->1	
) i e	r->1	
) i h	e->1	
) i ä	n->1	
) inf	ö->3	
) inn	e->1	
) int	e->1	
) lik	a->1	
) min	s->1	
) och	 ->12	
) om 	g->1	
) på 	g->1	
) sam	t->1	
) sin	 ->1	
) som	 ->2	
) täc	k->1	
) zon	 ->1	
) Ära	d->1	
) är 	d->1	p->1	
)(Gen	o->1	
)(Par	l->9	
)(Tal	m->1	
)) (U	t->2	
)) (f	ö->1	
)) in	f->2	
))(Ge	n->1	
))(Pa	r->7	
)). V	i->1	
)).. 	-->1	
))..(	D->1	E->1	
)).Fr	u->1	
)).Ja	g->1	
))Fru	 ->1	
))Her	r->1	
))och	I->1	
), bi	d->1	
), de	t->1	
), me	n->1	
), oc	h->2	
), rå	d->1	
), so	m->2	
), tj	ä->1	
), tv	å->1	
), vi	l->1	
), är	 ->1	
). Vi	l->1	
).(EN	)->1	
).)Be	t->1	
).. (	E->1	
).. -	(->1	
)..(D	E->1	
)..(E	L->1	
).De 	f->1	m->1	
).Det	 ->2	t->1	
).Fru	 ->1	
).Frå	g->1	
).För	 ->1	
).Her	r->5	
).Jag	 ->3	
).Kan	 ->1	
).Kom	m->1	
).Lik	v->1	
).Vid	a->1	
).Vil	k->1	
)0003	 ->2	
)0066	 ->1	
)0598	 ->2	
)0662	 ->1	
):Ang	å->19	
); an	n->1	
); en	 ->1	
)? Ha	r->1	
)Andr	a->2	
)Angå	e->2	
)Ansv	a->1	
)Betä	n->8	
)Det 	ä->1	
)Fru 	t->8	
)Förf	a->1	
)Förs	l->1	
)Geme	n->1	
)Heat	o->1	
)Herr	 ->2	
)Jag 	f->1	s->2	
)Just	e->1	
)Konr	a->1	
)Näst	a->3	
)Olje	b->1	
)Refo	r->1	
)Säke	r->1	
)Tack	 ->1	
)Uttj	ä->1	
)].) 	H->1	
)].He	r->2	
)ochI	I->1	
)Åter	u->1	
, "af	f->1	
, "en	 ->1	
, "ne	 ->1	
, "ov	i->1	
, "se	 ->1	
, (Br	y->1	
, , a	t->1	
, 1 p	r->1	
, 10,	 ->1	
, 11 	o->1	
, 11,	 ->2	
, 12 	j->1	
, 12,	 ->3	
, 13,	 ->1	
, 15 	m->1	
, 15,	 ->2	
, 16 	o->1	
, 16,	 ->1	
, 166	 ->1	
, 167	 ->1	
, 18,	 ->1	
, 199	3->2	4->1	
, 2 o	c->1	
, 20,	 ->1	
, 22,	 ->1	
, 24 	o->1	
, 245	 ->1	
, 248	,->1	
, 27,	 ->1	
, 28,	 ->2	
, 30,	 ->1	
, 31 	o->1	
, 32,	 ->2	
, 34,	 ->1	
, 36,	 ->1	
, 37,	 ->2	
, 38,	 ->1	
, 4, 	6->1	
, 40,	 ->1	
, 42 	o->2	
, 44 	o->1	
, 46 	o->1	
, 50 	m->1	
, 500	 ->1	
, 56 	p->1	
, 6, 	7->1	
, 7, 	9->1	o->1	
, 8, 	9->1	
, 88 	o->1	
, 9, 	a->1	f->1	
, 95/	3->1	
, Als	a->1	
, Amo	k->1	s->1	
, Anv	e->1	
, Ari	a->3	
, Asi	e->1	
, BNI	,->1	
, Bel	g->2	
, Ber	g->2	
, Bre	m->1	
, Bro	k->1	
, Bry	s->1	
, Bus	h->1	
, Cos	t->1	
, Cux	h->1	
, Dag	m->1	
, Dan	m->1	
, Dar	m->1	
, Dav	i->1	
, Dim	i->1	
, Dub	l->1	
, ECH	O->1	
, EDD	,->1	
, EEG	,->2	
, EG-	d->1	
, Eft	a->1	
, Eri	k->1	
, Erk	k->1	
, Eur	a->4	o->4	
, Eva	n->2	
, Fin	l->1	
, Fra	n->1	
, För	e->1	
, Gar	g->1	
, Gil	-->1	
, Gin	o->1	
, Gra	c->1	
, Hag	u->1	
, Hai	d->1	
, Hav	e->1	
, Hel	s->1	
, II 	-->1	
, III	 ->1	
, IV 	-->1	
, Ile	-->1	
, Ing	e->1	
, Irl	a->1	
, Ita	l->2	
, Jap	a->1	
, Jon	a->1	c->1	
, Jor	d->1	
, Kan	a->1	
, Kar	l->1	
, Kaz	a->1	
, Koc	h->1	
, Kor	e->1	
, Kul	t->1	
, Kvä	k->1	
, La 	R->1	
, Lan	g->4	
, Lei	n->1	
, Lis	s->1	
, Lom	é->1	
, Lor	r->1	
, Lux	e->1	
, Mar	k->1	
, Mis	t->1	
, Mit	t->1	
, Ned	e->1	
, Nor	d->1	
, OLA	F->1	
, Obe	r->1	
, Oly	m->1	
, PVC	,->1	
, Pal	a->2	e->2	
, Pei	j->1	
, Raf	a->1	
, Rap	k->1	
, Rea	d->1	
, Red	i->1	
, Rot	h->1	
, SEK	(->2	
, Sag	e->1	
, Sam	m->1	
, Sch	e->2	
, Sha	r->1	
, Slo	v->1	
, Soa	r->1	
, Spa	n->3	
, Sto	c->1	
, Sve	r->1	
, Tan	i->1	
, Thy	s->1	
, Tom	 ->1	
, Tot	a->1	
, Tys	k->3	
, Uzb	e->1	
, V -	 ->1	
, Vla	a->1	
, Waf	f->1	
, Wes	t->1	
, Wie	n->1	
, Wul	f->1	
, Wye	 ->1	
, Zim	e->1	
, acc	e->2	
, ade	k->1	
, adm	i->1	
, akt	i->1	
, alb	a->1	
, ald	r->1	
, all	 ->1	a->3	d->2	m->1	t->16	
, amb	a->1	
, ana	l->1	
, and	e->1	r->2	
, anf	ö->1	
, ang	å->4	
, ann	a->3	
, ans	e->13	l->1	t->1	v->2	
, ant	i->1	
, anv	ä->2	
, arb	e->5	
, arr	o->1	
, art	i->1	
, att	 ->174	
, av 	E->1	G->1	a->1	d->7	e->1	f->2	k->1	m->1	p->1	s->4	t->1	v->2	
, avf	a->1	
, avs	e->1	i->1	l->1	t->2	
, ban	k->1	
, bar	a->3	n->1	r->1	
, bed	r->1	
, beg	r->2	ä->1	
, beh	a->1	
, bek	r->1	
, bel	ä->1	
, ben	s->1	
, ber	 ->2	o->2	ö->1	
, bes	k->1	l->3	t->2	
, bet	o->1	r->3	
, bev	a->1	i->3	
, bid	r->2	
, bil	a->1	i->1	t->1	
, bl.	a->16	
, bla	n->10	
, bli	 ->1	r->3	
, bor	d->4	g->1	t->4	
, bri	s->3	
, bro	t->1	
, brö	t->1	
, byg	g->1	
, byr	å->1	
, bär	 ->1	s->1	
, bäs	t->5	
, båd	e->13	
, bör	 ->15	j->4	
, civ	i->1	
, com	p->1	
, de 	2->1	b->2	d->1	e->1	f->3	g->2	h->1	i->1	k->2	l->2	m->3	o->1	p->1	r->2	s->7	t->2	y->2	ä->2	
, dec	e->3	
, del	a->1	g->1	s->4	t->1	v->1	
, dem	 ->1	o->8	
, den	 ->46	n->4	s->1	
, der	a->3	
, des	s->11	t->1	
, det	 ->110	t->6	
, dia	l->1	
, dif	f->1	
, dis	c->1	k->1	
, dju	p->1	r->3	
, dri	f->1	
, du 	b->1	
, dvs	.->43	
, däc	k->1	
, där	 ->51	a->2	e->2	f->3	i->5	m->1	p->1	
, då 	D->1	b->4	d->1	f->2	h->1	i->1	j->1	k->5	m->2	p->1	r->1	s->4	v->3	
, dål	i->1	
, död	 ->1	a->1	
, döl	j->1	
, eff	e->2	
, eft	e->120	
, eko	n->2	s->1	
, ele	k->1	
, ell	e->30	
, eme	d->1	
, en 	a->4	b->3	d->2	e->1	f->4	g->6	h->4	i->2	k->4	m->6	n->3	o->7	p->3	r->4	s->16	t->1	u->3	v->3	z->1	ö->4	
, end	a->1	
, ene	r->3	
, enh	e->1	
, enk	e->1	
, enl	i->19	
, era	 ->1	
, erb	j->1	
, erk	ä->1	
, eta	b->1	
, etc	.->2	
, eti	k->1	
, etn	i->1	
, ett	 ->37	
, eur	o->3	
, exa	k->1	m->1	
, exe	m->5	
, exi	s->1	
, fac	k->1	
, fak	t->3	
, fas	t->7	
, fic	k->2	
, fin	a->2	n->8	
, fly	g->1	
, fol	k->7	
, for	m->1	s->5	t->2	
, fra	m->27	
, fre	d->2	
, fri	 ->1	h->5	
, fru	 ->55	
, frä	m->12	
, frå	g->9	n->11	
, ful	l->1	
, fun	g->1	
, får	 ->10	
, fåt	t->1	
, föd	e->1	
, för	 ->197	b->4	d->3	e->13	f->2	h->2	l->1	o->2	p->1	r->2	s->15	u->10	v->1	ä->1	
, gam	l->1	
, gan	s->1	
, gar	a->1	
, gav	 ->1	
, ge 	e->1	
, ged	i->1	
, gem	e->3	
, gen	o->22	
, ger	 ->2	
, giv	a->1	e->2	
, gjo	r->2	
, glö	m->1	
, god	 ->1	
, gra	n->1	
, gru	n->4	
, grä	n->1	
, gul	t->1	
, gyn	n->1	
, gäl	l->1	
, gå 	i->1	t->1	
, går	 ->4	
, gåt	t->1	
, gör	 ->6	a->3	
, ha 	o->1	
, had	e->2	
, haf	t->1	
, ham	n->3	
, han	 ->3	d->6	s->3	
, har	 ->75	
, hel	a->2	s->1	t->4	
, her	r->145	
, het	t->1	
, hjä	l->2	
, hop	p->2	
, hos	 ->1	
, hot	e->1	
, hum	l->1	
, hur	 ->13	
, hus	 ->1	
, huv	u->3	
, hyg	i->1	
, hyr	d->1	
, hys	e->1	
, häl	e->1	f->1	s->1	
, hän	v->2	
, här	 ->3	,->1	
, häv	d->1	
, hål	l->2	
, hög	 ->1	a->1	e->1	
, höj	d->2	
, i A	u->1	
, i B	r->1	
, i I	C->1	
, i P	a->1	
, i S	e->1	
, i T	a->1	
, i a	l->4	n->3	
, i b	e->2	u->1	å->1	ö->1	
, i d	a->1	e->20	i->1	
, i e	g->2	n->10	r->4	t->3	
, i f	o->1	r->1	ö->7	
, i h	j->1	u->1	ä->1	
, i i	n->1	
, i j	a->1	u->1	
, i k	l->1	o->1	
, i l	a->1	i->4	
, i m	i->1	o->2	å->1	
, i n	i->1	
, i p	l->1	r->2	
, i r	e->3	å->1	
, i s	a->3	i->2	j->3	k->1	l->1	t->7	y->26	
, i t	v->1	
, i u	r->1	
, i v	i->6	
, i ö	v->2	
, ibl	a->2	
, ick	e->1	
, idr	o->1	
, igå	n->1	
, inb	e->3	
, ind	u->1	
, inf	o->2	r->2	ö->5	
, ing	a->1	e->3	
, ink	l->15	
, inl	e->1	å->1	
, inn	a->7	e->5	o->1	
, ino	m->15	
, inr	e->1	
, ins	a->1	k->1	y->1	
, int	e->72	r->1	ä->1	
, inv	a->1	e->1	
, iro	n->1	
, ja 	e->1	n->1	t->1	
, jag	 ->36	
, jor	d->2	
, ju 	l->1	m->2	
, jus	t->13	
, jäm	f->1	l->1	
, jär	n->8	
, kad	m->2	
, kal	l->3	
, kam	p->1	
, kan	 ->29	a->1	s->7	
, kao	s->1	
, kat	o->1	
, kid	n->1	
, kla	r->1	s->1	
, kof	f->1	
, kol	l->14	
, kom	 ->2	m->53	p->3	
, kon	c->1	k->6	s->3	t->1	
, koo	p->1	
, kor	n->1	t->2	
, kos	t->2	
, kra	f->2	v->1	
, kri	m->2	
, kro	a->1	m->1	
, krä	v->6	
, kul	t->5	
, kun	d->2	
, kur	s->1	
, kvi	c->2	n->1	
, kän	d->1	n->1	
, kär	a->45	e->1	n->2	
, lad	e->2	
, lan	d->2	
, led	a->3	d->1	e->1	
, leg	a->1	i->2	
, lem	l->1	
, lid	e->1	
, lik	a->2	n->1	s->30	
, lit	e->1	
, liv	s->2	
, lju	d->1	
, lok	a->1	
, läg	e->1	g->2	
, läk	e->1	
, läm	n->2	p->2	
, län	d->1	
, läs	 ->1	
, lån	g->7	
, låt	 ->4	
, lön	s->1	
, mak	t->1	
, man	 ->4	i->1	
, mar	k->2	
, mat	p->1	
, med	 ->66	a->15	b->1	e->1	i->3	k->1	l->5	
, mel	l->1	
, men	 ->314	,->1	a->5	i->1	
, mer	 ->7	
, mes	t->1	
, mik	r->1	
, mil	i->1	j->9	
, min	 ->2	a->29	d->1	i->1	o->1	s->1	
, mis	s->3	
, mod	e->3	
, mon	o->1	
, mor	a->1	d->1	
, mot	 ->5	o->1	t->1	
, mul	t->1	
, mus	s->1	
, myc	k->6	
, myn	d->1	
, män	n->3	s->6	
, må 	v->1	
, mån	g->1	
, mås	t->25	
, nar	k->1	
, nat	i->3	u->8	
, naz	i->1	
, ned	l->1	m->1	r->1	
, nej	 ->1	
, nek	a->1	
, nep	o->1	
, ni 	a->1	h->1	t->1	ä->1	
, nog	g->1	
, nor	d->1	
, nu 	m->1	n->3	t->2	
, ny 	s->1	
, nya	 ->3	
, nyl	i->1	
, näm	l->34	n->2	
, när	 ->64	i->1	m->4	
, näs	d->1	
, någ	o->28	r->1	
, nöd	v->1	
, oak	t->1	
, oan	s->1	
, oav	s->4	
, obe	g->1	r->3	
, och	 ->668	
, ock	s->8	
, off	e->1	
, oft	a->1	
, oli	k->1	
, oly	c->1	
, om 	1->1	D->1	E->2	a->7	b->1	d->26	e->4	f->3	g->2	h->4	i->3	j->4	k->2	m->6	n->5	o->1	p->4	r->2	s->3	t->1	u->1	v->12	ä->4	
, omd	i->1	
, ome	d->1	
, omf	a->2	
, omv	a->1	
, opp	o->1	
, ord	 ->1	f->3	
, ore	g->1	
, org	a->4	
, ost	r->1	
, osv	.->2	
, oty	d->1	
, par	l->5	t->2	
, pen	n->1	
, per	s->3	
, pla	n->1	
, plu	n->1	s->1	
, pol	i->2	
, pra	k->1	
, pre	c->12	s->3	
, pri	n->1	o->2	v->4	
, pro	b->1	d->1	f->2	
, pub	l->1	
, på 	E->1	O->1	a->3	b->2	d->4	e->8	g->16	i->2	j->1	l->1	m->1	n->1	p->1	s->8	v->2	z->1	
, påg	å->1	
, påm	i->2	
, påp	e->1	
, rap	p->1	
, ras	i->5	
, rea	k->1	
, reg	e->4	i->6	
, rek	o->2	
, ren	t->1	
, res	p->2	u->1	
, rev	i->1	
, rik	t->3	
, rom	e->1	
, räd	d->1	s->1	
, räk	n->2	
, rät	t->9	
, råd	e->11	
, rör	 ->1	e->1	i->1	l->1	
, rös	t->1	
, sad	e->2	
, sak	e->1	n->1	
, sal	i->1	
, sam	a->1	h->1	m->3	o->2	r->1	t->23	
, san	n->1	
, sat	s->1	
, se 	f->1	t->2	
, sed	a->3	
, sek	r->1	
, ser	 ->2	
, set	t->1	
, sex	 ->2	
, sin	 ->5	a->1	
, sis	t->1	
, sju	,->1	k->2	
, sjä	l->1	
, ska	d->1	l->19	p->2	
, ske	p->2	
, ski	l->1	
, skj	u->1	
, sko	g->1	
, skr	e->1	i->2	o->1	
, sku	l->18	
, sky	l->1	
, skä	l->1	
, slu	t->3	
, slä	p->1	
, sma	k->1	
, små	 ->1	
, sna	r->5	
, sne	d->2	
, soc	i->5	
, sol	d->1	i->1	
, som	 ->381	
, spa	r->2	
, spe	c->7	l->1	
, spo	r->1	
, sta	b->1	d->1	r->1	t->3	
, sti	l->1	
, sto	r->1	
, str	a->2	i->1	u->3	ä->1	
, sty	m->1	
, stå	l->1	r->1	
, stö	d->4	
, sva	r->2	
, svå	r->1	
, syr	i->1	
, säg	a->2	e->2	
, säk	e->29	
, säl	j->1	
, sär	s->34	
, så 	a->55	b->3	d->6	f->3	h->1	k->8	l->3	m->3	s->18	u->1	v->3	ä->5	
, såd	a->2	
, såg	v->1	
, sås	o->17	
, såv	i->2	ä->18	
, sök	e->1	
, sön	d->1	
, t.e	x->8	
, tac	k->9	
, tak	,->1	
, tal	a->1	r->1	
, tar	 ->4	
, teo	r->1	
, til	l->58	
, tio	t->1	
, tit	t->1	
, tjä	n->6	
, tob	a->1	
, tog	 ->1	
, tol	k->1	
, ton	 ->1	
, tor	t->2	
, tot	a->1	
, tra	k->1	n->15	
, tre	 ->1	d->1	t->1	
, tro	l->1	r->6	t->20	
, trå	k->1	
, tul	l->1	
, tur	k->1	
, tvi	n->1	v->2	
, tvä	t->1	
, två	 ->5	
, ty 	E->1	d->4	i->1	n->2	p->2	v->2	
, tyc	k->1	
, tyd	l->1	
, tyv	ä->3	
, täc	k->1	
, tän	k->1	
, tåg	 ->1	
, tål	a->1	
, töm	m->1	
, und	e->19	r->1	
, ung	a->1	d->3	
, uni	o->2	
, upp	 ->1	b->1	f->2	l->2	m->6	n->1	r->1	
, ur 	e->1	m->1	v->1	
, uta	n->131	r->1	
, utb	i->5	
, utf	ä->1	
, utg	ö->2	
, uti	f->2	
, utm	ä->1	
, utn	y->1	
, uto	m->3	
, utr	i->4	y->1	
, uts	k->1	
, utt	a->1	r->4	
, utv	e->3	i->4	
, utö	v->1	
, vad	 ->15	
, val	t->1	u->1	
, van	 ->1	
, var	 ->11	a->4	e->6	f->9	i->2	j->1	k->2	s->11	v->1	
, vat	t->2	
, vek	h->1	
, vem	 ->1	
, ver	k->4	
, vet	 ->4	
, vi 	a->1	b->7	e->1	f->1	g->1	h->6	k->1	l->2	m->3	s->6	u->1	v->4	ä->1	
, via	 ->3	
, vic	e->2	
, vid	 ->10	a->1	t->1	
, vik	t->1	
, vil	j->2	k->165	l->21	
, vis	a->5	k->1	s->1	
, von	 ->1	
, vor	e->3	
, väc	k->2	
, väd	j->2	
, väg	l->1	m->1	r->1	
, väl	k->2	
, vär	d->4	
, våg	a->1	
, vål	d->1	
, vår	 ->3	a->3	
, ytt	e->1	
, Île	-->1	
, äga	r->2	
, än 	e->2	t->1	
, änd	a->2	r->2	å->5	
, är 	E->1	a->11	b->2	d->28	e->19	f->6	h->1	i->3	k->2	m->1	n->3	o->3	r->3	s->2	t->2	v->2	
, ära	d->21	
, ärl	i->1	
, äve	n->60	
, å a	n->1	
, åny	o->1	
, år 	2->1	
, åt 	d->1	
, åta	l->1	
, åte	r->17	
, åtf	ö->1	
, åtg	ä->1	
, åtm	i->7	
, ått	a->1	
, öka	 ->1	r->1	
, öpp	e->2	n->1	
, öve	r->6	
,07 m	i->1	
,2 mi	l->1	
,2 oc	h->1	
,2 pr	o->1	
,3 pr	o->1	
,4 tr	i->1	
,42 m	i->1	
,487 	m->1	
,5 mi	l->1	
,5 pr	o->2	
,6 pr	o->1	
,7 pr	o->1	
,8 mi	l->3	
,8 ti	l->1	
,9 pr	o->1	
- "de	n->1	
- 'Va	d->1	
- (DE	)->1	
- (PT	)->14	
- , v	i->1	
- 199	7->7	8->6	9->13	
- 2,8	 ->1	
- 31 	m->1	
- 6 m	i->1	
- 80 	p->1	
- Alt	e->2	
- C4-	0->6	
- C5-	0->14	
- Cam	r->1	
- Den	 ->1	
- Dom	s->1	
- EU-	k->1	
- Fru	 ->1	
- Her	r->3	
- Kal	e->1	
- Kom	m->1	
- Par	l->1	
- Rev	i->1	
- Rik	t->1	
- Råd	e->1	
- Sav	e->2	
- all	a->2	t->3	
- ans	e->1	
- anv	ä->1	
- arb	e->1	
- att	 ->27	
- av 	E->1	a->1	d->1	e->2	m->2	n->1	s->1	
- bet	y->1	
- bid	r->1	
- bli	 ->1	
- bör	 ->1	
- cen	t->1	
- de 	b->1	e->1	f->1	k->1	n->3	s->2	v->1	
- del	t->1	v->1	
- den	 ->5	
- des	s->1	
- det	 ->26	t->7	
- doc	k->1	
- dvs	.->2	
- där	 ->2	
- då 	t->2	
- eft	e->2	
- eko	n->1	
- ell	e->6	
- en 	a->1	e->1	f->1	m->2	p->1	s->1	y->1	
- ena	s->1	
- end	a->1	
- enh	ä->1	
- enl	i->1	
- ett	 ->3	
- eve	n->1	
- exe	m->1	
- exi	s->1	
- fat	t->1	
- fic	k->1	
- fra	m->1	
- frä	m->1	
- frå	g->1	
- få 	v->1	
- får	 ->1	
- fåt	t->1	
- för	 ->12	d->1	e->1	f->1	v->1	
- gen	d->1	
- ger	 ->1	
- gäl	l->1	
- gör	a->2	
- han	 ->1	
- har	 ->9	
- hos	 ->1	
- hur	 ->3	
- här	 ->1	
- i K	o->1	
- i a	t->1	
- i d	e->1	
- i f	ö->1	
- i m	i->1	
- i r	e->1	
- i s	a->1	t->1	y->1	
- i u	t->1	
- i v	å->1	
- ida	g->1	
- inf	ö->2	
- inn	e->1	
- ino	m->2	
- ins	a->1	
- int	e->10	
- ja 	i->1	
- ja,	 ->2	
- jag	 ->12	
- jus	t->1	
- kan	 ->1	
- kna	p->1	
- kom	m->6	
- kon	k->1	
- kos	t->2	
- krä	v->1	
- lik	s->1	
- lin	o->1	
- lys	s->1	
- låt	 ->2	
- man	 ->2	
- mar	k->1	
- med	 ->4	a->1	
- men	 ->8	
- mer	a->1	
- min	s->1	
- mis	s->1	
- mon	i->1	
- mot	 ->1	
- mån	g->1	
- mås	t->1	
- nat	u->1	
- ny 	r->1	
- näm	l->2	n->1	
- när	 ->3	
- någ	o->6	
- och	 ->159	
- ock	s->1	
- off	r->1	
- om 	d->1	m->2	r->1	s->1	t->1	v->2	
- omr	å->1	
- ord	r->1	
- par	l->1	
- pre	c->1	
- pri	n->1	
- pro	g->1	
- på 	E->1	d->1	h->1	s->1	
- påm	i->1	
- rap	p->1	
- reg	e->1	
- res	u->1	
- ris	k->1	
- råd	e->1	
- rör	a->1	
- sad	e->1	
- sam	l->1	m->1	t->2	
- se 	b->1	
- ser	 ->2	
- sit	t->1	
- ska	l->2	
- sku	l->1	
- sna	r->1	
- sne	d->1	
- som	 ->26	
- sta	t->2	
- sto	r->1	
- syf	t->1	
- sys	t->1	
- säg	e->1	
- sär	s->1	
- så 	a->1	h->2	s->2	
- sål	e->1	
- sök	a->1	
- tac	k->1	
- tek	n->1	
- til	l->3	
- tro	r->2	t->1	
- tve	t->1	
- tän	k->1	
- und	e->1	
- uta	n->7	
- utg	ö->1	
- uts	t->1	
- utt	r->1	
- var	 ->2	
- ver	k->1	
- vet	 ->1	
- vi 	h->2	k->1	s->1	ä->1	ö->1	
- vik	t->1	
- vil	k->10	
- vis	a->1	
- väl	k->1	
- Öst	e->1	t->1	
- är 	a->3	d->1	i->1	j->1	s->1	
- äve	n->10	
- åtm	i->2	
- öpp	e->1	
- öve	r->4	
-(EN)	 ->1	
-, Sa	g->1	
-, at	t->1	
-, dä	r->1	
-, fö	r->1	
-, i 	s->1	
-, in	t->1	
-, me	n->1	
-, sk	a->1	
-, tr	a->1	
-, ut	a->1	b->1	
-, är	 ->1	
-0001	/->1	
-0002	/->1	
-0003	/->4	
-0004	/->2	
-0006	/->4	
-0007	/->3	
-0009	/->2	
-0010	/->2	
-0011	/->2	
-0012	/->2	
-0018	/->3	
-0020	/->1	
-0022	/->2	
-0040	/->1	
-0041	/->1	
-0045	/->2	
-0050	/->1	
-0069	/->1	
-0073	/->1	
-0078	/->1	
-0087	/->1	
-0095	/->1	
-0104	/->2	
-0105	/->2	
-0106	/->1	
-0107	/->2	
-0108	/->2	
-0120	/->1	
-0122	/->1	
-0167	/->1	
-0180	/->2	
-0208	/->2	
-0212	/->1	
-0305	/->1	
-0327	/->2	
-0333	/->2	
-0334	/->2	
-0341	/->2	
-0350	/->1	
-0351	/->1	
-0352	/->1	
-0715	/->1	
-0778	/->1	
-0780	/->1	
-0781	/->1	
-0782	/->1	
-0785	/->1	
-0786	/->1	
-0788	/->1	
-0791	/->1	
-0793	/->1	
-0795	/->1	
-0796	/->1	
-0798	/->1	
-0801	/->1	
-0805	/->1	
-0807	/->1	
-0808	/->1	
-0813	/->1	
-0817	/->1	
-0819	/->1	
-0829	/->1	
-1995	 ->1	,->1	
-1997	,->1	
-1999	.->1	
-2 da	g->1	
-2-om	r->1	
-2000	.->1	
-2002	)->2	
-2004	 ->1	.->1	
-2006	 ->6	,->3	.->8	
-4 pr	o->1	
-98/0	3->1	
-Alpe	s->1	
-Alst	h->2	
-Arde	n->1	
-Atla	n->1	
-Behr	e->7	
-Carp	e->1	
-Clau	d->1	
-DE).	(->1	
-DE- 	o->2	
-DE-g	r->4	
-DE-l	e->1	
-Delg	a->1	
-Exup	é->1	
-Fina	 ->2	.->1	
-Fran	c->2	
-Harr	i->1	
-Hein	z->1	
-I); 	e->1	
-II) 	o->1	
-Isra	e->1	
-Jørg	e->2	
-Kees	 ->1	
-Le B	e->1	
-Loir	e->1	
-Mann	e->1	
-Math	i->2	
-Norm	a->1	
-PM s	o->1	
-Plat	h->4	
-Robl	e->1	
-Roma	g->1	
-SS:s	 ->1	
-Shar	a->1	
-Shei	k->5	
-Syri	e->1	
-affä	r->3	
-alba	n->1	
-anal	y->6	
-anpa	s->1	
-avta	l->3	
-avvi	s->1	
-belo	p->1	
-bene	f->5	
-best	ä->1	
-bila	r->1	
-bild	e->1	
-bile	n->1	
-bist	å->1	
-brit	t->1	
-budg	e->1	
-bugg	e->1	
-damm	a->1	
-dans	k->1	
-de-F	r->2	
-de-L	o->1	
-dire	k->3	
-disk	r->2	
-doms	t->22	
-effe	k->1	
-el-S	h->1	
-enhe	t->1	
-er r	a->1	
-fall	e->1	
-fond	e->1	
-foss	i->1	
-fran	s->1	
-free	-->2	.->1	
-fråg	a->1	
-förd	r->19	
-före	t->1	
-förk	a->1	l->1	
-förs	ä->1	
-geme	n->1	
-geno	m->1	
-grup	p->20	
-how 	t->1	
-init	i->2	
-inst	i->4	r->1	
-intä	k->2	
-irlä	n->1	
-isra	e->1	
-kana	l->1	
-kata	s->3	
-koli	b->1	
-komm	i->3	
-kort	 ->10	,->1	e->9	
-kost	n->1	
-kris	e->3	
-krit	e->1	
-lags	t->1	
-land	e->1	
-leda	m->1	r->1	
-leks	a->1	
-lite	r->2	
-lobb	y->1	
-länd	e->5	
-mail	 ->1	
-mant	r->1	
-medb	o->4	
-mede	l->1	
-medl	e->1	
-meta	l->1	
-nati	o->1	
-nivå	.->1	
-noti	s->1	
-nytt	o->1	
-olyc	k->1	
-områ	d->8	
-ordf	ö->1	
-orga	n->3	
-posi	t->1	
-prog	r->25	
-prot	o->2	
-ramp	r->1	
-rasi	s->1	
-rege	r->1	
-regi	m->1	o->5	
-rätt	 ->2	.->1	e->1	
-råde	t->4	
-shop	,->1	
-situ	a->1	
-skan	d->1	
-soci	a->2	
-spri	d->3	
-stat	e->2	l->9	u->2	
-stip	e->1	
-stop	-->1	
-stru	k->1	
-stöd	,->2	
-syst	e->1	
-sänd	a->1	e->2	
-tal 	p->1	
-tale	t->7	
-tals	k->1	
-test	e->1	
-text	e->1	
-tran	s->1	
-uppd	r->1	
-utvi	d->1	
-van 	G->1	
-värl	d->1	
-zon 	V->1	
-zone	n->1	r->1	
. (EL	)->1	
. (EN	)->23	
. (FI	)->1	
. (FR	)->12	
. (PT	)->1	
. -(E	N->1	
. 11 	m->1	
. 11,	3->1	
. 11.	0->3	A->1	E->1	K->1	
. 12.	0->6	
. 120	 ->1	
. 13.	0->1	
. 15.	0->2	
. 17.	3->1	
. 19.	5->1	
. 20.	2->1	
. 21.	0->1	5->1	
. 7 l	e->1	
. 7).	.->1	
. All	a->1	
. Av 	d->1	
. De 	h->1	s->1	
. Den	 ->5	n->4	
. Der	a->1	
. Des	s->3	
. Det	 ->31	t->8	
. Där	 ->3	e->1	f->2	
. Då 	b->1	t->1	
. Eft	e->2	
. En 	b->1	d->1	p->2	v->1	
. Enl	i->1	
. Equ	q->1	
. Ett	 ->1	
. Eur	o->4	
. Fog	 ->1	
. Fra	n->1	
. Fru	 ->2	
. Frä	m->1	
. Föl	j->1	
. För	 ->2	
. Gut	e->1	
. Han	 ->1	
. Her	r->3	
. Hon	 ->1	
. Hur	 ->1	
. Här	 ->3	
. Hål	l->1	
. I r	e->1	
. I s	t->1	
. Ing	a->1	
. Ini	t->1	
. Int	e->1	
. Jag	 ->10	
. Kom	m->1	
. Kos	t->1	
. Kär	a->1	
. Låt	 ->1	
. Man	 ->2	
. Men	 ->14	,->1	
. Ned	e->1	
. Ni 	h->1	
. Näs	t->1	
. Och	 ->4	
. Off	e->1	
. Om 	m->1	
. Par	l->1	
. Pro	c->1	
. På 	s->1	
. Råd	s->1	
. Sko	g->1	
. Skä	l->1	
. Som	 ->2	
. Syr	i->1	
. Så 	l->1	r->1	
. Tac	k->1	
. Til	l->1	
. USA	.->1	
. Var	f->1	j->1	k->1	
. Vi 	h->3	k->2	s->1	v->4	
. Vi,	 ->1	
. Vil	k->1	
. Vår	a->1	t->1	
. Wal	e->1	
. aid	s->1	
. ans	v->1	
. arb	e->1	
. art	i->1	
. att	 ->12	
. av 	v->1	
. avs	k->2	
. bet	o->1	
. de 	e->1	
. den	 ->3	
. des	s->2	
. det	 ->2	
. en 	t->1	
. enh	e->1	
. ert	,->1	
. ett	 ->3	
. for	d->1	
. får	 ->1	
. för	 ->4	d->1	s->3	
. gen	o->1	
. gra	n->1	
. gör	a->1	
. hos	 ->1	
. hur	 ->1	
. i M	e->1	
. i d	e->1	
. i e	n->1	
. i p	r->1	
. idé	n->1	
. inf	ö->1	
. inn	a->1	
. ino	m->1	
. int	e->3	
. jag	 ->1	
. kri	g->1	
. kun	n->1	
. kän	n->1	
. man	 ->2	
. med	 ->2	
. men	 ->1	
. min	d->1	
. mit	t->2	
. när	 ->5	
. nät	v->1	
. och	 ->2	
. olj	e->2	
. om 	d->1	n->1	v->1	
. på 	d->1	t->1	v->1	
. ska	l->2	
. sko	g->1	
. sof	t->1	
. spe	c->1	
. sto	r->1	
. säk	e->1	
. tra	n->1	
. und	e->1	
. utf	a->1	
. vad	 ->1	
. var	j->1	v->1	
. vi 	m->1	
. Ämn	a->1	
. Änd	å->1	
. Änn	u->1	
. Äve	n->1	
. Åtg	ä->1	
. Öst	t->1	
. änn	u->1	
. är 	v->1	
. öst	b->1	
." Är	a->1	
."Det	 ->1	
."I d	e->1	
."Jag	 ->1	
."Med	 ->1	
.(App	l->5	
.(Arb	e->1	
.(DA)	 ->2	
.(DE)	 ->2	
.(EL)	 ->2	
.(EN)	 ->10	
.(ES)	 ->1	
.(FR)	 ->6	
.(IT)	 ->3	
.(Ihå	l->1	
.(Liv	l->2	
.(NL)	 ->4	
.(PT)	 ->1	
.(Par	l->5	
.(Pro	t->1	
.(Sam	m->4	
.(Tal	m->7	
.) He	r->3	
.) Ta	l->1	
.).De	 ->1	
.).He	r->1	
.)And	r->2	
.)Ans	v->1	
.)Bet	ä->8	
.)Fru	 ->5	
.)För	f->1	s->1	
.)Gem	e->1	
.)Hea	t->1	
.)Her	r->1	
.)Jus	t->1	
.)Olj	e->1	
.)Ref	o->1	
.)Säk	e->1	
.)Åte	r->1	
., de	t->1	
., fr	å->1	
., äv	e->1	
.- (D	E->1	
.- (P	T->10	
.- De	n->1	
.- Fr	u->1	
.- He	r->2	
.. (E	L->1	N->15	
.. (F	I->1	R->9	
.. -(	E->1	
.. De	t->1	
.. Fr	u->1	
.. Fö	r->1	
.. He	r->1	
.. Pr	o->1	
.. Ta	c->1	
.. Vi	 ->1	
..(DA	)->2	
..(DE	)->2	
..(EL	)->1	
..(EN	)->5	
..(ES	)->1	
..(FR	)->5	
..(IT	)->1	
..(NL	)->3	
..(Ta	l->5	
..).D	e->1	
...(T	a->5	
...).	D->1	
....(	T->1	
...Fr	u->1	
...He	r->1	
...Lå	t->1	
..Fru	 ->1	
..Her	r->5	
..Låt	 ->1	
..Tac	k->1	
..Vi 	ä->1	
.00.(	S->2	
.00.)	A->1	O->1	
.00.D	e->1	
.00.F	a->1	ö->1	
.00.O	M->1	
.00.S	a->1	t->2	
.00.T	i->1	r->1	
.05 o	c->1	
.1 då	 ->1	
.1 i 	A->1	E->1	r->1	
.1 oc	h->2	
.1 vi	l->1	
.1 öv	e->1	
.1) e	f->1	
.1.1 	ö->1	
.1.Fö	r->1	
.1.Vi	 ->1	
.12.0	0->1	
.14 e	u->1	
.15 m	a->1	
.18 m	i->1	
.1998	 ->1	
.2 i 	A->2	S->1	a->1	f->1	
.2 oc	h->1	
.2).K	a->1	
.25.)	J->1	
.3 EG	-->1	
.3 bl	i->1	
.3 in	t->1	
.3, n	å->1	
.30, 	o->1	
.3; d	e->1	
.4 in	t->1	
.4.De	 ->1	
.4.Fö	r->1	
.50 o	c->1	
.55)U	t->1	
.8 i 	d->1	
.90 p	r->1	
.?Ans	e->1	
.Acce	p->1	
.Aher	n->1	
.Akti	v->1	
.Aldr	i->1	
.Alla	 ->21	
.Alld	e->1	
.Allm	ä->4	
.Allt	 ->16	f->1	s->1	
.Alte	n->2	
.Amer	i->1	
.Amst	e->1	
.Andr	a->4	
.Angå	e->1	
.Anhå	l->1	
.Anle	d->1	
.Anna	r->4	
.Anse	r->1	
.Ansv	a->3	
.Anta	l->2	
.Anvä	n->1	
.Arab	v->1	
.Arbe	t->2	
.Arti	k->2	
.Att 	a->1	b->1	d->2	f->1	g->2	h->1	i->1	k->1	l->2	m->2	r->1	s->1	t->2	u->3	v->1	
.Atta	c->1	
.Av 4	1->1	
.Av a	l->4	v->1	
.Av b	e->2	
.Av d	e->13	
.Av e	n->1	
.Av s	a->2	
.Av v	i->2	
.Avbr	o->1	
.Avgå	n->1	
.Avsa	t->1	
.Avse	r->1	
.Avsl	u->13	
.Bako	m->2	
.Bara	 ->4	
.Bedr	ä->2	
.Bedö	m->2	
.Befo	r->1	
.Bekv	ä->1	
.Bere	n->2	
.Bero	e->1	
.Besl	u->3	
.Betr	ä->6	
.Betä	n->16	
.Bevi	s->1	
.Bili	n->1	
.Bill	o->2	
.Bilt	i->2	
.Bist	å->1	
.Blan	d->7	
.Bord	e->2	
.Bosä	t->1	
.Bret	a->1	
.Bris	t->3	
.Brit	t->1	
.Brys	s->1	
.Budg	e->1	
.Bygg	e->1	
.Bäst	a->1	
.Båda	 ->5	
.CSU:	s->1	
.Cent	r->2	
.Corp	u->1	
.Cunh	a->1	
.DEBA	T->1	
.Dage	n->3	
.Dagl	i->2	
.Dala	i->1	
.Danm	a->1	
.De 1	4->1	5->1	
.De a	k->1	l->2	n->3	v->1	
.De b	e->4	i->1	
.De d	a->1	i->1	r->1	
.De e	u->2	
.De f	a->2	i->2	l->5	r->3	å->1	ö->7	
.De g	j->1	r->2	ä->1	
.De h	a->9	å->1	
.De i	n->1	
.De k	a->6	o->3	r->2	
.De l	a->1	ö->1	
.De m	i->1	y->1	å->5	
.De n	o->1	u->1	y->4	ä->1	
.De o	l->2	
.De p	e->1	o->2	
.De r	e->1	
.De s	e->4	i->2	k->5	l->1	o->3	t->7	
.De t	o->2	u->2	v->1	
.De u	p->2	t->2	
.De v	a->2	i->1	
.De ä	r->4	
.De å	t->2	
.Dels	 ->1	
.Delv	i->1	
.Den 	1->1	2->1	a->20	b->4	c->1	e->15	f->17	g->9	h->16	i->2	k->13	l->2	m->10	n->7	o->5	p->3	r->5	s->16	t->10	u->2	v->8	ä->9	å->3	ö->1	
.Denn	a->47	e->1	
.Dera	s->1	
.Dess	 ->2	a->30	u->24	
.Det 	a->11	b->28	c->2	d->2	e->9	f->97	g->30	h->51	i->11	j->1	k->45	l->5	m->27	n->2	o->1	p->9	r->22	s->66	t->6	u->2	v->40	ä->316	å->3	ö->3	
.Det,	 ->1	
.Deta	l->1	
.Dets	a->1	
.Dett	a->196	
.Dire	k->7	
.Disk	u->1	
.Dock	 ->2	
.Doku	m->1	
.Doms	t->2	
.Där 	b->1	f->2	h->3	k->1	l->1	m->1	ä->1	
.Dära	v->2	
.Däre	f->4	m->5	
.Därf	ö->91	
.Däri	 ->1	g->2	
.Därm	e->4	
.Däru	t->1	
.Därv	i->1	
.Då d	e->1	
.Då f	i->1	r->1	å->1	
.Då g	i->1	
.Då h	a->2	
.Då k	a->3	o->4	
.Då m	å->1	
.Då o	c->1	
.Då s	k->1	y->1	
.Då v	a->1	i->1	
.Då ä	r->2	
.Då ö	v->1	
.EG-d	o->3	
.EKSG	-->1	
.EU m	å->1	
.EU ä	r->1	
.EU-k	o->2	
.EU-o	r->1	
.Effe	k->5	
.Efte	r->36	
.Ekon	o->2	
.Emel	l->8	
.En a	l->3	n->6	s->1	v->5	
.En b	o->2	ä->1	
.En d	e->6	
.En f	r->2	ö->2	
.En g	e->1	
.En k	a->1	n->1	o->3	
.En m	a->1	e->1	
.En r	a->2	e->2	
.En s	a->1	i->1	u->1	y->1	ä->1	å->4	
.En u	p->1	
.En v	a->1	e->1	i->3	ä->2	
.En ö	k->1	v->1	
.Enba	r->1	
.Enda	s->9	
.Enke	l->1	
.Enli	g->31	
.Er a	n->1	
.Erfa	r->2	
.Erik	a->4	
.Ert 	p->1	
.Ett 	a->10	d->2	e->4	f->4	h->1	l->1	m->1	n->2	o->2	p->1	s->9	t->2	v->3	å->1	
.Euro	j->2	n->1	p->47	s->1	
.Even	t->1	
.Exce	p->1	
.Exem	p->1	
.Expe	r->2	
.FEO 	b->1	
.FPÖ 	h->1	ä->1	
.FPÖ:	s->2	
.Fack	f->3	
.Fakt	u->4	
.Farl	i->1	
.Fasc	i->1	
.Fela	k->1	
.Fem 	l->1	
.Fina	n->2	
.Finn	s->2	
.Fler	a->3	t->1	
.Flor	e->3	
.Folk	 ->2	
.Fors	k->2	
.Fram	 ->1	f->2	s->2	t->2	å->1	
.Fran	s->2	
.Fred	s->1	
.Frih	e->1	
.Fru 	B->1	L->1	M->1	P->1	k->3	l->1	t->46	
.Frut	e->1	
.Fråg	a->31	e->2	o->1	
.Från	 ->2	
.Fyrt	i->1	
.Får 	j->1	
.Följ	a->4	d->1	
.För 	1->1	a->28	b->1	d->90	e->2	f->2	i->1	k->1	m->7	n->7	o->5	p->1	s->3	t->4	u->1	v->7	å->1	ö->3	
.Förb	u->2	
.Förd	e->1	r->2	
.Före	b->1	d->7	n->4	t->2	
.Förh	o->3	
.Förl	u->1	
.Förm	o->1	
.Förp	a->1	
.Förs	i->1	l->6	t->17	ö->1	
.Fört	j->1	r->1	
.Föru	t->7	
.Förv	a->1	i->2	ä->1	
.Förä	n->1	
.Geme	n->3	
.Gene	r->1	
.Geno	m->25	
.Ger 	d->1	
.Give	t->2	
.Gola	n->1	
.Grat	u->1	
.Grek	l->2	
.Grun	d->1	
.Grup	p->2	
.Gäll	a->1	
.Gå h	e->1	
.Gör 	v->2	
.Hade	 ->2	
.Haid	e->1	
.Han 	a->1	b->1	h->7	s->3	t->1	ä->3	
.Hand	e->1	l->2	
.Hans	 ->2	
.Har 	m->1	r->1	v->1	
.Hela	 ->3	
.Helt	 ->2	
.Herr	 ->268	
.Hist	o->2	
.Hit 	h->3	
.Hitt	i->2	
.Hon 	h->2	s->1	
.Hopp	e->1	
.Hult	e->1	
.Hur 	f->2	g->1	h->1	k->1	l->1	m->2	s->16	
.Huru	v->1	
.Huvu	d->7	
.Hyck	l->1	
.Händ	e->2	
.Här 	b->4	f->3	g->1	h->4	i->1	k->5	m->2	r->1	s->1	t->2	v->3	ä->1	
.Härm	e->1	
.Häro	m->1	
.Höge	r->1	
.I Am	s->1	
.I Eu	r->4	
.I Fr	a->1	
.I He	l->1	
.I Ir	l->2	
.I It	a->1	
.I Ne	d->1	
.I Ra	p->1	
.I Ti	b->1	
.I Ty	s->1	
.I al	l->3	
.I an	d->1	n->2	
.I ap	r->1	
.I ar	t->1	
.I av	s->1	v->2	
.I be	t->4	
.I da	g->17	
.I de	 ->2	n->18	t->31	
.I di	r->1	
.I eg	e->4	
.I en	 ->7	l->3	
.I et	t->2	
.I fl	e->1	
.I fo	r->1	
.I fr	a->1	å->5	
.I fö	r->6	
.I gå	r->2	
.I ju	n->1	
.I kl	a->1	
.I ko	m->2	n->1	
.I li	k->6	
.I mi	n->1	t->1	
.I mo	r->2	t->2	
.I må	l->1	
.I no	v->2	
.I nä	s->2	
.I oc	h->4	
.I pa	r->1	
.I pr	i->1	o->1	
.I ra	p->2	
.I re	a->1	g->1	s->4	v->1	
.I rä	t->1	
.I rå	d->1	
.I sa	m->3	
.I si	n->1	t->1	
.I sj	ä->4	
.I sl	u->2	
.I st	i->1	r->1	ä->8	
.I sy	n->1	s->1	
.I så	 ->2	d->1	
.I tj	u->1	
.I up	p->1	
.I ut	b->1	
.I va	r->2	
.I ve	r->1	
.I vi	l->2	s->2	t->2	
.I vo	n->1	
.I vä	n->2	
.I vå	r->6	
.I än	d->1	
.I öv	r->3	
.Ibla	n->3	
.Idén	 ->1	
.Ille	g->1	
.Immi	g->1	
.Indu	s->1	
.Infö	r->4	
.Inga	 ->1	
.Inge	n->9	t->2	
.Init	i->1	
.Inne	b->1	h->1	
.Inom	 ->10	
.Inre	 ->1	s->1	
.Inrä	t->1	
.Insa	t->2	
.Inte	 ->11	r->1	
.Irla	n->1	
.Isra	e->1	
.Ital	i->1	
.Ja e	l->1	
.Ja t	i->1	
.Ja, 	f->1	j->1	s->1	
.Jack	s->1	
.Jacq	u->1	
.Jag 	a->51	b->31	d->7	e->1	f->40	g->9	h->86	i->8	k->42	l->3	m->23	n->3	o->1	p->5	r->10	s->98	t->115	u->25	v->154	ä->46	ö->7	
.Jonc	k->1	
.Jord	b->1	
.Ju m	i->1	
.Just	 ->8	e->1	
.Jämf	ö->1	
.Jäms	t->1	
.Kafo	r->1	
.Kan 	k->4	m->1	n->4	v->1	
.Kans	k->6	
.Karl	 ->1	
.Kata	s->1	
.Kinn	o->3	
.Knap	p->1	
.Koch	 ->1	
.Kode	n->1	
.Kom 	i->1	
.Komm	e->4	i->97	u->1	
.Komp	r->1	
.Konk	r->1	u->12	
.Kons	e->1	t->1	u->3	
.Konv	e->1	
.Kort	 ->2	
.Koso	v->1	
.Kost	n->3	
.Krav	 ->1	e->2	
.Kult	u->7	
.Kvan	t->1	
.Kvin	n->1	
.Kära	 ->4	
.Kärn	a->1	k->1	
.La R	é->1	
.Land	s->1	
.Lang	e->1	
.Leda	m->2	
.Ledn	i->1	
.Lika	 ->1	s->2	
.Likr	i->1	
.Liks	o->6	
.Likv	ä->1	
.Litt	e->1	
.Livs	m->3	
.Lyck	a->1	l->1	
.Lynn	e->1	
.Lägg	 ->2	
.Länd	e->1	
.Lån 	a->1	
.Lång	r->1	
.Låt 	e->1	i->1	m->31	o->14	v->1	
.Majo	r->1	
.Malt	a->2	
.Man 	b->8	f->2	g->2	h->4	i->1	j->1	k->11	l->1	m->12	r->1	s->3	t->2	u->3	v->1	
.Mann	e->1	
.Marg	a->1	
.Mark	n->4	
.Maxi	m->2	
.Med 	a->3	d->8	e->2	f->1	h->5	o->2	s->2	t->6	
.Meda	n->4	
.Medb	e->1	o->2	
.Medg	e->1	
.Medl	e->9	
.Mell	a->3	
.Men 	-->2	C->1	E->1	a->5	b->2	d->52	e->4	f->7	g->1	h->6	i->8	j->28	k->5	m->4	n->5	o->4	p->4	s->12	t->2	u->4	v->28	ä->3	å->1	
.Men,	 ->2	
.Ment	a->1	
.Mer 	s->1	v->1	ä->1	
.Milj	ö->1	
.Min 	a->6	f->5	g->5	k->1	p->1	s->4	t->2	u->1	å->1	ö->1	
.Mina	 ->16	
.Minn	s->1	
.Mins	k->1	
.Mitt	 ->2	
.Mora	l->1	
.Mot 	b->4	d->4	
.Myll	e->1	
.Mynd	i->3	
.Männ	i->4	
.Märk	l->1	
.Måhä	n->1	
.Måle	t->2	
.Mång	a->10	
.Möjl	i->2	
.Nati	o->3	
.Natu	r->14	
.Nej,	 ->1	
.Ni a	g->1	
.Ni b	e->2	o->1	
.Ni f	r->1	ö->2	
.Ni h	a->7	
.Ni k	a->2	o->3	ä->2	
.Ni l	ä->1	
.Ni m	å->4	
.Ni s	a->2	k->2	ä->1	
.Ni t	a->2	
.Ni v	e->2	
.Niel	s->1	
.Nivå	n->1	
.Norm	e->1	
.Nu a	n->2	
.Nu b	e->1	
.Nu f	i->1	ö->1	
.Nu h	a->6	o->1	
.Nu k	a->2	
.Nu m	å->1	
.Nu t	i->1	
.Nu v	e->1	ä->1	
.Nu ä	r->7	
.Nu å	t->1	
.Nume	r->1	
.Nuva	r->1	
.Nya 	r->1	
.Nyli	g->1	
.När 	a->2	b->2	d->30	e->1	f->1	j->6	k->1	m->6	p->1	s->1	t->1	v->12	
.Näst	a->1	
.Någo	n->1	t->1	
.Någr	a->2	
.Nåja	,->1	
.Nödv	ä->1	
.OK, 	d->1	
.OLAF	,->2	
.OMRÖ	S->2	
.Oavs	e->2	
.Ober	o->2	
.Och 	E->1	S->1	a->2	d->20	e->2	g->1	i->2	j->8	k->1	m->1	n->4	o->1	s->6	t->1	v->8	ä->1	
.Ocks	å->2	
.Offe	n->2	
.Ofta	 ->1	
.Om 5	0->1	
.Om E	u->1	
.Om S	c->1	y->1	
.Om a	l->3	
.Om b	e->1	
.Om d	e->21	o->1	
.Om e	n->1	r->1	t->2	
.Om f	o->1	
.Om g	e->1	i->1	
.Om i	n->1	
.Om j	a->2	
.Om k	a->1	o->4	
.Om l	a->1	
.Om m	a->10	
.Om n	i->6	
.Om p	a->2	
.Om r	e->1	å->1	
.Om s	l->1	y->1	
.Om t	r->1	v->1	
.Om u	p->1	
.Om v	i->22	
.Omrö	s->15	
.Onöd	i->1	
.Ord 	s->1	
.Orde	n->1	r->1	t->1	
.Ordf	ö->7	
.Orka	n->2	
.Oron	 ->1	
.Orov	ä->1	
.Orsa	k->2	
.Oz h	a->1	
.PPE-	D->2	
.Para	g->1	
.Parl	a->21	
.Pers	o->4	
.Plan	e->1	
.Plas	t->2	
.Pläd	e->1	
.Port	u->2	
.Prec	i->5	
.Pres	e->1	
.Prob	l->8	
.Proc	e->2	
.Prod	i->3	u->2	
.Prog	r->1	
.Proj	e->2	
.Punk	t->2	
.På a	l->1	
.På d	e->19	
.På e	t->1	
.På g	r->1	
.På l	a->1	
.På m	a->1	i->1	å->1	
.På o	m->2	
.På p	a->1	
.På s	a->3	i->3	å->4	
.På u	p->1	
.På v	i->2	
.Rapp	o->3	
.Rasi	s->1	
.Reak	t->1	
.Reda	n->3	
.Refo	r->6	
.Rege	r->4	
.Regi	o->1	
.Rent	 ->2	
.Rest	e->2	
.Resu	l->5	
.Retr	o->1	
.Revi	s->2	
.Rika	 ->1	
.Rikt	l->3	
.Risk	e->1	
.Rope	t->1	
.Roth	-->2	
.Rumä	n->1	
.Räkn	a->1	
.Rätt	s->2	
.Råde	t->16	
.Samh	ä->2	
.Samm	a->7	
.Samo	r->1	
.Samt	i->14	
.Sann	i->4	o->1	
.Save	 ->1	N->1	
.Schr	o->1	
.Schu	l->1	
.Schü	s->1	
.Seda	n->15	
.Sett	 ->1	
.Sist	 ->2	
.Situ	a->3	
.Sju 	ä->1	
.Själ	v->2	
.Skad	o->1	
.Skal	l->3	
.Skot	t->1	
.Skul	l->4	
.Skyd	d->1	
.Slut	l->34	r->1	s->3	
.Små 	o->1	
.Småf	ö->1	
.Snab	b->1	
.Snar	a->1	
.Soci	a->3	
.Som 	E->1	a->2	b->1	e->7	f->3	h->1	j->7	k->3	l->2	m->1	n->6	p->2	s->3	u->1	v->2	
.Soml	i->3	
.Stab	i->1	
.Stat	e->5	i->1	l->2	
.Stor	a->2	m->2	
.Stra	f->1	
.Stru	k->1	
.Strä	v->1	
.Stäm	m->1	
.Stål	s->1	
.Stöd	 ->2	e->3	s->1	
.Stör	r->2	s->2	
.Subv	e->2	
.Svep	e->1	
.Syft	e->6	
.Syri	e->1	
.Säg 	m->1	
.Säke	r->1	
.Särs	k->2	
.Så b	l->1	
.Så d	e->3	
.Så e	n->1	r->1	
.Så f	r->1	
.Så h	ä->1	
.Så j	a->3	
.Så k	a->1	o->1	
.Så l	ä->3	å->1	
.Så n	å->1	
.Så s	e->1	o->2	ä->1	
.Så t	i->1	
.Så v	a->1	i->4	å->1	
.Så ä	r->1	v->2	
.Såda	n->2	
.Såle	d->4	
.Sång	e->1	
.Såso	m->2	
.Såvä	l->1	
.TV-b	i->1	
.Ta d	ä->1	
.Tack	 ->14	,->13	.->1	
.Tadz	j->1	
.Tala	r->1	
.Tank	e->3	
.Terr	o->1	
.Thea	t->2	
.Thys	s->1	
.Tidi	g->1	
.Till	 ->23	s->2	v->3	ä->3	å->6	
.Titt	a->1	
.Tong	i->1	
.Topp	m->2	
.Torv	 ->1	e->1	
.Tran	s->2	
.Tre 	ä->1	
.Tror	 ->1	
.Trot	s->16	
.Trov	ä->1	
.Träd	 ->1	
.Tuse	n->1	
.Tvär	t->3	
.Två 	v->1	ä->1	
.Ty e	n->1	
.Ty i	n->1	
.Ty s	o->1	
.Ty u	n->1	
.Ty v	a->1	i->2	
.Tydl	i->1	
.Tyvä	r->9	
.Tänk	 ->1	
.Unda	n->3	
.Unde	r->27	
.Ungd	o->1	
.Unge	f->2	
.Unio	n->5	
.Uppe	n->1	
.Uppf	ö->1	
.Uppg	i->3	
.Uppr	ä->1	
.Ur d	e->2	
.Ur e	n->1	
.Ur p	a->1	
.Utan	 ->3	
.Utbi	l->2	
.Utde	l->1	
.Utes	t->1	
.Utfo	r->2	
.Utfö	r->1	
.Utgi	f->1	
.Utif	r->1	
.Utma	n->2	
.Utnä	m->1	
.Utsk	o->2	
.Utve	c->1	
.Utvi	d->1	
.Vad 	a->2	b->9	d->1	e->1	f->1	g->14	h->1	j->3	k->6	m->1	s->8	t->1	u->1	v->6	ä->3	
.Vada	n->1	
.Vale	n->2	t->1	
.Van 	H->1	
.Vanl	i->1	
.Var 	d->1	f->2	h->1	o->2	s->1	
.Vare	 ->2	
.Varf	ö->11	
.Varj	e->5	
.Vem 	b->1	v->1	
.Vems	 ->2	
.Verk	s->1	
.Vete	n->1	r->1	
.Vi a	c->1	l->1	n->17	r->1	v->5	
.Vi b	e->23	i->1	o->1	ö->11	
.Vi d	e->2	i->5	r->1	
.Vi e	r->1	u->1	
.Vi f	a->1	i->3	o->2	ä->1	å->9	ö->10	
.Vi g	e->1	j->1	o->2	r->1	ö->3	
.Vi h	a->80	o->6	y->1	ä->2	å->1	
.Vi i	 ->6	n->7	
.Vi j	a->1	
.Vi k	a->25	o->19	r->8	u->1	ä->3	
.Vi l	a->2	i->1	ö->1	
.Vi m	e->4	o->1	å->73	
.Vi o	r->1	
.Vi p	a->1	l->1	
.Vi r	a->1	e->1	i->1	ä->2	ö->1	
.Vi s	a->1	e->5	i->1	k->19	o->1	t->7	v->2	ä->3	
.Vi t	a->5	i->2	r->2	v->2	y->4	ä->2	
.Vi u	n->1	p->6	t->1	
.Vi v	a->3	e->15	i->28	ä->7	
.Vi ä	n->1	r->28	
.Vi ö	n->1	
.Via 	s->1	
.Vid 	E->1	b->1	d->3	e->2	l->1	m->2	s->2	
.Vida	r->7	
.Vikt	e->1	
.Vilj	a->1	
.Vilk	a->9	e->1	
.Vill	 ->4	k->1	
.Vind	e->1	
.Viss	a->10	e->2	t->1	
.Vitb	o->3	
.Von 	W->1	
.Värd	e->1	
.Väst	m->1	r->1	
.Vår 	e->1	g->5	i->2	o->1	r->2	u->2	ö->1	
.Våra	 ->7	
.Vårt	 ->5	
.Worl	d->1	
.Ytte	r->3	
.a. a	r->1	t->1	
.a. b	e->1	
.a. d	e->1	
.a. e	n->1	t->1	
.a. f	å->1	ö->4	
.a. g	e->1	ö->1	
.a. i	 ->2	
.a. k	r->1	
.a. m	e->1	
.a. n	ä->3	
.a. o	l->1	m->1	
.a. p	å->1	
.a. s	k->2	t->1	
.a. u	n->1	
.a. v	a->1	
.d. Ö	s->1	
.d. ö	s->1	
.d., 	f->1	
.ex. 	E->1	F->1	N->1	U->1	a->2	d->2	e->1	i->1	k->2	m->2	n->2	o->1	p->1	u->1	v->1	
.g.a.	 ->1	
.k. a	n->1	
.k. i	n->1	
.k. s	k->1	o->1	
.komm	i->1	
.m. a	v->2	
.m. d	e->1	
.m. i	 ->1	
.m. ä	n->1	r->1	
.m., 	d->1	
.m.Oc	h->1	
.o.m.	 ->6	,->1	
.Än e	n->3	
.Ända	 ->1	
.Ändr	a->1	i->13	
.Ändå	 ->4	
.Ännu	 ->1	
.Äntl	i->1	
.Är I	s->1	
.Är d	e->11	
.Är k	o->1	
.Är r	å->1	
.Är s	t->1	
.Ärad	e->3	
.Även	 ->31	
.Å ED	D->1	
.Å an	d->10	
.Å en	a->2	
.År 1	9->4	
.År 2	0->1	
.Året	 ->1	
.Åtag	a->1	
.Åter	i->1	v->1	
.Åtgä	r->2	
.ÖVP 	(->1	
.Ögon	b->2	
.Ökad	 ->1	
.Öste	r->2	
.Över	 ->1	v->1	
.Övri	g->1	
/00 -	 ->1	
/00) 	f->1	
/00):	A->1	
/0012	(->1	
/0013	(->1	
/0083	 ->1	
/0090	(->1	
/0106	(->2	
/0169	(->2	
/0194	(->2	
/0228	(->1	
/0240	(->2	
/0318	(->1	
/0352	(->1	
/0370	(->2	
/0371	(->2	
/0803	(->1	
/0805	(->1	
/0825	(->2	
/1/19	9->2	
/1998	,->2	
/1999	 ->25	)->14	
/2000	 ->2	)->24	
/2123	(->1	
/2127	(->1	
/3 av	 ->1	
/35/E	G->4	
/409 	o->1	
/43.T	y->1	
/55/E	G->2	
/591/	E->2	
/60/9	2->1	
/71 a	n->1	
/71/E	G->1	
/728/	E->1	
/75 o	m->1	
/92 o	c->1	
/95.F	r->1	
/98 -	 ->1	
/98-9	8->1	
/99 (	H->1	
/99 -	 ->1	
/99 b	e->1	
/99 o	c->2	
/99) 	f->1	o->1	
/99):	A->18	
/99)A	n->2	
/99.J	a->1	
/EG a	t->1	
/EG o	m->2	
/EG s	k->1	
/EG u	p->1	
/EG, 	E->1	f->1	v->1	
/EKSG	,->2	
/Euro	p->1	
/NGL-	g->2	
/Nord	i->2	
/Oil-	p->1	
/den 	b->1	
/elle	r->1	
/halv	o->1	
/intä	k->1	
/rike	d->1	
/samm	a->1	
/år)?	 ->1	
/år, 	n->1	
0 - 1	9->3	
0 - C	4->1	5->1	
0 - d	e->1	
0 000	 ->11	
0 Enl	i->1	
0 ans	t->1	
0 arb	e->2	
0 arr	a->1	
0 att	 ->1	
0 bar	a->1	
0 bil	j->1	
0 det	a->1	
0 dol	l->1	
0 dom	a->1	
0 död	a->1	
0 ell	e->2	
0 ens	k->1	
0 eur	o->1	
0 fra	m->1	
0 frå	n->4	
0 fåg	l->2	
0 för	 ->1	
0 gul	d->1	
0 gån	g->1	
0 han	d->1	
0 har	 ->2	
0 hek	t->1	
0 i a	r->3	
0 i f	ö->4	
0 inn	e->3	
0 jan	u->1	
0 jun	i->1	
0 jur	i->1	
0 kan	 ->1	
0 kil	o->4	
0 km 	l->1	m->1	
0 km,	 ->1	
0 km.	T->1	
0 läg	g->1	
0 med	 ->1	l->1	
0 mil	j->17	
0 min	u->2	
0 mot	 ->1	
0 nya	 ->1	
0 när	 ->1	
0 och	 ->7	
0 oli	k->1	
0 pro	c->37	
0 på 	f->1	
0 rim	m->1	
0 ska	d->1	
0 sku	l->1	
0 som	 ->2	
0 stå	r->1	
0 tib	e->1	
0 ton	 ->8	/->2	
0 uta	n->1	r->1	
0 var	 ->1	
0 º C	.->1	
0 änd	r->7	
0 är 	h->1	l->1	s->2	v->1	
0 år 	a->1	e->2	i->1	o->1	s->1	ä->1	
0 år.	J->1	Ä->1	
0 års	 ->1	
0 åtg	ä->1	
0" so	m->1	
0" ti	l->2	
0".De	 ->1	
0".Vi	 ->1	
0(CNS	)->2	
0(COD	)->3	
0) av	 ->20	
0) fr	å->1	
0) fö	r->1	
0) oc	h->1	
0).Fr	å->1	
0).Ja	g->1	
0):An	g->1	
0, 12	,->1	
0, 22	,->1	
0, 32	,->1	
0, 46	 ->1	
0, dä	r->1	
0, fö	r->1	
0, i 	d->1	
0, mo	t->1	
0, må	s->1	
0, oc	h->1	
0, sk	j->1	
0, så	 ->1	
0, äv	e->1	
0- oc	h->1	
0-200	4->1	6->16	
0-bug	g->1	
0-pro	g->4	
0-tal	 ->1	e->7	s->1	
0.(Sa	m->2	
0.)An	s->1	
0.)Ol	j->1	
0.25.	)->1	
0.4.F	ö->1	
0.Den	 ->1	
0.Det	 ->2	t->3	
0.Fas	c->1	
0.Fru	 ->1	
0.För	 ->1	s->1	
0.Jag	 ->2	
0.Kom	m->1	
0.Man	 ->1	
0.Men	 ->1	
0.OMR	Ö->1	
0.Sam	o->1	
0.Sto	r->1	
0.Str	a->1	
0.Til	l->1	
0.Tra	n->1	
0.Vi 	d->1	
0/199	8->1	9->3	
0/200	0->3	
0/92 	o->1	
0/99 	-->1	b->1	
0/99)	 ->1	:->1	
00 - 	1->3	d->1	
00 00	0->6	
00 En	l->1	
00 ar	b->2	r->1	
00 at	t->1	
00 ba	r->1	
00 bi	l->1	
00 do	l->1	
00 få	g->2	
00 fö	r->1	
00 ha	n->1	r->2	
00 he	k->1	
00 in	n->2	
00 ki	l->4	
00 km	 ->2	,->1	.->1	
00 lä	g->1	
00 me	d->1	
00 mi	l->4	
00 mo	t->1	
00 nä	r->1	
00 oc	h->4	
00 ol	i->1	
00 pr	o->1	
00 på	 ->1	
00 sk	a->1	u->1	
00 so	m->1	
00 st	å->1	
00 ti	b->1	
00 to	n->10	
00 ut	a->1	
00 va	r->1	
00 än	d->4	
00 är	 ->4	
00 år	 ->1	
00" s	o->1	
00" t	i->2	
00".D	e->1	
00".V	i->1	
00) a	v->20	
00) f	r->1	ö->1	
00) o	c->1	
00).F	r->1	
00).J	a->1	
00):A	n->1	
00, d	ä->1	
00, f	ö->1	
00, i	 ->1	
00, m	o->1	å->1	
00, s	å->1	
00, ä	v->1	
00-20	0->17	
00-bu	g->1	
00-pr	o->4	
00-ta	l->4	
00.(S	a->2	
00.)A	n->1	
00.)O	l->1	
00.De	n->1	t->4	
00.Fa	s->1	
00.Fr	u->1	
00.Fö	r->2	
00.Ja	g->2	
00.Ma	n->1	
00.Me	n->1	
00.OM	R->1	
00.Sa	m->1	
00.St	o->1	r->1	
00.Ti	l->1	
00.Tr	a->1	
00.Vi	 ->1	
000 -	 ->3	
000 E	n->1	
000 a	r->2	t->1	
000 b	a->1	
000 f	å->2	ö->1	
000 h	a->2	e->1	
000 i	n->2	
000 k	i->1	m->3	
000 l	ä->1	
000 m	e->1	i->1	o->1	
000 n	ä->1	
000 o	c->2	
000 p	å->1	
000 s	k->1	o->1	t->1	
000 t	i->1	o->10	
000 u	t->1	
000 v	a->1	
000 ä	r->4	
000" 	s->1	t->2	
000".	D->1	V->1	
000) 	a->20	f->1	o->1	
000).	F->1	J->1	
000, 	d->1	f->1	i->1	m->2	s->1	ä->1	
000-2	0->17	
000-b	u->1	
000-p	r->4	
000-t	a->4	
000.D	e->4	
000.F	r->1	ö->1	
000.J	a->2	
000.M	a->1	e->1	
000.V	i->1	
0001/	2->1	
0002/	2->1	
0003 	-->2	
0003/	2->4	
0004/	1->1	2->1	
0006/	0->2	2->2	
0007/	2->3	
0009/	2->2	
000Nä	s->1	
001 ä	n->1	
001, 	m->1	
001/2	0->1	
0010/	2->2	
0011/	2->2	
0012(	C->1	
0012/	2->2	
0013(	C->1	
0018/	2->2	9->1	
002 (	K->1	
002 f	a->1	
002) 	-->2	
002, 	k->1	s->1	
002. 	J->1	
002.H	e->1	
002.M	i->1	
002.P	å->1	
002.V	i->1	
002/2	0->1	
0020/	1->1	
0022/	2->2	
003 -	 ->2	
003/2	0->4	
003?H	e->1	
004 i	n->1	
004.D	e->1	
004.K	o->1	
004/1	9->1	
004/2	0->1	
0040/	9->1	
0041/	9->1	
0045/	0->1	2->1	
0050/	2->1	
006 [	K->1	
006 f	ö->2	
006 g	ä->1	
006 k	o->1	
006 l	i->1	
006 o	c->1	
006 s	å->1	
006 t	a->1	o->1	
006 å	t->1	
006, 	f->1	m->1	n->1	s->2	
006.D	e->2	
006.E	n->1	
006.F	r->1	
006.H	e->1	
006.J	a->2	
006.M	a->1	
006.T	a->1	
006/0	0->2	
006/2	0->2	
0066 	-->1	
0069/	1->1	
007, 	r->1	
007/2	0->3	
0073/	1->1	
0078/	1->1	
008 t	o->2	
0083 	(->1	
0087/	1->1	
009/2	0->2	
0090(	C->1	
0095/	1->1	
00Näs	t->1	
01 än	t->1	
01, m	å->1	
01/20	0->1	
01/99	)->1	
010 e	l->1	
010/2	0->2	
0104/	1->2	
0105/	1->2	
0106(	C->2	
0106/	1->1	
0107/	1->2	
0108/	1->2	
011/2	0->2	
0113 	-->1	
012 e	n->1	
012(C	O->1	
012/2	0->2	
0120/	9->1	
0122/	1->1	
013(C	N->1	
0167/	1->1	
0169(	C->2	
018/2	0->2	
018/9	8->1	
0180/	1->2	
0194(	C->2	
02 (K	O->1	
02 fa	k->1	
02) -	 ->2	
02, k	o->1	
02, s	o->1	
02. J	a->1	
02.He	r->1	
02.Mi	n->1	
02.På	 ->1	
02.Vi	 ->1	
02/20	0->1	
020/1	9->1	
0208/	1->2	
0212/	1->1	
022/2	0->2	
0228(	C->1	
0240(	C->2	
03 - 	C->2	
03(CN	S->1	
03/20	0->4	
0305/	1->1	
0318(	S->1	
0327/	1->2	
0333/	1->2	
0334/	1->2	
0341/	1->2	
0350/	1->1	
0351/	1->1	
0352(	C->1	
0352/	1->1	
0370(	C->2	
0371(	C->2	
03?He	r->1	
04 in	l->1	
04.De	t->1	
04.Ko	m->1	
04/19	9->3	
04/20	0->1	
040/9	9->1	
041/9	9->1	
045/0	0->1	
045/2	0->1	
05 i 	E->1	
05 oc	h->1	
05 ti	l->1	
05(CN	S->1	
05/19	9->3	
05/99	)->1	
050/2	0->1	
0550 	-->1	
0598 	-->2	
06 [K	O->1	
06 fö	r->2	
06 gä	l->1	
06 ko	m->1	
06 li	g->1	
06 oc	h->1	
06 så	 ->1	
06 ta	s->1	
06 to	t->1	
06 åt	e->1	
06(CO	D->2	
06, f	ö->1	
06, m	e->1	
06, n	ä->1	
06, s	o->2	
06.De	t->2	
06.En	l->1	
06.Fr	å->1	
06.He	r->1	
06.Ja	g->2	
06.Ma	n->1	
06.Ta	c->1	
06/00	)->2	
06/19	9->1	
06/20	0->2	
0652 	-->1	
066 -	 ->1	
0662 	-->1	
069/1	9->1	
07 mi	l->1	
07, r	e->1	
07/19	9->2	
07/20	0->3	
07/99	)->1	
0715/	9->1	
073/1	9->1	
0778/	9->1	
078/1	9->1	
0780/	9->1	
0781/	9->1	
0782/	9->1	
0785/	9->1	
0786/	9->1	
0788/	9->1	
0791/	9->1	
0793/	9->1	
0795/	9->1	
0796/	9->1	
0798/	9->1	
08 to	n->2	
08/19	9->4	
08/99	)->1	
0801/	9->1	
0803(	C->1	
0805(	C->1	
0805/	9->1	
0807/	9->1	
0808/	9->1	
0813/	9->1	
0817/	9->1	
0819/	9->1	
0825(	C->2	
0829/	9->1	
083 (	C->1	
087/1	9->1	
09 oc	h->1	
09/20	0->2	
090(C	O->1	
094/1	9->2	
095/1	/->2	9->1	
0Näst	a->1	
1 000	 ->2	
1 400	 ->1	
1 ang	å->1	
1 då 	a->1	
1 eft	e->1	
1 frå	n->3	
1 ger	 ->1	
1 i A	m->1	
1 i E	G->1	
1 i a	r->1	
1 i k	a->1	
1 i r	a->1	
1 jan	u->9	
1 jul	i->1	
1 jun	i->1	
1 maj	 ->1	
1 mar	s->3	
1 men	 ->1	
1 mil	j->1	
1 och	 ->18	
1 ock	s->1	
1 om 	d->1	
1 pro	c->7	
1 ris	k->1	
1 sep	t->1	
1 sta	t->2	
1 ur 	e->1	
1 urv	a->1	
1 uta	n->1	
1 vil	k->1	
1 änt	l->1	
1 är 	n->1	
1 år 	e->1	
1 öve	r->1	
1(COD	)->2	
1) ef	t->1	
1, 12	,->2	
1, 2 	o->1	
1, 4,	 ->1	
1, at	t->1	
1, fö	r->1	
1, må	s->1	
1, oc	h->1	
1, sk	a->1	
1,2 o	c->1	
1,2 p	r->1	
1,3 p	r->1	
1,4 t	r->1	
1-2 d	a->1	
1-omr	å->4	
1-reg	i->5	
1-sta	t->2	
1.00.	(->1	)->1	F->1	T->1	
1.1 d	å->1	
1.1 o	c->2	
1.1 ö	v->1	
1.1.F	ö->1	
1.1.V	i->1	
1.3 E	G->1	
1.3 b	l->1	
1.3 i	n->1	
1.3, 	n->1	
1.3; 	d->1	
1.55)	U->1	
1.Alt	e->1	
1.Exc	e->1	
1.För	 ->1	
1.Jag	 ->1	
1.Kul	t->1	
1.Vi 	a->1	
1/199	8->1	9->4	
1/200	0->3	
1/3 a	v->1	
1/99)	 ->1	:->2	A->1	
1/EG 	o->1	
1/EKS	G->2	
10 00	0->2	
10 el	l->2	
10 fr	a->1	
10 i 	a->1	
10 ja	n->1	
10 ka	n->1	
10 mi	l->2	
10 pr	o->4	
10 ri	m->1	
10 so	m->1	
10 än	d->1	
10 är	 ->1	
10 år	.->1	
10, 1	2->1	
10.Ko	m->1	
10/20	0->2	
100 d	o->1	
100 k	i->1	
100 m	i->1	
100 o	l->1	
100 p	r->1	
100 ä	n->4	
104/1	9->2	
105 i	 ->1	
105 t	i->1	
105/1	9->2	
106(C	O->2	
106/1	9->1	
107/1	9->2	
108/1	9->2	
11 i 	a->1	
11 ja	n->2	
11 mi	l->1	
11 oc	h->1	
11 st	a->1	
11, 1	2->2	
11, f	ö->1	
11,3 	p->1	
11.00	.->3	
11.Al	t->1	
11.Ex	c->1	
11.Ku	l->1	
11/20	0->2	
110 i	 ->1	
113 -	 ->1	
115 m	i->1	
12 en	l->1	
12 fr	å->1	
12 in	n->1	
12 ja	n->1	
12 mi	l->1	
12 må	n->1	
12 oc	h->1	
12 pr	o->1	
12 st	a->1	
12(CO	D->1	
12, 1	3->1	5->1	
12, d	v->1	
12, t	r->1	
12.00	.->7	
12/19	9->1	
12/20	0->2	
12/99	 ->2	.->1	
120 m	i->1	
120/9	9->1	
122/1	9->1	
123 p	e->1	
123(C	O->1	
1244 	o->1	
1244.	I->1	J->1	
125 m	i->1	
1260/	9->1	
127(C	O->1	
13 (E	U->1	
13 - 	C->1	
13 00	0->1	
13 Am	s->1	
13 fe	b->1	
13 i 	E->1	f->1	
13 ja	n->1	
13 ny	a->1	
13 ok	t->1	
13 pr	o->2	
13 sa	m->1	
13 är	 ->1	
13(CN	S->1	
13, 2	8->2	
13.05	 ->1	
13.Fö	r->1	
13/19	9->1	
13/99	)->1	
130 d	o->1	
133.2	 ->1	
138.4	.->1	
14 eu	r->1	
14 fe	b->5	
14 le	d->1	
14 me	d->5	
14 oc	h->1	
14 se	p->1	
14 ti	l->1	
14, e	l->1	
14/19	9->1	
140 j	u->1	
14094	/->2	
143 o	m->1	
15 av	 ->1	
15 ma	r->2	
15 mi	l->1	
15 ol	i->2	
15 om	 ->1	
15 pr	o->3	
15 rä	c->1	
15 se	p->1	
15 st	a->1	
15 år	.->1	
15, 1	6->2	
15.00	.->2	
15/98	-->1	
150 g	u->1	
150 o	c->1	
158 -	 ->1	
158 i	 ->1	
158).	D->1	
158.1	 ->1	
16 00	0->1	
16 oc	h->3	
16 pe	r->1	
16 pr	o->1	
16 ra	d->1	
16) s	a->1	
16, 2	0->1	
164 r	ö->1	
166 e	m->1	
167 m	i->3	
167/1	9->1	
169(C	O->2	
17 de	c->2	
17 mi	l->1	
17 oc	h->1	
17 ok	t->1	
17 så	 ->1	
17, 1	8->1	
17, s	å->1	
17.30	,->1	
17.Sl	u->1	
17/99	)->1	
170 m	i->1	
174 t	u->1	
1762 	u->1	
1762.	M->1	
18 de	c->1	
18 hä	n->1	
18 i 	b->1	
18 mi	l->2	
18 må	n->1	
18 no	v->3	
18(SY	N->1	
18, 2	7->1	
18/20	0->2	
18/98	 ->1	
180 m	i->1	
180/1	9->2	
19 - 	C->1	
19 de	p->1	
19 ma	r->1	
19 pr	o->1	
19 so	m->1	
19 är	 ->1	
19.50	 ->1	
19/99	)->1	
1917 	o->1	
1923,	 ->1	
193 o	c->1	
1930-	t->1	
194(C	O->2	
194.D	e->1	
1945.	F->1	
1948.	D->1	
195 m	i->1	
1957 	(->1	
1957.	E->1	
1967 	h->1	i->1	m->1	o->2	
1967,	 ->1	
1969 	o->1	
1976 	e->1	
1977 	-->1	
1982,	 ->1	
1982.	I->1	
1986 	h->1	o->1	
1986.	Å->1	
1989,	 ->1	
1990 	u->1	
1990.	D->1	
1991 	e->1	g->1	o->1	
1992 	s->2	å->1	
1992,	 ->1	
1993 	h->1	o->1	u->1	
1993,	 ->1	
1993-	1->2	
1993.	O->1	
1993?	F->1	
1994 	e->1	h->1	o->2	
1994,	 ->1	
1994-	1->1	
1995 	(->1	h->1	k->1	r->1	s->1	å->1	
1995,	 ->2	
1995-	1->1	
1996 	-->1	e->1	h->1	i->1	l->1	o->1	v->2	ä->1	å->2	
1996,	 ->2	
1996.	D->1	E->1	J->1	M->1	O->1	
1997 	(->1	-->1	d->1	f->1	h->2	i->1	l->1	o->6	p->1	t->2	u->1	ä->1	å->1	
1997)	 ->1	
1997,	 ->2	
1997.	-->1	.->1	B->1	D->2	I->1	M->1	N->1	V->2	
1997/	0->7	
1997?	D->1	
1997N	ä->1	
1998 	g->1	h->1	k->1	o->6	r->1	s->1	u->3	v->2	ä->2	
1998)	 ->3	
1998,	 ->3	
1998-	2->2	
1998.	 ->1	P->1	S->1	
1998/	0->4	
1999 	-->26	a->4	d->1	e->1	f->2	g->1	h->5	i->4	j->1	k->4	n->1	o->4	p->1	r->1	s->1	t->1	u->3	v->3	ä->1	å->1	ö->1	
1999"	.->1	
1999)	 ->17	.->1	0->3	
1999,	 ->7	
1999-	2->2	
1999.	 ->1	.->1	D->3	E->2	F->3	J->1	K->1	U->1	V->1	
1999/	0->11	2->2	
1999:	 ->1	
1:a å	r->1	
2 (KO	M->1	
2 - C	4->3	
2 - v	i->1	
2 000	 ->1	
2 400	 ->1	
2 av 	P->1	
2 bla	n->1	
2 bli	r->1	
2 dag	a->1	
2 dec	e->1	
2 ell	e->1	
2 enl	i->1	
2 eur	o->1	
2 fak	t->1	
2 frå	n->2	
2 har	 ->1	
2 i A	m->2	
2 i S	c->1	
2 i a	r->3	
2 i f	ö->3	
2 i r	e->1	
2 i s	y->1	
2 i t	j->1	
2 inn	e->2	
2 jan	u->1	
2 mil	j->5	
2 mån	a->1	
2 och	 ->9	
2 pro	c->4	
2 pun	k->1	
2 rik	t->1	
2 skr	e->1	
2 som	 ->2	
2 sta	t->1	
2 und	e->1	
2 upp	h->1	
2 års	 ->1	
2(CNS	)->1	
2(COD	)->1	
2) - 	A->1	S->1	
2) fö	r->1	
2).Ka	n->1	
2, 11	,->1	
2, 13	,->1	
2, 15	,->1	
2, 24	 ->1	8->1	
2, 37	,->2	
2, de	t->1	
2, dv	s->1	
2, el	l->1	
2, en	 ->1	
2, fr	a->1	
2, i 	a->1	r->1	
2, ko	m->1	
2, lä	g->1	
2, sk	ä->1	
2, so	m->2	
2, ti	l->1	
2, tr	e->1	
2, vi	l->2	
2,487	 ->1	
2,5 m	i->1	
2,6 p	r->1	
2,8 m	i->1	
2-omr	å->3	
2-stö	d->1	
2. Ja	g->1	
2.00.	(->1	D->1	O->1	S->3	T->1	
2.1 i	 ->1	
2.2 i	 ->1	
2.Det	 ->1	
2.Her	r->1	
2.I e	n->1	
2.Isr	a->1	
2.Jag	 ->1	
2.Man	 ->1	
2.Men	 ->1	
2.Min	a->1	
2.På 	d->1	
2.Vi 	p->1	
2.Äve	n->1	
2/199	9->3	
2/200	0->5	
2/43.	T->1	
2/99 	o->2	
2/99)	:->1	
2/99.	J->1	
20 - 	C->1	
20 00	0->1	
20 eu	r->1	
20 fr	å->1	
20 gå	n->1	
20 mi	l->2	n->1	
20 ny	a->1	
20 pr	o->3	
20 º 	C->1	
20 än	d->1	
20 år	 ->5	
20, 2	2->1	
20.25	.->1	
20/19	9->1	
20/99	 ->1	
200 0	0->4	
200 å	r->1	
2000 	-->3	E->1	a->2	f->1	h->2	i->1	l->1	m->2	n->1	o->2	s->2	u->1	v->1	ä->4	
2000"	 ->3	.->2	
2000)	 ->22	.->2	
2000,	 ->7	
2000-	2->17	b->1	p->4	t->4	
2000.	D->4	F->2	J->2	M->1	V->1	
2000N	ä->1	
2001 	ä->1	
2001,	 ->1	
2002 	(->1	f->1	
2002)	 ->2	
2002,	 ->2	
2002.	 ->1	H->1	M->1	P->1	V->1	
2003?	H->1	
2004 	i->1	
2004.	D->1	K->1	
2006 	[->1	f->2	g->1	k->1	l->1	o->1	s->1	t->2	å->1	
2006,	 ->5	
2006.	D->2	E->1	F->1	H->1	J->2	M->1	T->1	
2007,	 ->1	
2010 	e->1	
2012 	e->1	
208/1	9->2	
21 ja	n->1	
21 ju	l->1	
21 oc	k->1	
21 om	 ->1	
21 st	a->1	
21 är	 ->1	
21 år	 ->1	
21.00	.->1	
21.55	)->1	
212/1	9->1	
2123(	C->1	
2127(	C->1	
21:a 	å->1	
22 - 	C->1	
22 av	 ->1	
22 ri	k->1	
22, 2	4->1	
22, i	 ->1	
22, v	i->1	
22,5 	m->1	
22.Äv	e->1	
22/19	9->1	
22/20	0->2	
226 i	 ->1	
228(C	N->1	
23 de	c->1	
23 in	n->1	
23 pe	r->1	
23(CO	S->1	
23, e	f->1	
23,7 	p->1	
24 ny	a->2	
24 oc	h->1	
24 ok	t->1	
24 pr	o->1	
240(C	N->2	
244 o	c->1	
244.I	 ->1	
244.J	a->1	
245 o	c->1	
248, 	2->1	
25 gr	a->1	
25 me	s->1	
25 mi	l->1	n->1	
25 om	r->1	
25 pr	o->7	
25 ti	l->1	
25(CN	S->2	
25.)J	u->1	
25.De	s->1	
250 m	i->1	
255 i	 ->3	n->1	
26 "p	å->1	
26 i 	a->1	
26 in	d->1	
26 me	d->1	
26 no	v->1	
26 oc	h->1	
26 pr	o->1	
260/9	9->1	
262 e	u->1	
27 de	c->1	
27 fa	l->1	
27 lä	n->1	
27 oc	h->1	
27 pr	o->2	
27(CO	S->1	
27, 3	4->1	
27/19	9->2	
28 fr	å->1	
28 ju	l->1	
28 ny	a->1	
28 pr	o->1	
28(CN	S->1	
28, 3	0->1	2->1	
28/EG	,->1	
280 i	 ->4	
280.4	.->1	
28:e 	å->1	
29 dö	d->1	
29 fr	å->1	
29 lä	n->1	
29 mi	n->1	
29, 3	1->1	
29/99	)->1	
299.2	 ->2	
3 (CO	D->1	
3 (EU	-->1	
3 - C	4->1	5->2	
3 000	 ->5	
3 Ams	t->1	
3 EG-	f->1	
3 av 	s->1	t->1	
3 bli	r->1	
3 dec	e->1	
3 feb	r->2	
3 frå	n->1	
3 för	 ->1	
3 har	 ->1	
3 hör	 ->1	
3 i E	U->1	
3 i d	i->1	
3 i f	ö->1	
3 inn	e->1	
3 int	e->1	
3 jan	u->2	
3 maj	 ->1	
3 nya	 ->1	
3 och	 ->4	
3 okt	o->2	
3 om 	a->1	
3 per	s->2	
3 pro	c->6	
3 pun	k->1	
3 sam	t->1	
3 ute	s->1	
3 är 	v->1	
3(CNS	)->2	
3(COS	)->1	
3, 19	9->1	
3, 28	,->2	
3, 7,	 ->1	
3, ef	t->1	
3, nå	g->1	
3,7 p	r->1	
3,8 m	i->1	
3,8 t	i->1	
3,9 p	r->1	
3-199	5->2	
3-4 p	r->1	
3-lit	e->2	
3.05 	o->1	
3.1) 	e->1	
3.2 o	c->1	
3.8 i	 ->1	
3.Frå	g->1	
3.För	b->1	
3.I ö	v->1	
3.Om 	a->1	
3.Tyd	l->1	
3/199	9->4	
3/200	0->4	
3/75 	o->1	
3/99)	:->2	
30 do	m->1	
30 fr	å->1	
30 i 	a->1	
30 in	n->1	
30 ju	n->1	
30 me	d->1	
30 mi	l->1	
30 oc	h->1	
30 pr	o->3	
30, 3	2->1	
30, o	c->1	
30-ta	l->1	
300 s	k->1	
305/1	9->1	
31 fr	å->1	
31 ja	n->1	
31 ma	j->1	r->1	
31 oc	h->2	
314 l	e->1	
318(S	Y->1	
32 mi	l->1	
32, 2	4->1	
32, 3	7->2	
32.Ja	g->1	
327/1	9->2	
33 00	0->2	
33 av	 ->1	
33 fr	å->1	
33 fö	r->1	
33 i 	d->1	
33 oc	h->1	
33.2 	o->1	
33/19	9->2	
332, 	2->1	
333/1	9->2	
334/1	9->2	
34 i 	a->1	
34 sk	a->1	
34 ti	l->1	
34 år	 ->1	
34, 3	6->1	
34.1.	1->1	
34/19	9->2	
341/1	9->2	
344 -	 ->1	
35 fr	å->1	
35 mi	l->5	
35.Så	d->1	
35/EG	 ->3	,->1	
350 m	i->1	
350/1	9->1	
351/1	9->1	
352(C	N->1	
352/1	9->1	
36 fr	å->1	
36, 3	8->1	
367 0	0->1	
37 fr	å->1	
37 i 	a->1	
37 pr	o->1	
37, 4	2->2	
37.2 	i->1	
37/60	/->1	
370 m	i->1	
370(C	O->2	
371(C	O->2	
38 fr	å->1	
38 fö	r->1	
38 oc	h->2	
38, 4	4->1	
38.4.	D->1	
38: f	o->1	
39 fr	å->1	
39 i 	M->1	
39 pr	o->1	
39, 4	0->1	
3: fö	r->1	
3; de	t->1	
3?Frå	g->1	
3?Her	r->1	
4 - C	5->1	
4 000	 ->1	
4 c i	 ->1	
4 en 	a->1	
4 ett	 ->1	
4 eur	o->1	
4 feb	r->5	
4 frå	n->1	
4 har	 ->1	
4 i E	G->1	K->1	
4 i a	n->1	
4 i d	e->2	i->1	
4 inl	e->1	
4 int	e->1	
4 jun	i->2	
4 led	a->1	
4 lik	s->1	
4 med	l->5	
4 nya	 ->2	
4 när	 ->1	
4 och	 ->8	
4 okt	o->1	
4 pro	c->5	
4 rös	t->1	
4 sep	t->1	
4 ska	t->1	
4 til	l->2	
4 tri	l->1	
4 tus	e->1	
4 år 	s->1	
4(COD	)->2	
4, 11	 ->1	,->1	
4, 36	,->1	
4, 6,	 ->1	
4, el	l->1	
4, fö	r->1	
4, ko	n->1	
4, oc	h->1	
4-001	8->1	
4-021	2->1	
4-035	0->1	1->1	2->1	
4-071	5->1	
4-199	9->1	
4.1.1	 ->1	
4.2).	K->1	
4.De 	h->1	
4.Det	 ->2	
4.För	 ->1	
4.I d	e->3	
4.Jag	 ->2	
4.Kom	m->1	
4/199	9->8	
4/200	0->1	
4/55/	E->2	
4/728	/->1	
40 fr	å->1	
40 ju	r->1	
40 mi	l->1	n->1	
40 pr	o->6	
40 år	 ->1	.->1	s->1	
40(CN	S->2	
40, 4	6->1	
40/99	)->1	
400 0	0->1	
400 k	i->2	m->1	
400 m	i->2	
409 o	c->1	
4094/	1->2	
41 fr	å->1	
41 pr	o->1	
41 ri	s->1	
41 ur	v->1	
41/19	9->2	
41/99	)->1	
410 f	r->1	
42 fr	å->1	
42 i 	f->1	
42 mi	l->1	
42 oc	h->2	
43 hö	r->1	
43 om	 ->1	
43.Fr	å->1	
43.Ty	d->1	
44 - 	C->1	
44 fr	å->1	
44 oc	h->3	
44.I 	d->1	
44.Ja	g->1	
45 av	 ->1	
45 ce	n->1	
45 fr	å->1	
45 gä	l->1	
45 oc	h->1	
45, d	e->1	
45. D	ä->1	
45."I	 ->1	
45.Fr	u->1	
45.He	r->1	
45.Vi	 ->1	
45/00	 ->1	
45/20	0->1	
46 oc	h->2	
462 u	n->1	
47 gä	l->1	
48 gä	l->1	
48 i 	f->2	
48 in	n->1	
48 än	d->1	
48, 2	4->1	
48.De	t->1	
487 m	i->1	
5 (en	 ->1	
5 - 8	0->1	
5 000	 ->2	.->1	
5 008	 ->2	
5 av 	d->1	e->1	
5 cen	t->1	
5 frå	n->3	
5 gra	d->1	
5 gäl	l->2	
5 har	 ->1	
5 i A	m->1	
5 i E	G->1	
5 i f	ö->3	
5 int	e->1	
5 kom	 ->1	
5 mar	s->2	
5 mes	t->1	
5 mil	j->16	
5 min	s->1	
5 mor	d->1	
5 och	 ->4	
5 okt	o->1	
5 oli	k->2	
5 om 	d->1	m->1	
5 omr	å->1	
5 pro	c->13	j->1	
5 rik	t->1	
5 räc	k->1	
5 sep	t->1	
5 slu	t->1	
5 sta	t->1	
5 til	l->4	
5 vis	a->1	
5 år.	D->1	L->1	
5 års	 ->1	
5(CNS	)->3	
5)Utt	j->1	
5, 16	 ->1	,->1	
5, de	 ->1	
5, dä	r->1	
5, nå	g->1	
5, oc	h->2	
5, ut	o->1	
5,5 p	r->1	
5,8 m	i->1	
5-000	1->1	2->1	3->4	4->2	6->3	7->3	9->2	
5-001	0->2	1->2	2->2	8->2	
5-002	0->1	2->2	
5-004	0->1	1->1	5->2	
5-005	0->1	
5-006	9->1	
5-007	3->1	8->1	
5-008	7->1	
5-009	5->1	
5-010	4->2	5->2	6->1	7->2	8->2	
5-012	0->1	2->1	
5-016	7->1	
5-018	0->2	
5-020	8->2	
5-030	5->1	
5-032	7->2	
5-033	3->2	4->2	
5-034	1->2	
5-199	7->1	
5. Dä	r->1	
5."I 	d->1	
5.)Ju	s->1	
5.00.	)->1	F->1	
5.4 i	n->1	
5.Des	s->1	
5.Eme	l->1	
5.Fru	 ->1	
5.Frå	g->1	
5.Her	r->1	
5.Såd	a->1	
5.Vi 	i->1	
5/00 	-->1	
5/1/1	9->2	
5/199	9->4	
5/200	0->1	
5/35/	E->1	
5/95.	F->1	
5/98-	9->1	
5/99)	:->2	A->1	
5/EG 	a->1	o->1	s->1	u->1	
5/EG,	 ->2	
50 - 	C->1	
50 00	0->1	
50 gu	l->1	
50 i 	a->1	
50 mi	l->4	
50 oc	h->2	
50 pr	o->3	
50, s	k->1	
50- o	c->1	
50-ta	l->2	
50/19	9->1	
50/20	0->1	
500 0	0->1	
51/19	9->1	
519 -	 ->1	
52 - 	C->1	
52 i 	t->1	
52(CN	S->1	
52/19	9->1	
520 -	 ->1	
520 f	r->1	
522 -	 ->1	
53 pr	o->1	
540 m	i->1	
55 i 	A->1	f->2	
55 in	t->1	
55 mo	r->1	
55 pr	o->1	
55)Ut	t->1	
55/EG	 ->1	,->1	
550 -	 ->1	
56 pr	o->1	
56, s	o->1	
57 (m	e->1	
57,5 	p->1	
57.Eu	r->1	
5713/	1->1	
58 - 	C->1	
58 i 	E->1	
58).D	e->1	
58.1 	i->1	
591/E	K->2	
598 -	 ->2	
5b ka	n->1	
5b-om	r->1	
5b.De	t->1	
6 "på	p->1	
6 - C	5->1	
6 - s	a->1	
6 000	 ->1	
6 [KO	M->1	
6 dec	e->1	
6 eft	e->1	
6 ell	e->1	
6 emo	t->1	
6 frå	n->2	
6 för	 ->2	
6 gäl	l->1	
6 had	e->1	
6 har	 ->1	
6 i E	G->1	
6 i a	v->1	
6 i f	ö->6	
6 i h	ö->1	
6 i u	n->1	
6 ind	i->1	
6 kom	m->1	
6 lig	g->1	
6 låg	 ->1	
6 med	 ->1	
6 mil	j->1	
6 nov	e->1	
6 och	 ->15	
6 om 	a->1	
6 per	s->1	
6 pro	c->6	
6 rad	e->1	
6 så 	s->1	
6 tas	 ->1	
6 tot	a->1	
6 var	 ->1	
6 vil	k->1	
6 är 	s->1	
6 års	 ->2	
6 åte	r->1	
6(COD	)->2	
6) sa	m->1	
6, 20	,->1	
6, 38	,->1	
6, 7,	 ->1	
6, fö	r->1	
6, ha	r->1	
6, me	n->1	
6, nä	r->1	
6, so	m->3	
6, ta	r->1	
6, vi	l->1	
6,07 	m->1	
6.Det	 ->3	
6.Enl	i->2	
6.Frå	g->1	
6.Her	r->1	
6.Jag	 ->3	
6.Man	 ->1	
6.Men	 ->1	
6.Och	 ->1	
6.Så 	s->1	
6.Tac	k->1	
6.År 	1->1	
6/00)	 ->1	:->1	
6/199	9->1	
6/200	0->2	
6/35/	E->3	
6/71 	a->1	
6/71/	E->1	
6/99)	:->2	
60 00	0->1	
60 fr	å->1	
60-ta	l->1	
60/92	 ->1	
60/99	 ->1	
600 b	i->1	
614/1	9->1	
62 - 	C->1	
62 eu	r->1	
62 i 	f->1	
62 un	d->1	
62 up	p->1	
62.Ma	n->1	
64 rö	s->1	
652 -	 ->1	
66 - 	C->1	
66 em	o->1	
662 -	 ->1	
67 00	0->1	
67 ha	r->1	
67 i 	A->1	u->1	
67 me	d->1	
67 mi	l->3	
67 oc	h->2	
67, o	c->1	
67/19	9->1	
68 at	t->1	
685/9	5->1	
69 oc	h->1	
69(CO	D->2	
69/19	9->1	
7 (av	s->1	
7 (me	r->1	
7 - d	v->1	
7 - i	n->2	
7 000	 ->1	
7 dec	e->4	
7 där	 ->1	
7 fal	l->1	
7 frå	n->1	
7 för	e->1	t->1	
7 gra	d->1	
7 gäl	l->1	
7 har	 ->2	
7 här	r->1	
7 i A	m->3	
7 i a	r->1	v->1	
7 i b	e->1	
7 i d	e->1	
7 i f	ö->3	
7 i u	t->1	
7 i v	i->1	
7 led	a->1	
7 lyd	e->1	
7 län	d->1	
7 med	a->1	
7 mil	j->7	
7 näm	n->1	
7 och	 ->11	
7 okt	o->1	
7 om 	t->1	
7 pro	c->5	
7 på 	R->1	n->1	
7 så 	s->1	
7 tro	l->1	t->1	
7 upp	,->1	
7 är 	i->1	
7 års	 ->1	
7(COS	)->1	
7) 06	5->1	
7).. 	(->1	
7, 18	,->1	
7, 34	,->1	
7, 42	 ->2	
7, 88	 ->1	
7, 9,	 ->1	
7, dv	s->1	
7, me	n->1	
7, oc	h->2	
7, om	 ->1	
7, re	s->1	
7, so	m->1	
7, så	 ->1	
7, va	r->1	
7,2 m	i->1	
7,42 	m->1	
7,5 p	r->1	
7.- D	e->1	
7.. (	E->1	
7.1 i	 ->1	
7.2 i	 ->2	
7.30,	 ->1	
7.Bet	ä->1	
7.Det	 ->2	
7.Eur	o->1	
7.Frå	g->1	
7.I v	å->1	
7.Man	 ->1	
7.Nu 	ä->1	
7.Sed	a->1	
7.Slu	t->1	
7.Vi 	h->1	m->1	
7/019	4->2	
7/035	2->1	
7/037	0->2	1->2	
7/199	9->6	
7/200	0->3	
7/60/	9->1	
7/99 	(->1	
7/99)	:->2	
70 an	s->1	
70 mi	l->2	
70 pr	o->1	
70(CO	D->2	
700 a	r->1	
700 h	a->1	
700 o	c->2	
71 an	g->1	
71(CO	D->2	
71/EG	 ->1	
713/1	9->1	
715/9	8->1	
728/E	G->1	
73,9 	p->1	
73/19	9->1	
74 tu	s->1	
75 - 	8->1	
75 mi	l->2	
75 om	 ->1	
76 el	l->1	
76 pr	o->1	
762 u	p->1	
762.M	a->1	
77 - 	i->1	
77 mi	l->1	
778/9	9->1	
78/19	9->1	
78/99	)->1	
780/9	9->1	
781/9	9->1	
782/9	9->1	
785/9	9->1	
786/9	9->1	
788/9	9->1	
79/40	9->1	
791/9	9->1	
793/9	9->1	
795/9	9->1	
796/9	9->1	
798/9	9->1	
7?De 	p->1	
7Näst	a->1	
8 - 1	9->1	
8 - C	5->3	
8 462	 ->1	
8 att	 ->1	
8 beh	ö->1	
8 dec	e->1	
8 frå	n->3	
8 för	e->1	
8 god	k->1	
8 gäl	l->1	
8 had	e->1	
8 hän	v->1	
8 i E	G->1	K->1	
8 i b	e->1	
8 i d	i->1	
8 i f	ö->2	
8 inn	e->1	
8 jul	i->1	
8 kos	t->1	
8 mil	j->6	
8 mån	a->1	
8 nov	e->3	
8 nya	 ->1	
8 och	 ->12	
8 pro	c->1	
8 reg	i->1	
8 res	o->1	
8 ska	l->1	
8 til	l->2	
8 ton	 ->1	,->1	
8 und	e->1	
8 utb	e->1	
8 utg	ö->1	
8 var	 ->2	
8 änd	r->1	
8 är 	g->1	i->1	k->1	r->1	
8(CNS	)->1	
8(SYN	)->1	
8) 51	9->1	
8) 52	0->1	2->1	
8).De	t->1	
8)066	2->1	
8, 24	5->1	
8, 27	,->1	
8, 30	,->1	
8, 32	,->1	
8, 44	 ->1	
8, 9,	 ->1	
8, SE	K->2	
8, dä	r->1	
8, så	v->1	
8-200	2->2	
8-98/	0->1	
8. De	s->1	
8.1 i	 ->1	
8.4.D	e->1	
8.Det	 ->1	
8.Pre	c->1	
8.Sto	r->1	
8/010	6->2	
8/016	9->2	
8/031	8->1	
8/199	9->5	
8/200	0->2	
8/591	/->2	
8/98 	-->1	
8/99)	:->4	
8/EG,	 ->1	
80 en	s->1	
80 i 	f->4	
80 mi	l->1	
80 pr	o->11	
80 än	d->1	
80 åt	g->1	
80.4.	F->1	
80/19	9->2	
80/99	)->1	
801/9	9->1	
803(C	N->1	
805(C	N->1	
805/9	9->1	
807/9	9->1	
808/9	9->1	
8095/	1->2	
81 oc	h->5	
81 pr	o->1	
81.1 	d->1	o->2	
81.1.	F->1	V->1	
81.3 	E->1	b->1	i->1	
81.3,	 ->1	
81.3;	 ->1	
81/99	)->1	
813/9	9->1	
817/9	9->1	
819/9	9->1	
82 ha	r->1	
82 in	n->1	
82) f	ö->1	
82, d	e->1	
82, e	l->1	
82, f	r->1	
82, l	ä->1	
82, t	i->1	
82.I 	e->1	
82.Is	r->1	
82/99	)->1	
825(C	N->2	
829/9	9->1	
83 (C	O->1	
83 pr	o->1	
85 oc	h->2	
85 pr	o->1	
85 ti	l->1	
85/95	.->1	
85/99	)->1	
86 ha	d->1	
86 i 	E->1	f->1	
86 oc	h->1	
86 pr	o->1	
86.År	 ->1	
86/99	)->1	
87 mi	l->1	
87, 8	8->1	
87.1 	i->1	
87.2 	i->1	
87/19	9->1	
88 i 	E->1	
88 oc	h->1	
88 är	 ->1	
88/59	1->2	
88/99	)->1	
89 i 	f->1	
89 ti	l->1	
89, 1	9->1	
8: fo	r->1	
8:e å	r->1	
9 (Ho	w->1	
9 - 1	9->20	
9 - 3	1->1	
9 - C	4->1	5->6	
9 ant	o->3	
9 avs	a->1	
9 bet	y->1	
9 dec	e->1	
9 dep	a->1	
9 där	 ->1	
9 död	a->1	
9 erh	ö->1	
9 fal	l->1	
9 feb	r->1	
9 fra	m->2	
9 frå	n->3	
9 god	k->1	
9 had	e->1	
9 ham	n->1	
9 har	 ->3	
9 i M	a->1	
9 i f	ö->1	
9 i h	a->1	
9 i s	t->1	
9 i v	a->1	
9 inn	e->1	
9 int	e->1	
9 jäm	n->1	
9 kan	 ->1	
9 kom	m->2	
9 kun	d->1	
9 län	d->1	
9 mar	s->1	
9 mil	j->3	
9 min	u->1	
9 när	 ->1	
9 och	 ->6	
9 ock	s->1	
9 om 	a->1	
9 pro	c->3	
9 prä	g->1	
9 ras	a->1	
9 ska	l->1	
9 som	 ->1	
9 til	l->2	
9 upp	g->1	m->1	
9 ut 	e->1	
9 var	 ->2	
9 vis	a->1	
9 är 	o->1	
9 äve	n->1	
9 års	 ->1	
9 öve	r->1	
9".Bå	d->1	
9(COD	)->2	
9) 01	1->1	
9) 05	5->1	
9) 15	8->1	
9) 34	4->1	
9) av	 ->12	
9) fr	å->2	
9) oc	h->1	
9).Ko	m->1	
9)000	3->2	
9)006	6->1	
9)059	8->2	
9):An	g->18	
9)Ang	å->2	
9, 19	9->1	
9, 31	 ->1	
9, 40	,->1	
9, an	d->1	
9, av	 ->1	
9, be	s->1	
9, dv	s->1	
9, fö	r->1	
9, ha	r->1	
9, nä	r->1	
9, oc	h->2	
9-200	4->1	6->1	
9. Vi	 ->1	
9..(F	R->1	
9.1 v	i->1	
9.2 i	 ->2	
9.50 	o->1	
9.De 	l->1	
9.Des	s->1	
9.Det	 ->1	
9.En 	r->1	
9.Eur	o->1	
9.Frå	n->1	
9.För	u->1	ä->1	
9.Jag	 ->2	
9.Kom	m->1	
9.Und	e->1	
9.Vi 	m->1	
9/001	2->1	3->1	
9/008	3->1	
9/009	0->1	
9/022	8->1	
9/024	0->2	
9/080	3->1	5->1	
9/082	5->2	
9/199	9->1	
9/200	0->2	
9/212	3->1	7->1	
9/409	 ->1	
9/99)	:->2	
90 de	t->1	
90 dö	d->1	
90 pr	o->4	
90 ut	a->1	
90(CO	D->1	
90-ta	l->1	
90.De	t->1	
91 ef	t->1	
91 ge	r->1	
91 oc	h->1	
91 pr	o->1	
91/99	)->1	
91/EK	S->2	
917 o	c->1	
92 oc	h->1	
92 sk	r->1	
92 so	m->1	
92 år	s->1	
92, e	n->1	
92/43	.->1	
923, 	e->1	
93 ha	r->1	
93 oc	h->2	
93 pe	r->1	
93 ut	e->1	
93, 1	9->1	
93-19	9->2	
93.Om	 ->1	
93/75	 ->1	
93/99	)->1	
930-t	a->1	
93?Fr	å->1	
94 et	t->1	
94 ha	r->1	
94 nä	r->1	
94 oc	h->2	
94 pr	o->2	
94(CO	D->2	
94, f	ö->1	
94, k	o->1	
94-19	9->1	
94.De	t->1	
94/19	9->2	
94/55	/->2	
94/72	8->1	
945.F	r->1	
948.D	e->1	
95 (e	n->1	
95 ha	r->1	
95 i 	f->1	
95 ko	m->1	
95 mi	l->3	
95 ri	k->1	
95 sl	u->1	
95 ti	l->1	
95 år	s->1	
95, n	å->1	
95, o	c->1	
95-19	9->1	
95.Fr	å->1	
95/1/	1->2	
95/19	9->1	
95/35	/->1	
95/99	)->1	
957 (	m->1	
957.E	u->1	
96 - 	s->1	
96 ef	t->1	
96 ha	r->1	
96 i 	h->1	
96 lå	g->1	
96 oc	h->1	
96 va	r->1	
96 vi	l->1	
96 är	 ->1	
96 år	s->2	
96, h	a->1	
96, v	i->1	
96.De	t->1	
96.En	l->1	
96.Ja	g->1	
96.Me	n->1	
96.Oc	h->1	
96/35	/->3	
96/71	 ->1	/->1	
96/99	)->1	
9614/	1->1	
967 h	a->1	
967 i	 ->1	
967 m	e->1	
967 o	c->2	
967, 	o->1	
969 o	c->1	
97 (a	v->1	
97 - 	i->1	
97 dä	r->1	
97 fö	r->1	
97 ha	r->1	
97 hä	r->1	
97 i 	a->1	
97 ly	d->1	
97 oc	h->5	
97 om	 ->1	
97 på	 ->1	
97 tr	o->2	
97 up	p->1	
97 är	 ->1	
97 år	s->1	
97) 0	6->1	
97, m	e->1	
97, v	a->1	
97.- 	D->1	
97.. 	(->1	
97.Be	t->1	
97.De	t->2	
97.I 	v->1	
97.Ma	n->1	
97.Nu	 ->1	
97.Se	d->1	
97.Vi	 ->2	
97/01	9->2	
97/03	5->1	7->4	
97/99	 ->1	
976 e	l->1	
977 -	 ->1	
97?De	 ->1	
97Näs	t->1	
98 - 	1->1	C->2	
98 go	d->1	
98 ha	d->1	
98 ko	s->1	
98 mi	l->1	
98 oc	h->6	
98 re	g->1	
98 sk	a->1	
98 un	d->1	
98 ut	b->1	g->1	
98 va	r->2	
98 är	 ->2	
98) 5	1->1	2->2	
98)06	6->1	
98, S	E->2	
98, d	ä->1	
98-20	0->2	
98-98	/->1	
98. D	e->1	
98.Pr	e->1	
98.St	o->1	
98/01	0->2	6->2	
98/03	1->1	
98/99	)->1	
982, 	d->1	
982.I	s->1	
986 h	a->1	
986 o	c->1	
986.Å	r->1	
989, 	1->1	
99 (H	o->1	
99 - 	1->20	3->1	C->6	
99 an	t->3	
99 av	s->1	
99 be	t->1	
99 dä	r->1	
99 er	h->1	
99 fr	a->2	
99 go	d->1	
99 ha	d->1	m->1	r->3	
99 i 	h->1	s->1	v->1	
99 in	n->1	
99 jä	m->1	
99 ka	n->1	
99 ko	m->2	
99 ku	n->1	
99 nä	r->1	
99 oc	h->4	k->1	
99 om	 ->1	
99 pr	ä->1	
99 ra	s->1	
99 sk	a->1	
99 ti	l->1	
99 up	p->2	
99 ut	 ->1	
99 va	r->2	
99 vi	s->1	
99 äv	e->1	
99 år	s->1	
99 öv	e->1	
99".B	å->1	
99) 0	1->1	5->1	
99) 1	5->1	
99) 3	4->1	
99) a	v->12	
99) f	r->2	
99) o	c->1	
99).K	o->1	
99)00	0->2	6->1	
99)05	9->2	
99):A	n->18	
99)An	g->2	
99, a	v->1	
99, b	e->1	
99, d	v->1	
99, h	a->1	
99, n	ä->1	
99, o	c->2	
99-20	0->2	
99. V	i->1	
99..(	F->1	
99.2 	i->2	
99.De	 ->1	s->1	t->1	
99.En	 ->1	
99.Eu	r->1	
99.Fr	å->1	
99.Fö	r->2	
99.Ja	g->2	
99.Ko	m->1	
99.Un	d->1	
99.Vi	 ->1	
99/00	1->2	8->1	9->1	
99/02	2->1	4->2	
99/08	0->2	2->2	
99/21	2->2	
990 u	t->1	
990.D	e->1	
991 e	f->1	
991 g	e->1	
991 o	c->1	
992 s	k->1	o->1	
992 å	r->1	
992, 	e->1	
993 h	a->1	
993 o	c->1	
993 u	t->1	
993, 	1->1	
993-1	9->2	
993.O	m->1	
993?F	r->1	
994 e	t->1	
994 h	a->1	
994 o	c->2	
994, 	f->1	
994-1	9->1	
995 (	e->1	
995 h	a->1	
995 k	o->1	
995 r	i->1	
995 s	l->1	
995 å	r->1	
995, 	n->1	o->1	
995-1	9->1	
996 -	 ->1	
996 e	f->1	
996 h	a->1	
996 i	 ->1	
996 l	å->1	
996 o	c->1	
996 v	a->1	i->1	
996 ä	r->1	
996 å	r->2	
996, 	h->1	v->1	
996.D	e->1	
996.E	n->1	
996.J	a->1	
996.M	e->1	
996.O	c->1	
997 (	a->1	
997 -	 ->1	
997 d	ä->1	
997 f	ö->1	
997 h	a->1	ä->1	
997 i	 ->1	
997 l	y->1	
997 o	c->5	m->1	
997 p	å->1	
997 t	r->2	
997 u	p->1	
997 ä	r->1	
997 å	r->1	
997) 	0->1	
997, 	m->1	v->1	
997.-	 ->1	
997..	 ->1	
997.B	e->1	
997.D	e->2	
997.I	 ->1	
997.M	a->1	
997.N	u->1	
997.V	i->2	
997/0	1->2	3->5	
997?D	e->1	
997Nä	s->1	
998 g	o->1	
998 h	a->1	
998 k	o->1	
998 o	c->6	
998 r	e->1	
998 s	k->1	
998 u	n->1	t->2	
998 v	a->2	
998 ä	r->2	
998) 	5->3	
998, 	S->2	d->1	
998-2	0->2	
998. 	D->1	
998.P	r->1	
998.S	t->1	
998/0	1->4	
999 -	 ->26	
999 a	n->3	v->1	
999 d	ä->1	
999 e	r->1	
999 f	r->2	
999 g	o->1	
999 h	a->5	
999 i	 ->3	n->1	
999 j	ä->1	
999 k	a->1	o->2	u->1	
999 n	ä->1	
999 o	c->3	m->1	
999 p	r->1	
999 r	a->1	
999 s	k->1	
999 t	i->1	
999 u	p->2	t->1	
999 v	a->2	i->1	
999 ä	v->1	
999 å	r->1	
999 ö	v->1	
999".	B->1	
999) 	0->2	1->1	3->1	a->12	f->1	
999).	K->1	
999)0	0->2	5->1	
999, 	a->1	b->1	d->1	h->1	n->1	o->2	
999-2	0->2	
999. 	V->1	
999..	(->1	
999.D	e->3	
999.E	n->1	u->1	
999.F	r->1	ö->2	
999.J	a->1	
999.K	o->1	
999.U	n->1	
999.V	i->1	
999/0	0->4	2->3	8->4	
999/2	1->2	
999: 	"->1	
99: "	j->1	
9: "j	a->1	
: "At	t->1	
: "De	t->4	
: "Ja	,->1	
: "Mi	n->1	
: "Om	 ->1	
: "al	d->1	
: "de	t->1	
: "he	l->1	
: "in	 ->1	
: "ja	 ->1	
: "va	r->1	
: Anl	ä->1	
: Anm	ä->1	
: Arb	e->1	
: Art	i->1	
: Ast	u->1	
: Att	 ->1	
: De 	d->1	n->1	s->1	
: Des	s->1	
: Det	 ->4	t->1	
: Eft	e->1	
: Eri	k->1	
: Eur	o->1	
: Fin	n->1	
: Fir	m->1	
: Flo	r->1	
: Fri	h->2	
: Frä	m->1	
: För	 ->2	h->1	s->2	
: Gem	e->1	
: Gen	o->1	
: Gre	k->1	
: Ham	b->1	
: Han	d->1	
: Hol	z->1	
: I b	ö->1	
: I m	o->1	
: I s	l->1	
: Ing	e->1	
: Jag	 ->7	
: Jor	d->1	
: Koc	h->1	
: Kom	m->4	
: Kon	v->1	
: Kän	n->1	
: Kär	n->1	
: Mai	n->1	
: Nar	k->1	
: Nyt	t->1	
: När	 ->3	
: Om 	E->1	
: Osl	o->1	
: Par	l->1	
: Por	t->1	
: På 	g->1	
: Rev	i->1	
: Sta	d->1	
: Stö	d->1	
: Tur	k->1	
: Tåg	k->1	
: Und	e->1	
: Uni	o->1	
: Utn	ä->1	
: Utv	ä->1	
: Vad	 ->3	
: Vap	e->1	
: Vem	 ->3	
: Vi 	b->1	f->2	h->1	m->2	ä->1	
: ang	i->1	
: ant	i->3	
: att	 ->8	
: bal	a->1	
: bes	t->1	
: de 	h->1	s->1	
: def	i->1	
: del	s->1	
: den	 ->7	n->1	
: det	 ->9	t->4	
: dir	e->1	
: dub	b->1	
: där	i->1	
: en 	e->1	f->2	l->1	m->1	r->1	s->1	t->1	
: ett	 ->2	
: for	d->1	s->1	
: frå	g->2	
: för	 ->9	e->1	s->2	
: gem	e->1	
: gen	o->1	
: gör	 ->1	
: han	d->1	s->1	
: hur	 ->4	
: hög	s->1	
: i F	r->1	
: i l	e->1	
: i r	e->1	
: ino	m->1	
: ins	p->1	t->1	
: ja,	 ->1	
: jag	 ->4	
: kan	d->1	
: kom	m->3	
: man	 ->1	
: med	 ->1	l->1	
: min	i->1	
: nu 	s->1	
: när	 ->1	,->1	
: om 	E->1	e->1	k->1	r->1	
: ope	r->1	
: par	a->1	
: pro	g->1	
: rät	t->1	
: ska	l->1	
: sys	t->1	
: tan	k->1	
: til	l->1	
: tol	k->1	
: und	e->1	
: upp	b->1	
: utb	y->2	
: utn	y->1	
: utv	i->1	
: vad	 ->2	
: var	f->2	k->1	
: vem	 ->3	
: vi 	h->2	k->1	l->1	m->1	s->3	v->2	
: vil	k->2	
: våg	a->1	
: vår	t->1	
: Är 	k->1	
: Äve	n->1	
: Åtg	ä->2	
: Öpp	e->1	
: å e	n->1	
: öns	k->1	
:Angå	e->19	
:Den 	s->1	
:Det 	e->1	
:För 	d->1	
:Föro	r->1	
:a år	h->1	
:e ra	p->2	
:e år	s->1	
:s (f	i->1	
:s Ba	r->1	
:s Eu	r->1	
:s an	s->1	
:s ar	b->2	g->1	
:s be	f->1	s->2	
:s bi	l->1	s->1	
:s bu	d->2	
:s by	r->1	
:s de	l->1	
:s di	r->1	
:s do	g->1	
:s eg	e->1	
:s ek	o->1	
:s eu	r->1	
:s fr	a->2	
:s fö	r->2	
:s ga	r->1	
:s ge	m->1	
:s gi	v->1	
:s ha	m->1	
:s he	l->1	
:s in	g->1	s->5	
:s ko	n->1	
:s ku	s->1	
:s la	g->1	
:s li	v->2	
:s me	d->3	
:s mi	l->1	n->1	
:s nu	v->1	
:s nä	s->1	
:s oc	h->3	
:s om	r->1	
:s or	d->1	g->1	
:s pa	r->1	
:s po	l->3	
:s re	g->1	s->1	
:s sa	k->1	
:s si	d->1	
:s st	r->4	y->1	
:s sä	k->1	
:s te	r->1	
:s tj	ä->1	
:s up	p->1	
:s ur	s->1	
:s ut	r->1	
:s ve	r->1	
:s.Le	d->1	
; Dan	m->1	
; Jav	e->1	
; all	a->1	
; ann	a->1	
; ant	i->1	
; art	i->1	
; att	 ->3	
; av 	k->1	
; b) 	m->1	
; de 	ä->1	
; den	 ->4	
; des	s->4	
; det	 ->21	t->1	
; där	 ->1	
; då 	b->1	
; en 	a->1	d->1	k->1	s->2	
; end	a->1	
; enl	i->1	
; fis	k->1	
; for	t->1	
; fri	h->1	
; för	 ->4	b->1	o->1	u->1	
; här	 ->1	
; i F	ö->1	
; i d	a->1	
; i e	g->1	
; inf	o->1	
; inl	e->1	
; ins	y->1	
; int	e->1	
; jag	 ->4	
; kom	m->1	
; loj	a->1	
; man	 ->1	
; men	 ->2	
; min	 ->1	a->1	
; och	 ->5	
; pun	k->3	
; sam	h->1	
; sko	g->1	
; slu	t->1	
; und	a->1	
; vi 	b->1	f->1	h->2	m->1	
; vid	 ->1	
; änn	u->1	
; å e	n->1	
; öve	r->1	
? 21 	å->1	
? Den	 ->2	
? Har	 ->2	
? Int	e->1	
? Med	 ->1	
? Och	:->1	
? Råd	e->1	
?"Ja 	E->1	
?, rå	d->2	
?- (P	T->3	
?. (E	N->8	
?. (F	R->1	
?.(EN	)->2	
?.Her	r->2	
?Anse	r->3	
?Ansl	a->1	
?Att 	d->1	h->1	
?Av t	r->1	
?Avsl	u->1	
?Bord	e->1	
?Dage	n->1	
?De h	a->1	
?De p	r->1	
?De t	y->1	
?Den 	2->1	a->1	f->2	k->1	s->3	
?Dess	a->1	
?Det 	b->2	d->1	e->1	f->2	h->1	k->2	ä->9	
?Dett	a->1	
?Där 	h->1	
?Därf	ö->2	
?Efte	r->1	
?Elle	r->1	
?Enda	s->1	
?Enli	g->1	
?Ett 	E->1	e->1	s->1	
?Euro	p->2	
?Finn	s->1	
?Folk	 ->1	
?Fru 	l->1	t->5	
?Fråg	a->3	
?För 	a->1	d->4	e->1	o->1	
?Förs	t->1	
?Har 	o->1	r->1	v->2	
?Heml	i->1	
?Herr	 ->15	
?Hur 	b->1	k->2	l->1	m->2	s->2	t->1	ä->1	
?Här 	ä->1	
?Härm	e->1	
?I Fr	a->1	
?I da	g->2	
?I er	a->1	
?I fj	o->1	
?I me	d->1	
?I så	 ->1	
?I vi	l->1	
?Init	i->1	
?Inte	 ->1	
?Ja, 	h->1	n->1	
?Jag 	a->1	f->1	j->1	k->1	r->2	s->3	t->3	v->6	ö->3	
?Jo d	å->1	
?Jo, 	d->1	i->1	s->1	
?Kan 	k->1	u->1	
?Kans	k->3	
?Koll	e->1	
?Komm	e->4	i->2	
?Kära	 ->1	
?Man 	f->1	
?Men 	p->1	v->1	
?Mena	r->1	
?Natu	r->1	
?Nej,	 ->5	
?Nej.	I->1	
?Ni k	o->2	
?Ni n	ä->1	
?När 	d->1	k->1	t->1	
?Näst	a->1	
?Och 	j->1	o->1	s->1	
?Olik	a->1	
?Om i	n->2	
?Parl	a->1	
?Prob	l->1	
?På d	e->1	
?På v	i->1	
?RINA	 ->1	
?Rege	r->1	
?Seda	n->1	
?Seri	ö->1	
?Skul	l->3	
?Som 	p->1	s->1	
?Svar	e->1	
?Tack	 ->1	
?Till	 ->1	
?Tyck	e->1	
?Tänk	 ->1	
?Utgi	f->1	
?Vad 	b->1	f->1	g->1	k->1	s->1	t->2	
?Vem 	d->1	k->1	
?Vets	k->1	
?Vi b	e->2	
?Vi f	å->1	
?Vi h	a->1	
?Vi m	å->2	
?Vi s	e->1	v->1	
?Vi t	r->1	
?Vi ä	r->2	
?Vilk	a->6	e->7	
?Viss	a->2	
?Är d	e->8	
?Är h	y->1	
?Är i	n->1	
?Är v	i->1	
?Även	 ->2	
A - o	c->1	
A OCH	 ->1	
A att	 ->1	
A ell	e->1	
A har	 ->3	
A på 	b->1	
A var	 ->1	
A) De	 ->1	
A) Ve	n->1	
A, Ka	n->1	
A, ef	t->1	
A, so	m->1	
A-ins	t->1	
A-stö	d->1	
A. Gu	t->1	
A.Jag	 ->1	
A.Vi 	s->1	
A5-00	0->13	1->8	2->2	6->1	7->2	8->1	
A5-01	0->9	
A:s.L	e->1	
ABB A	l->1	
ABB-A	l->2	
ABC d	e->1	
ADR) 	o->1	
AF gö	r->1	
AF i 	e->1	r->1	
AF ka	n->1	
AF ko	n->1	
AF sk	a->1	
AF, E	u->1	
AF, d	e->1	
AF, e	n->1	
AF, k	o->1	
AF, s	å->2	
AF, v	i->1	
AF, ö	v->1	
AF.Al	l->1	
AF.Fö	r->1	
AF.He	r->1	
AF.Me	n->1	
AF:s 	(->1	u->1	
AKTUE	L->1	
ANDE 	F->1	
ARPOL	 ->1	
AS (I	n->1	
ASP m	å->1	
ATT O	M->1	
Accep	t->1	
Act. 	D->1	
Adana	 ->1	
Adena	u->1	
Adolf	 ->2	
Adria	t->1	
Afrik	a->4	
Agrif	i->1	
Agust	a->1	
Ahern	 ->5	,->3	
Aids,	 ->1	
Akkuy	u->2	
Akköy	 ->1	
Aktiv	i->1	
Alava	n->2	
Albac	è->1	
Alban	i->1	
Alber	t->1	
Albri	g->1	
Aldri	g->1	
Alexa	n->2	
Alger	i->1	
Alica	n->1	
Alla 	a->1	b->3	d->5	g->2	h->4	i->2	l->1	m->1	s->2	t->1	u->1	v->2	
Allde	l->1	
Allmä	n->4	
Allt 	d->11	f->2	s->2	t->1	
Alltf	ö->1	
Allts	e->2	å->2	
Alper	n->1	
Alpes	 ->1	
Alsac	e->3	
Alsth	o->3	
Alten	e->18	
Ameri	k->2	
Amoco	,->1	
Amoko	 ->5	
Amos 	O->1	
Amste	r->39	
Andra	 ->4	b->3	
Angel	i->1	
Angåe	n->22	
Anhål	l->1	
Ankar	a->1	
Anled	n->1	
Anläg	g->1	
Anmäl	n->1	
Anna 	T->1	
Annar	s->4	
Anser	 ->4	
Ansla	g->1	
Ansva	r->4	
Antal	e->2	
Antón	i->1	
Anver	s->1	
Använ	d->1	
Apari	c->1	
Applå	d->5	
Arabr	e->1	
Arabv	ä->1	
Arafa	t->1	
Arbet	s->4	
Arden	n->1	
Ari V	a->1	
Arian	e->3	
Artik	e->2	l->1	
Asien	 ->1	,->1	
Assad	 ->1	,->1	
Astur	i->1	
Atatu	r->1	
Atatü	r->1	
Atlan	t->4	
Att F	l->1	
Att a	v->1	
Att b	i->1	
Att d	e->3	ö->1	
Att f	r->1	
Att g	a->1	e->2	
Att h	j->1	u->1	
Att i	 ->1	n->1	
Att k	u->1	
Att l	å->2	
Att m	a->2	
Att r	a->1	
Att s	å->1	
Att t	a->1	i->1	
Att u	t->3	
Att v	i->1	
Attac	k->1	
Ausch	w->1	
Auto/	O->1	
Auver	g->1	
Av 41	0->1	
Av al	l->4	
Av av	g->1	
Av be	s->1	t->1	
Av de	n->11	t->4	
Av en	 ->1	
Av om	f->1	
Av sa	m->2	
Av tr	e->1	
Av vi	l->1	s->1	
Avbro	t->1	
Avfal	l->1	
Avgån	g->1	
Avian	o->1	
Avsat	t->1	
Avser	 ->1	
Avsev	ä->1	
Avslu	t->14	
Azore	r->2	
B Als	t->1	
B och	 ->1	
B ta 	u->1	
B-Als	t->2	
B5-00	0->2	4->2	
BATT 	O->1	
BB Al	s->1	
BB-Al	s->2	
BC de	n->1	
BI - 	d->1	
BNI b	e->1	
BNI i	 ->1	
BNI o	c->2	
BNI p	e->2	
BNI, 	e->1	
BNP j	ä->1	
BNP m	i->1	
BNP p	e->3	å->1	
BNP å	r->1	
BNP, 	i->1	m->1	
BP, e	f->1	
BRÅDS	K->1	
BSE o	c->2	
BSE-k	r->3	
BSE-t	e->1	
Bakom	 ->2	
Balfo	r->1	
Balka	n->7	
Bank 	e->1	
Bara 	g->1	m->1	n->1	s->1	
Barak	 ->5	.->1	s->3	
Barce	l->2	
Baren	t->1	
Barnh	i->1	
Barni	e->14	
Barón	 ->2	
Baski	e->2	
Basse	-->1	
Bedrä	g->2	
Bedöm	n->2	
Befor	d->1	
Behre	n->7	
Bekvä	m->1	
Belgi	e->9	
Benel	u->1	
Beren	d->12	g->2	
Berg 	g->1	
Berge	r->12	
Berli	n->7	
Berna	r->1	
Bernd	 ->3	
Berni	é->1	
Beroe	n->1	
Berth	u->1	
Berti	n->1	
Beslu	t->4	
Besqu	e->1	
Beträ	f->7	
Betän	k->25	
Bevis	e->1	
Big b	r->1	
Bilin	d->1	
Billo	b->2	
Bilti	l->2	
Bisca	y->6	
Bistå	n->1	
Blak 	s->1	
Bland	 ->8	
Blok 	o->1	
Boett	i->1	
Bolke	s->1	
Bonde	 ->1	
Borde	 ->3	a->1	
Borto	m->1	
Bosät	t->1	
Bourl	a->6	
Bowe.	E->1	V->1	
Bowis	 ->2	
Brand	e->2	
Brasi	l->1	
Brave	r->1	
Breme	n->1	
Breta	g->8	
Brist	 ->2	e->1	
Briti	s->1	
Britt	i->1	
Brok 	d->1	f->2	g->1	o->1	s->1	
Brok,	 ->3	
Bruno	 ->1	
Bryss	e->19	
Budap	e->1	
Budge	t->1	
Bulga	r->1	
Bush,	 ->1	
Busqu	i->1	
Bygge	t->1	
Byrne	 ->1	,->1	
Byrån	 ->1	
Bästa	 ->1	
Båda 	d->1	f->1	g->1	h->1	p->1	
C den	 ->1	
C, at	t->1	
C-lek	s->1	
C. De	t->1	
C. Ef	t->1	
C.Vi 	d->1	
C4-00	1->1	
C4-02	1->1	
C4-03	5->3	
C4-07	1->1	
C5-00	0->1	2->1	4->2	5->1	9->1	
C5-01	2->2	6->1	8->2	
C5-02	0->2	
C5-03	0->1	2->2	3->4	4->2	
CAF:s	 ->1	
CECAF	:->1	
CEN e	l->1	
CEN h	a->1	
CEN k	o->1	
CEN o	c->1	
CEN) 	i->1	s->1	
CEN, 	a->1	s->1	
CEN:s	 ->4	
CERN)	 ->1	
CES) 	ä->1	
CES-z	o->3	
CH BR	Å->1	
CHO i	 ->1	
CHO, 	a->1	
CHO.D	e->1	
CK nu	 ->1	
CLAF 	s->1	
CM.At	t->1	
CNS))	 ->1	(->4	.->2	F->1	o->1	
COD))	 ->4	(->4	.->3	H->1	
COD)]	.->1	
COS)]	.->2	
CSU-g	r->1	
CSU:s	 ->2	
Cadiz	 ->3	,->1	-->1	
Cadou	 ->1	
Camre	 ->1	
Camus	 ->1	
Canad	a->1	
Candu	t->1	
Canyo	n->3	
Carpe	g->1	
Carth	y->1	
Casab	l->1	
Casac	a->1	
Caudr	o->1	
Caval	e->1	
Centr	a->13	
Cermi	s->1	
Ceyhu	n->1	
Champ	a->1	
Chiqu	i->1	
Claud	e->1	
Clint	o->1	
Coca 	C->1	
Cocil	o->1	
Cola,	 ->1	
Conak	r->1	
Const	a->1	
Corbe	t->1	
Corpu	s->1	
Costa	 ->7	,->2	
Counc	i->1	
Cox o	c->1	
Cox s	a->1	
Cox!J	a->1	
Cox, 	j->1	
Cresp	o->2	
Cunha	s->1	
Curie	-->1	
Cusí 	ä->1	
Cuxha	v->1	
Cyper	n->1	
D bör	 ->1	
D för	 ->1	
D krä	v->1	
D)) (	U->1	f->1	
D)) i	n->2	
D))(P	a->4	
D))..	 ->1	(->1	
D)).F	r->1	
D))He	r->1	
D)].)	 ->1	
D, oc	h->1	
D-gru	p->2	
DA) D	e->1	
DA) V	e->1	
DD, o	c->1	
DD-gr	u->2	
DDR.S	e->1	
DE FR	Å->1	
DE) H	e->1	
DE) J	a->1	
DE) Ä	r->1	
DE).(	E->1	
DE- o	c->2	
DE-gr	u->4	
DE-le	d->1	
DEBAT	T->1	
DR an	s->1	
DR) o	c->1	
DR-gr	u->1	
DR.Se	d->1	
DR:s 	u->1	
DSKAN	D->1	
Da Co	s->3	
Dagen	s->5	
Dagli	g->2	
Dagma	r->1	
Dalai	 ->7	
Dam b	e->1	
Dam s	a->1	
Damas	k->1	
Danma	r->26	
Darms	t->1	
David	 ->3	
De 14	 ->1	
De 15	 ->1	
De Gr	ö->1	
De Pa	l->1	
De Ro	o->1	
De ak	t->1	
De al	l->2	
De an	d->2	s->1	t->1	
De av	 ->1	
De be	d->1	h->2	r->1	
De bi	l->1	
De da	n->2	
De di	s->2	
De dr	ö->1	
De eu	r->2	
De fa	r->1	t->1	
De fi	c->1	n->1	
De fl	e->5	
De fr	a->1	å->2	
De få	r->1	
De fö	r->9	
De gj	o->1	
De gr	u->2	ö->6	
De gä	l->1	
De ha	n->1	r->10	
De hå	l->1	
De in	t->1	
De ka	n->6	
De ko	l->1	m->3	
De kr	i->1	ä->1	
De la	n->1	
De lö	s->1	
De mi	n->1	
De my	c->1	
De må	s->5	
De no	r->2	
De nu	v->1	
De ny	a->3	h->1	
De nä	r->1	
De ol	i->3	
De pe	r->1	
De po	l->2	
De pr	o->1	
De re	l->1	
De se	n->4	r->1	
De si	s->2	
De sk	a->4	y->1	
De sl	u->1	
De so	c->1	m->4	
De st	a->4	o->1	r->1	ö->2	
De to	g->1	t->1	
De tu	r->2	
De tv	å->2	
De ty	s->1	
De up	p->2	
De ut	g->1	t->1	
De va	r->2	
De vi	l->1	
De är	 ->4	
De åt	g->2	
Delga	d->1	
Delor	s->3	
Dels 	a->1	
Delvi	s->1	
Demin	i->1	
Demok	r->1	
Den 1	3->1	4->1	
Den 2	3->1	6->1	
Den a	n->18	s->1	v->3	
Den b	e->1	y->1	ö->2	
Den c	e->1	
Den e	n->7	u->8	
Den f	e->1	i->1	j->3	r->3	u->1	å->2	ö->13	
Den g	e->8	r->1	ä->1	
Den h	a->11	o->1	ä->4	ö->1	
Den i	 ->1	n->3	s->1	
Den k	a->5	o->8	r->1	
Den l	i->1	å->1	
Den m	y->1	ä->1	å->7	ö->1	
Den n	e->2	o->1	y->3	ö->1	
Den o	b->2	e->1	m->2	r->2	
Den p	o->2	å->1	
Den r	e->3	i->1	ä->1	ö->2	
Den s	e->1	i->3	j->1	k->4	o->7	t->9	
Den t	a->2	e->1	i->1	r->4	v->2	y->1	
Den u	p->1	t->1	
Den v	a->1	e->2	i->4	ä->1	
Den ä	n->1	r->8	
Den å	t->3	
Den ö	s->1	
Denna	 ->56	
Denne	 ->1	
Deras	 ->2	
Dess 	l->1	s->1	
Dessa	 ->34	
Dessu	t->25	
Det a	l->1	n->10	
Det b	e->23	l->2	r->1	ä->3	ö->6	
Det c	e->1	i->1	
Det d	a->2	e->1	i->1	j->1	å->1	
Det e	g->1	k->1	n->7	u->1	x->1	
Det f	a->10	i->69	r->3	å->7	ö->23	
Det g	e->2	l->5	r->1	y->1	ä->18	å->5	ö->6	
Det h	a->48	i->1	ä->6	ö->1	
Det i	n->12	
Det j	u->1	
Det k	a->16	o->19	r->11	u->2	v->1	
Det l	a->1	i->2	ä->1	ö->1	
Det m	e->1	o->3	å->28	
Det n	u->1	y->1	
Det o	r->1	
Det p	l->1	o->7	r->2	
Det r	i->1	ä->10	å->9	ö->4	
Det s	a->6	e->2	i->2	k->26	l->2	m->1	n->2	o->15	t->16	v->1	y->1	ä->1	å->1	
Det t	i->2	r->1	v->1	y->1	å->1	
Det u	p->1	t->1	
Det v	a->14	e->3	i->21	o->5	ä->1	
Det ä	c->1	n->1	r->359	
Det å	l->1	r->1	t->2	
Det ö	v->3	
Det, 	h->1	
Detal	j->1	
Detsa	m->1	
Detta	 ->208	,->3	
Deuts	c->1	
Dimit	r->5	
Direk	t->9	
Disku	s->1	
Dock 	e->1	g->1	
Dokum	e->1	
Domst	o->3	
Doris	 ->1	
Dubli	n->7	
Duham	e->1	
Duise	n->3	
Dutro	u->1	
Där b	e->1	
Där d	r->1	
Där f	i->2	
Där h	a->4	å->1	
Där j	a->1	
Där k	r->1	
Där l	y->1	
Där m	å->1	
Där v	ä->1	
Där ä	r->1	
Därav	 ->2	
Däref	t->4	
Därem	o->6	
Därfö	r->96	
Däri 	v->1	
Därig	e->2	
Därme	d->4	
Därut	ö->1	
Därvi	d->1	
Då bö	r->1	
Då de	s->1	
Då fi	n->1	
Då fr	a->1	
Då få	r->1	
Då gi	v->1	
Då ha	n->1	r->1	
Då ka	n->3	
Då ko	m->4	
Då må	s->1	
Då oc	h->1	
Då sk	a->1	
Då sy	f->1	
Då ta	l->1	
Då va	r->1	
Då vi	l->1	
Då är	 ->2	
Då öv	e->1	
Díez 	G->1	
Dührk	o->1	
E FRÅ	G->1	
E har	 ->2	
E och	 ->2	
E til	l->1	
E är 	a->1	
E) He	r->1	
E) Ja	g->1	
E) Är	a->1	
E).(E	N->1	
E)Jag	 ->1	
E- oc	h->2	
E-DE)	.->1	
E-DE-	 ->2	g->4	l->1	
E-gru	p->12	
E-kol	i->1	
E-kri	s->3	
E-led	a->1	
E-tes	t->1	
E/NGL	-->2	
EBATT	 ->1	
ECAF:	s->1	
ECHO 	i->1	
ECHO,	 ->1	
ECHO.	D->1	
EDD, 	o->1	
EDD-g	r->2	
EEG t	i->1	
EEG, 	E->2	
EG at	t->1	
EG om	 ->2	
EG sk	u->1	
EG ti	l->2	
EG up	p->1	
EG, E	u->4	
EG, f	ö->1	
EG, o	m->1	
EG, v	i->1	
EG-di	r->2	
EG-do	m->22	
EG-fö	r->8	
EG-in	i->1	
EG-ko	r->16	
EG-rä	t->3	
EG.Vi	 ->1	
EG:s 	d->1	l->1	m->1	
EG?, 	r->1	
EIF h	a->1	
EIF),	 ->1	
EK (d	e->1	
EK(19	9->3	
EK(99	)->1	
EKSG,	 ->2	
EKSG-	f->6	
EL) F	P->1	
EL) H	e->1	
EL) J	a->1	
ELDR 	a->1	
ELDR-	g->1	
ELDR:	s->1	
ELLA 	O->1	
EM-20	0->1	
EMU, 	t->1	
EMU-a	n->1	
EMU-k	r->1	
EMU:s	 ->3	
EN el	l->1	
EN ha	r->1	
EN ko	m->1	
EN oc	h->1	
EN) D	e->2	
EN) F	r->4	å->1	ö->1	
EN) H	e->4	
EN) I	 ->3	
EN) J	a->7	
EN) K	o->1	
EN) L	å->2	
EN) M	i->1	
EN) S	e->1	
EN) T	a->3	i->1	
EN) U	n->1	
EN) V	a->2	
EN) i	n->1	
EN) s	o->1	
EN, a	l->1	
EN, s	o->1	
EN-gr	u->1	
EN:s 	a->2	s->1	v->1	
EO be	f->1	s->1	
EO är	 ->1	
EP ("	d->1	
EP re	p->1	
ERN) 	i->1	
ERREG	,->1	-->1	?->1	
ES) -	 ->1	
ES) ä	r->1	
ES-zo	n->3	
EU "c	o->1	
EU I 	e->1	
EU ag	e->1	
EU at	t->2	
EU bl	a->1	
EU bö	r->1	
EU dä	r->1	
EU fr	a->1	
EU ge	r->1	
EU gö	r->1	
EU ha	r->2	
EU i 	d->1	
EU in	f->2	t->1	
EU ka	n->3	
EU me	r->1	
EU my	c->1	
EU må	s->1	
EU oc	h->4	
EU på	 ->1	
EU re	d->1	
EU sk	a->1	
EU so	m->4	
EU sy	s->1	
EU ut	s->1	v->1	
EU är	 ->2	
EU, f	ö->1	
EU, l	å->1	
EU, m	e->1	
EU, p	å->1	
EU, v	i->1	
EU-bi	s->1	
EU-bu	d->1	
EU-en	h->1	
EU-fo	n->1	
EU-fö	r->5	
EU-ge	n->1	
EU-in	i->1	s->4	
EU-ko	m->2	r->4	
EU-la	g->1	n->1	
EU-lä	n->3	
EU-ma	n->1	
EU-me	d->5	
EU-ni	v->1	
EU-or	d->1	
EU-pr	o->2	
EU-re	g->1	
EU-rä	t->1	
EU-st	r->1	
EU-sä	n->2	
EU-te	x->1	
EU-ut	v->1	
EU-vä	r->1	
EU.. 	(->1	
EU.Al	l->1	
EU.Da	g->1	
EU.De	 ->1	t->1	
EU.Fr	å->1	
EU.Nu	 ->1	
EU.Ro	p->1	
EU.Vi	 ->3	
EU:s 	B->1	b->6	e->1	f->3	g->1	h->1	i->6	k->2	l->2	m->4	n->1	o->5	p->3	r->1	s->4	t->2	u->1	
EU?He	r->1	
EUGFJ	)->2	:->1	
Ecemi	s->1	
Edinb	u->1	
Effek	t->5	
Eftar	l->2	
Efter	 ->20	s->28	
Egypt	e->2	
Ehud 	B->2	
Eieck	 ->1	
Ekofi	n->2	
Ekono	m->3	
Elisa	b->1	
Eller	 ->1	
Elles	 ->3	
Elmar	 ->2	
Elst.	D->1	
Emell	e->8	
Emili	a->1	
En al	l->3	
En an	d->1	n->5	
En as	p->1	
En av	 ->6	
En be	l->1	
En bo	e->1	m->1	
En bä	t->1	
En de	l->7	
En fr	i->1	å->1	
En fö	r->2	
En ge	n->1	
En ka	t->1	
En kn	a->1	
En ko	m->1	n->2	
En ma	j->1	
En me	d->1	
En pe	r->1	
En pr	o->1	
En ra	d->2	
En re	s->1	v->1	
En sa	k->1	
En si	s->1	
En su	c->1	
En sy	s->1	
En sä	r->1	
En så	 ->1	d->3	
En up	p->1	
En va	r->1	
En ve	r->1	
En vi	k->3	t->1	
En vä	l->1	s->2	x->1	
En ök	a->1	
En öv	e->1	
Enbar	t->1	
Endas	t->11	
Enkel	t->1	
Enlig	t->37	
Equal	 ->6	"->1	,->1	
Equqa	l->2	
Er an	s->1	
Era t	v->1	
Erfar	e->2	
Erika	 ->14	,->5	-->1	.->2	s->7	
Eritr	e->1	
Erkki	 ->2	
Ert b	e->1	
Ert p	a->1	
Etiop	i->3	
Ett E	u->1	
Ett a	n->6	s->1	v->4	
Ett d	i->2	
Ett e	f->1	x->4	
Ett f	e->2	l->1	ö->1	
Ett h	ö->1	
Ett l	ä->1	
Ett m	y->1	
Ett n	y->3	
Ett o	m->2	
Ett p	å->1	
Ett s	a->1	e->1	i->2	o->1	t->1	y->2	å->2	
Ett t	r->1	y->1	
Ett v	e->1	i->2	
Ett å	r->1	
Eurat	o->4	
Euro-	r->1	
Eurod	a->5	
Euroj	u->6	
Euron	s->1	
Europ	a->459	e->357	o->16	
Euros	k->1	t->1	
Evans	 ->3	,->4	
Event	u->1	
Excep	t->1	
Exemp	e->1	
Exper	t->2	
Exupé	r->1	
Exxon	 ->3	
F gör	a->1	
F har	 ->1	
F i e	t->1	
F i r	ä->1	
F kan	 ->1	
F kon	t->1	
F ska	p->1	
F) är	 ->1	
F), b	i->1	
F, Eu	r->1	
F, de	n->1	
F, en	 ->1	
F, ko	m->1	
F, så	 ->2	
F, vi	l->1	
F, öv	e->1	
F.All	t->1	
F.För	 ->1	
F.Her	r->1	
F.Men	 ->1	
F:s (	f->1	
F:s u	t->1	
FAF, 	s->1	
FBI -	 ->1	
FEO b	e->2	
FEO ä	r->1	
FI) J	a->1	
FIL, 	f->1	
FIPOL	)->1	
FJ) f	i->1	
FJ), 	ä->1	
FJ:s 	g->1	
FMI d	ä->1	
FN, s	o->1	
FN-up	p->1	
FN.He	r->1	
FN:s 	a->1	b->2	e->1	g->1	r->1	s->2	
FOP).	V->1	
FPÖ (	Ö->2	
FPÖ f	ö->1	
FPÖ h	ä->1	
FPÖ i	n->1	
FPÖ m	i->1	
FPÖ o	c->2	m->1	
FPÖ s	o->1	
FPÖ v	i->1	
FPÖ ä	r->1	
FPÖ).	J->1	
FPÖ-l	e->1	
FPÖ-m	e->1	
FPÖ:s	 ->4	
FR) "	T->1	
FR) D	e->4	
FR) E	f->1	
FR) F	r->1	
FR) H	e->1	
FR) I	 ->2	
FR) J	a->3	ö->1	
FR) N	e->1	ä->2	
FR) T	h->1	
FRÅGO	R->1	
FSR -	 ->1	
FUF) 	ä->1	
Fackf	ö->3	
Facto	r->1	
Faktu	m->4	
Farli	g->1	
Farou	k->1	
Fasci	s->1	
Feira	,->2	
Felak	t->1	
Fem l	ä->1	
Fina 	f->1	o->1	s->1	
Fina.	H->1	
Finan	s->2	
Finla	n->6	
Finns	 ->4	
Firma	n->1	
Fisch	l->4	
Flaut	r->2	
Flera	 ->3	
Flert	a->1	
Flore	n->19	
Fléch	a->1	
FoU, 	n->1	
FoU-r	a->1	
Fog f	ö->1	
Folk 	r->1	s->1	t->1	
Folkf	r->1	
Folkr	e->2	
Fonta	i->1	
Ford,	 ->1	
Fores	t->1	
Forsk	a->1	n->1	
Fraga	.->1	
Fram 	t->1	
Framf	ö->2	
Framl	ä->1	
Frams	t->2	
Framt	a->1	i->1	
Framå	t->1	
Franc	e->2	i->1	
Frank	r->39	
Frano	i->1	
Frans	m->2	
Franz	 ->3	
Franç	o->1	
Frass	o->1	
Freds	p->1	
Frihe	t->3	
Fru A	h->1	
Fru B	e->1	
Fru L	y->1	
Fru M	c->1	
Fru P	l->1	
Fru S	c->1	
Fru k	o->4	
Fru l	e->2	
Fru t	a->70	
Frute	a->3	
Främj	a->1	
Främs	t->1	
Fråga	 ->21	n->16	
Fråge	s->2	
Frågo	r->3	
Från 	k->1	o->1	
Fund 	L->1	
Fyrti	o->1	
Fästn	i->1	
Får j	a->3	
Följa	k->5	
Följd	e->1	
För 1	9->2	
För a	t->31	
För b	a->1	
För d	e->100	
För e	g->1	n->3	
För f	ö->2	
För i	 ->1	
För k	o->1	
För l	e->1	
För m	a->1	e->1	i->6	å->1	
För n	ä->7	å->1	
För o	m->2	s->4	
För p	e->1	
För s	t->2	ä->1	
För t	i->2	v->2	
För u	n->1	
För v	a->1	i->4	å->2	
För å	t->1	
För ö	g->1	r->1	v->1	
Förbu	d->2	n->3	
Förde	l->1	
Fördr	a->2	
Föreb	y->1	
Föred	r->8	
Fören	a->15	l->1	t->28	
Föret	a->1	r->1	
Förfa	r->1	
Förhi	n->1	
Förho	p->3	
Förin	t->2	
Förlu	s->1	
Förmo	d->1	
Föror	e->1	
Förpa	c->1	
Försi	k->1	
Försl	a->8	
Först	 ->25	a->2	å->1	
Försä	m->1	
Försö	k->1	
Förtj	ä->1	
Förtr	o->1	
Förut	o->6	s->1	
Förva	l->1	
Förvi	s->2	
Förvä	n->1	
Förän	d->1	
G att	 ->1	
G om 	t->1	u->1	
G sku	l->1	
G til	l->2	
G upp	f->1	
G(Par	l->1	
G, EE	G->2	
G, Eu	r->4	
G, fö	r->1	
G, om	 ->1	
G, vi	l->1	
G-dir	e->2	
G-dom	s->22	
G-för	d->14	
G-ini	t->1	
G-kor	t->16	
G-rät	t->3	
G.(EN	)->1	
G.Vi 	v->1	
G:s d	i->1	
G:s l	a->1	
G:s m	i->1	
G?, r	å->1	
GA-st	ö->1	
GASP 	m->1	
GFJ) 	f->1	
GFJ),	 ->1	
GFJ:s	 ->1	
GL-gr	u->2	
GORNä	s->1	
GUE/N	G->2	
GUSP 	o->1	
Galeo	t->1	
Galic	i->2	
Gama 	-->1	p->1	u->1	
Garga	n->5	
Gaza 	o->1	
Gaza,	 ->1	
Gaza.	D->1	S->1	
Gazar	e->2	
Gemel	l->1	
Gemen	s->5	
Gener	a->9	e->1	
Genom	 ->24	f->3	s->1	
Genèv	e->3	
Ger d	e->1	
Gil-D	e->1	
Gil-R	o->1	
Gino,	 ->1	
Givet	v->2	
Goebb	e->1	
Golan	 ->3	.->1	?->1	h->4	
Golfs	t->3	
Golln	i->1	
Gomes	,->1	
Gonzá	l->1	
Goodw	i->1	
Gorse	l->1	
Gott 	n->1	
Graca	 ->3	
Graco	-->1	
Gratu	l->1	
Graça	 ->5	
Grekl	a->14	
Gross	e->2	t->1	
Grund	e->1	
Grupp	e->10	
Gröna	/->1	
Gröni	t->1	
Guate	m->1	
Guigo	u->1	
Gulfk	r->1	
Gusp"	,->1	
Guter	r->2	
Gälla	n->1	
Gå he	m->1	
Gör v	i->2	
Göteb	o->1	
H BRÅ	D->1	
H-000	6->1	
H-077	8->1	
H-078	0->1	1->1	2->1	5->1	6->1	8->1	
H-079	1->1	3->1	5->1	6->1	8->1	
H-080	1->1	5->1	7->1	8->1	
H-081	3->1	7->1	9->1	
H-082	9->1	
HO i 	b->1	
HO, a	k->1	
HO.De	t->1	
Haard	e->1	
Hade 	d->1	v->1	
Hader	a->1	
Hague	,->1	
Haide	r->37	
Hambu	r->1	
Han a	v->1	
Han b	e->1	
Han h	a->6	ä->1	
Han k	a->1	
Han n	ä->1	
Han s	a->3	
Han t	a->1	
Han ä	r->3	
Hande	l->1	
Handi	k->1	
Handl	i->2	
Hans 	H->1	f->1	h->1	
Har k	o->3	
Har m	a->2	
Har o	r->1	
Har r	e->1	å->1	
Har v	i->3	
Harri	s->1	
Hatzi	d->2	
Haven	,->1	
Heato	n->1	
Hebro	n->1	
Hedge	 ->1	
Hedkv	i->1	
Heinz	 ->2	
Hela 	f->1	p->1	s->1	
Helig	h->1	
Helsi	n->20	
Helt 	k->1	n->1	
Hemli	g->1	
Henry	 ->1	
Herr 	A->1	B->2	G->1	P->2	S->1	W->1	f->1	k->12	l->5	m->1	o->3	p->2	r->5	t->292	
Hicks	.->1	
Hilto	n->1	
Himal	a->1	
Histo	r->2	
Hit h	ö->3	
Hitle	r->6	
Hitti	l->3	
Holly	w->1	
Holzm	a->2	
Hon h	a->2	
Hon l	i->1	
Hon s	ä->1	
Hoppe	t->1	
Howit	t->1	
Huhne	,->1	
Hulte	n->19	
Hulth	e->6	
Hur b	e->1	
Hur f	ö->2	
Hur g	ö->1	
Hur h	a->1	
Hur k	a->1	o->2	
Hur l	i->1	ä->1	
Hur m	y->1	å->3	
Hur s	e->3	k->6	o->8	t->1	v->1	
Hur t	ä->1	
Hur ä	r->1	
Huruv	i->1	
Huvud	a->2	d->1	f->1	l->1	m->2	
Hyckl	e->1	
Hände	l->2	
Hänsc	h->2	
Här b	e->3	ä->1	ö->1	
Här f	i->1	ö->2	
Här g	e->1	
Här h	a->4	
Här i	n->1	
Här k	a->3	o->2	
Här m	å->2	
Här n	ö->1	
Här r	i->1	ä->1	
Här s	k->1	
Här t	a->1	i->1	r->1	
Här v	i->3	
Här ä	g->1	r->1	
Härme	d->2	
Härom	 ->1	
Hålle	r->1	
Höger	e->1	
I - K	o->1	
I - P	a->1	
I - R	å->1	
I - d	e->1	
I Ams	t->1	
I Eur	o->4	
I Fra	n->2	
I Hel	s->1	
I Irl	a->2	
I Ita	l->1	
I Ned	e->1	
I Rap	k->1	
I Sch	r->1	
I Tib	e->1	
I Tur	k->1	
I Tys	k->1	
I all	a->3	
I and	r->1	
I ann	a->2	
I apr	i->1	
I art	i->1	
I avs	a->1	
I avv	a->2	
I bet	r->1	ä->5	
I bud	g->1	
I bör	j->2	
I dag	 ->22	s->2	
I de 	k->1	n->1	
I den	 ->18	n->5	
I det	 ->22	t->13	
I dir	e->1	
I där	 ->1	
I ege	n->7	
I en 	b->1	c->1	r->1	s->1	t->3	
I enl	i->4	
I era	 ->1	
I ett	 ->2	
I fjo	l->1	
I fle	r->1	
I for	t->1	
I fra	m->1	
I frå	g->5	
I för	h->1	p->1	r->1	s->3	
I går	 ->2	d->1	
I har	 ->2	
I i E	U->1	
I i a	n->1	
I i f	ö->1	
I jun	i->1	
I kla	r->1	
I kom	m->2	
I kon	s->1	
I kri	t->1	
I lik	h->7	
I med	d->1	
I min	a->1	
I mit	t->1	
I mor	g->2	s->1	
I mot	s->3	
I mål	 ->1	
I nov	e->2	
I näs	t->2	
I och	 ->8	
I okt	o->1	
I par	l->1	
I per	 ->2	
I pri	n->1	
I pro	g->1	
I rap	p->2	
I rea	l->1	
I reg	i->1	
I res	o->5	
I rev	i->1	
I rät	t->1	
I råd	e->1	
I sam	b->3	
I sin	 ->1	
I sit	t->2	
I sjä	l->4	
I ska	l->1	
I slu	t->3	
I sti	l->1	
I str	u->1	
I stä	l->9	
I syn	n->1	
I sys	t->1	
I så 	f->1	m->2	
I såd	a->1	
I tju	g->1	
I upp	f->1	
I utb	y->1	
I uts	k->1	
I var	j->2	
I ver	k->1	
I vil	k->3	
I vis	s->2	
I vit	b->2	
I von	 ->1	
I vän	t->2	
I vår	 ->1	a->3	t->2	
I änd	r->1	
I övr	i->3	
I) Ja	g->1	
I) oc	h->1	
I); e	n->1	
I, et	t->1	
I, ha	n->1	
I-pro	g->3	
I. fö	r->2	
I:e r	a->2	
ICES)	 ->1	
ICES-	z->3	
IF ha	r->1	
IF), 	b->1	
IFIL,	 ->1	
IFOP)	.->1	
II - 	K->1	R->1	
II ha	r->2	
II i 	f->1	
II kr	i->1	
II sk	a->1	
II) o	c->1	
II, h	a->1	
II-pr	o->2	
II. f	ö->1	
II:e 	r->2	
III -	 ->1	
III h	a->1	
III k	r->1	
III s	k->1	
III:e	 ->1	
IK, v	i->1	
IK.De	t->2	
IL, f	i->1	
IMO).	F->1	
IMO.D	e->1	
IMO:s	 ->1	
INA h	a->1	
INA v	a->1	
INA, 	e->1	
ING(P	a->1	
ING.(	E->1	
INTE 	h->1	
INTER	R->3	
IPOL)	,->1	
IRA h	a->1	
ISPA-	i->1	
IT) D	e->1	
IT) H	e->1	
IT) O	m->1	
IV - 	D->1	
IV i 	E->1	f->1	
IX oc	h->1	
IX, f	a->1	
Iblan	d->3	
Idén 	o->1	
Ihåll	a->1	
Ile-d	e->1	
Illeg	a->1	
Imben	i->3	
Immig	r->1	
Indie	n->5	
Indus	t->1	
Inför	 ->4	
Inga 	g->1	m->1	
Ingen	 ->8	,->1	t->1	
Inger	 ->1	
Inget	 ->2	d->1	
Ingle	w->2	
Initi	a->3	
Inneb	ö->1	
Inneh	å->1	
Inom 	E->1	d->3	e->1	j->1	r->3	u->1	
Inre 	m->1	
Inres	a->1	
Inrät	t->1	
Insat	s->2	
Inte 	b->1	e->3	f->2	h->3	m->2	p->1	s->1	u->1	ä->1	
Inter	n->21	
Irlan	d->22	
Isabe	l->2	
Islan	d->1	
Israe	l->38	
Istan	b->1	
Itali	e->18	
Izqui	e->1	
J) fi	n->1	
J), ä	r->1	
J:s g	a->1	
Ja Er	i->1	
Ja el	l->1	
Ja ti	l->1	
Ja, d	e->1	
Ja, f	r->1	
Ja, h	e->2	
Ja, j	a->1	
Ja, n	a->1	
Ja, s	o->1	
Ja, v	i->1	
Jacks	o->2	
Jacob	 ->2	
Jacqu	e->3	
Jag a	c->1	n->61	v->2	
Jag b	a->1	e->26	l->6	o->1	
Jag d	e->6	r->2	
Jag e	r->1	
Jag f	i->1	r->7	å->2	ö->38	
Jag g	e->2	l->7	o->1	r->3	
Jag h	a->47	o->38	ä->3	å->9	ö->1	
Jag i	n->9	
Jag j	ä->1	
Jag k	a->33	o->11	ä->6	
Jag l	a->1	y->1	ä->1	
Jag m	e->5	i->4	o->3	ä->1	å->13	
Jag n	o->2	ä->2	
Jag o	m->1	
Jag p	e->1	l->1	r->1	å->2	
Jag r	e->4	ä->5	ö->5	
Jag s	a->2	e->4	k->109	o->1	t->9	y->2	ä->3	å->1	
Jag t	a->19	i->3	r->72	v->1	y->27	ä->11	
Jag u	n->5	p->20	t->6	
Jag v	a->2	e->18	i->173	ä->18	å->1	
Jag ä	r->56	
Jag ö	n->5	v->6	
Jan-K	e->1	
Japan	 ->2	,->1	
Javet	t->1	
Jean-	C->1	
Jerus	a->2	
Jo då	,->1	
Jo, d	e->1	
Jo, i	 ->1	
Jo, s	y->1	
Jonas	 ->2	
Jonck	h->14	
Jorda	n->2	
Jordb	r->2	
Jospi	n->1	
Ju mi	n->1	
Jugos	l->1	
Junke	r->1	
Just 	a->1	d->1	h->1	i->2	n->2	p->1	
Juste	r->2	
Jämfö	r->2	
Jämst	ä->1	
Jörg 	H->14	
Jørge	n->2	
K (de	t->1	
K nu 	ä->1	
K(199	8->3	
K(99)	0->1	
K, de	t->1	
K, vi	 ->1	
K.Det	 ->2	
KANDE	 ->1	
KOM(1	9->8	
KOM(9	8->1	9->1	
KSG, 	E->2	
KSG-f	ö->6	
KTUEL	L->1	
Kafor	 ->1	
Kalei	d->2	
Kalej	d->1	
Kan k	o->5	
Kan m	a->1	
Kan n	i->4	
Kan r	å->1	
Kan u	n->1	
Kan v	i->1	
Kanad	a->1	
Kansk	e->9	
Kanta	b->3	
Karas	 ->3	
Karl 	H->1	v->3	
Karl-	H->1	
Karls	r->2	
Karte	l->2	
Kaspi	s->1	
Katas	t->1	
Kaufm	a->1	
Kauka	s->3	
Kazak	s->1	
Kees 	W->1	
Kfor 	s->1	
Kina 	a->2	e->1	f->1	g->1	i->1	o->1	
Kina,	 ->1	
Kina.	U->1	
Kinas	 ->1	
Kinno	c->24	
Kirgi	z->5	
Knapp	t->1	
Koch 	f->3	h->1	t->2	
Koch)	D->1	
Koch,	 ->5	
Koch.	J->1	
KochI	 ->1	
Kochs	 ->1	
Koden	 ->1	
Kolle	g->1	
Kom i	h->1	
Komme	r->12	
Kommi	s->106	t->1	
Kommu	n->1	
Kompr	o->1	
Konkr	e->1	
Konku	r->13	
Konra	d->1	
Konse	k->1	
Konst	i->1	
Konsu	m->3	
Konve	n->2	
Korea	 ->2	
Kort 	s->2	
Kosov	o->60	
Kostn	a->4	
Kouch	n->12	
Krav 	p->1	
Krave	n->1	t->1	
Kultu	r->25	
Kumar	 ->1	
Kungl	i->1	
Kvant	i->1	
Kvinn	o->5	
Kväka	r->1	
Kyoto	 ->2	-->1	.->1	p->2	s->1	
Känne	r->1	
Kära 	k->6	
Kärna	n->1	
Kärnk	r->2	
Kärnt	e->1	
Köln 	a->1	i->1	
Köpen	h->1	
L (en	 ->1	
L) At	t->1	
L) FP	Ö->1	
L) He	r->4	
L) Ja	g->1	
L), m	e->1	
L, fi	n->1	
L-gru	p->2	
LA OC	H->1	
LAF g	ö->1	
LAF i	 ->2	
LAF k	a->1	o->1	
LAF s	k->1	
LAF, 	E->1	d->1	e->1	k->1	s->1	v->1	ö->1	
LAF.A	l->1	
LAF.F	ö->1	
LAF.H	e->1	
LAF.M	e->1	
LAF:s	 ->1	
LAS (	I->1	
LDR a	n->1	
LDR-g	r->1	
LDR:s	 ->1	
LFAF,	 ->1	
LLA O	C->1	
LTCM.	A->1	
La Ré	u->2	
Laan 	f->1	
Laan.	V->1	
Laans	 ->5	
Lama 	h->1	o->1	s->1	
Lama.	J->1	V->1	
Lamas	 ->2	
Landi	s->1	
Lands	b->1	
Lange	 ->11	,->1	n->17	s->1	
Lanka	 ->2	.->1	
Lappl	a->2	
Le Be	s->1	
Leade	r->5	
Ledam	o->3	ö->1	
Ledni	n->1	
Leine	n->6	
Leins	t->2	
Leoni	 ->1	
Liban	o->5	
Liber	a->2	
Libye	n->1	
Liika	n->3	
Lika 	v->1	
Likas	å->2	
Likri	k->1	
Likso	m->8	
Likvä	l->1	
Lille	 ->1	
Lissa	b->8	
Litau	e->1	
Litte	r->1	
Livli	g->2	
Livsm	e->3	
Lloyd	s->1	
Loire	 ->1	,->1	-->1	
Loméa	v->1	
Lomék	o->1	
Londo	n->4	
Lord 	I->2	
Lorra	i->2	
Lotha	r->3	
Louse	w->1	
Loyol	a->2	
Lutte	 ->1	
Luxem	b->6	
Lycka	s->1	
Lyckl	i->1	
Lynne	 ->1	!->1	s->2	
Lägg 	d->1	m->1	
Lände	r->1	
Lån a	v->1	
Långr	a->1	
Låt e	r->1	
Låt i	n->1	
Låt m	i->40	
Låt o	s->18	
Låt v	å->1	
Lööw 	f->1	
M AKT	U->1	
M som	 ->1	
M(199	7->1	9->7	
M(98)	0->1	
M(99)	0->1	
M-200	0->1	
M.Att	 ->1	
MARPO	L->1	
MI dä	r->1	
MIK, 	v->1	
MIK.D	e->2	
MO).F	ö->1	
MO.De	t->1	
MO:s 	n->1	
MRÖST	N->2	
MU, t	y->1	
MU-an	p->1	
MU-kr	i->1	
MU:s 	d->1	h->1	o->1	
Maast	r->6	
Macao	 ->1	
Madag	a->1	
Madei	r->2	
Madri	d->3	
Mains	t->1	
Major	i->1	
Malta	 ->5	,->1	s->1	
Man b	e->1	ö->7	
Man f	o->1	r->1	å->1	
Man g	å->1	ö->1	
Man h	a->4	
Man i	n->1	
Man j	a->1	
Man k	a->10	o->2	
Man l	ä->1	
Man m	å->14	
Man r	ö->1	
Man s	a->1	k->2	
Man t	e->1	i->1	
Man u	p->3	
Man v	i->1	
Manne	n->1	s->1	
Marga	r->1	
Margo	t->1	
Maria	 ->1	
Marie	 ->1	
Marin	h->6	
Markn	a->4	
Marko	v->1	
Marpo	l->1	
Marse	i->1	
Marti	n->1	
Mathi	e->2	
Maxim	a->1	i->1	
McCar	t->1	
McNal	l->5	
Med a	n->2	v->1	
Med d	e->12	
Med e	n->2	
Med f	ö->1	
Med h	j->1	ä->5	
Med o	m->2	
Med s	a->1	t->1	
Med t	a->6	i->1	
Medan	 ->3	,->1	
Medbe	s->1	
Medbo	r->2	
Medel	h->3	
Medge	r->1	
Medle	m->9	
Mella	n->20	
Men -	 ->2	
Men C	E->1	
Men E	u->1	
Men F	E->1	
Men a	l->1	n->1	t->2	v->1	
Men b	o->1	å->1	
Men d	e->52	i->1	ä->2	
Men e	f->2	n->3	r->1	
Men f	o->1	r->1	ö->5	
Men g	e->1	
Men h	a->3	o->1	u->3	
Men i	 ->4	d->1	n->4	
Men j	a->31	u->2	
Men k	a->2	o->2	v->1	
Men m	a->1	e->3	
Men n	u->2	ä->2	å->1	
Men o	a->1	m->3	
Men p	e->1	l->1	o->2	å->1	
Men s	a->5	e->1	o->3	t->1	ä->1	å->2	
Men t	r->1	y->2	
Men u	n->1	p->1	r->2	
Men v	a->1	e->2	i->29	
Men ä	v->3	
Men å	 ->1	
Men, 	f->2	h->1	
Menar	 ->1	
Menta	l->1	
Mer s	p->1	
Mer v	o->1	
Mer ä	n->1	
Mexik	o->1	
Michi	e->1	
Midde	l->1	
Midla	n->1	
Miljö	m->1	
Min a	n->3	v->3	
Min d	e->1	
Min f	r->4	ö->1	
Min g	r->9	
Min k	o->1	
Min p	e->1	
Min s	i->3	p->1	
Min t	r->2	
Min u	p->1	
Min å	s->1	
Min ö	n->1	
Mina 	d->11	f->1	k->3	s->1	u->1	ä->1	
Mindr	e->1	
Minis	t->1	
Minns	 ->1	
Minsk	a->1	
Minuc	 ->1	
Miste	r->2	
Mitro	v->1	
Mitt 	l->1	p->2	
Mitte	r->2	
Monti	 ->10	!->3	,->2	.->2	
Montr	e->2	
Moral	,->1	
Morat	i->4	
Morbi	h->1	
Morga	n->4	
Moskv	a->1	
Mot b	a->4	
Mot d	e->4	
Moura	 ->6	,->2	
Mousk	o->1	
Mulde	r->1	
Mycke	t->1	
Mylle	r->1	
Myndi	g->3	
Männi	s->5	
Märkl	i->1	
Måhän	d->1	
Målet	 ->2	
Många	 ->10	
Möjli	g->2	
Münch	e->1	
N ell	e->1	
N har	 ->1	
N kom	m->1	
N och	 ->1	
N) De	n->2	
N) Fr	u->4	
N) Få	r->1	
N) Fö	r->1	
N) He	r->4	
N) I 	S->1	d->1	g->1	
N) Ja	,->1	g->6	
N) Ko	m->1	
N) Lå	t->2	
N) Mi	t->1	
N) Se	d->1	
N) Ta	c->3	
N) Ti	d->1	
N) Un	d->1	
N) Va	d->2	
N) i 	G->1	
N) in	t->1	
N) so	m->1	
N)). 	V->1	
N, al	l->1	
N, so	m->2	
N-gru	p->1	
N-upp	d->1	
N.Her	r->1	
N:s a	n->1	r->2	
N:s b	e->2	
N:s e	k->1	
N:s g	i->1	
N:s r	e->1	
N:s s	a->1	i->1	ä->1	
N:s v	e->1	
NA ha	r->1	
NA va	r->1	
NA, e	f->1	
NDE F	R->1	
NG(Pa	r->1	
NG.(E	N->1	
NGL-g	r->2	
NI be	t->1	
NI i 	a->1	
NI oc	h->2	
NI pe	r->2	
NI, e	t->1	
NIFIL	,->1	
NING(	P->1	
NING.	(->1	
NL) A	t->1	
NL) H	e->3	
NMIK,	 ->1	
NMIK.	D->2	
NP jä	m->1	
NP mi	n->1	
NP pe	r->3	
NP på	 ->1	
NP år	 ->1	
NP, i	 ->1	
NP, m	e->1	
NS)) 	(->1	
NS))(	G->1	P->3	
NS)).	.->1	J->1	
NS))F	r->1	
NS))o	c->1	
NTE h	a->1	
NTERR	E->3	
Nally	 ->1	!->1	.->1	b->1	s->1	
Nana 	M->1	
Napol	i->1	
Narko	t->1	
Natio	n->7	
Nato 	i->1	
Natoa	k->1	
Natob	a->1	
Natos	 ->2	
Natur	l->15	
Neder	l->9	
Nej, 	b->1	d->1	h->1	j->1	m->1	n->1	s->1	
Nej.I	 ->1	
New Y	o->1	
Ni ag	e->1	
Ni be	g->1	s->1	t->1	
Ni bo	r->1	
Ni fr	a->1	
Ni fö	r->2	
Ni ha	r->11	
Ni ka	n->2	
Ni ko	m->5	
Ni kä	n->2	
Ni lä	t->1	
Ni må	s->4	
Ni nä	m->1	
Ni sa	d->3	
Ni sk	a->2	
Ni sä	g->1	
Ni ta	l->2	
Ni ve	t->2	
Ni vi	l->1	
Niels	e->1	o->5	
Nikit	i->2	
Nivån	 ->1	
Nogue	i->1	
Noirm	o->1	
Nordi	s->2	t->1	
Norge	 ->1	,->1	
Norma	n->1	
Norme	r->1	
Nu an	g->1	m->1	
Nu be	h->1	
Nu fi	n->1	
Nu få	r->1	
Nu fö	r->1	
Nu ha	r->6	
Nu ho	t->1	
Nu ka	n->2	
Nu må	s->1	
Nu ti	l->1	
Nu ve	r->1	
Nu vä	n->1	
Nu är	 ->7	
Nu åt	e->1	
Numer	a->1	
Nuvar	a->1	
Nya Z	e->2	
Nya r	e->1	
Nylig	e->1	
Nytt 	I->1	
När a	l->3	
När b	a->1	l->1	
När d	e->35	
När e	t->1	
När f	e->1	
När j	a->7	
När k	o->6	
När m	a->6	e->1	
När n	ä->1	
När p	l->1	
När s	e->1	
När t	i->1	ä->1	
När v	i->15	ä->1	
Nästa	 ->26	
Någon	s->1	t->1	
Något	 ->1	
Några	 ->2	
Nåja,	 ->1	
Nödvä	n->1	
O bef	i->1	
O bes	t->1	
O i b	u->1	
O är 	p->1	
O).Fö	r->1	
O, ak	t->1	
O.Det	 ->2	
O:s n	u->1	
O?End	a->1	
OCH B	R->1	
OD)) 	(->2	i->2	
OD))(	P->4	
OD)).	.->2	F->1	
OD))H	e->1	
OD)].	)->1	
OFSR 	-->1	
OK, d	e->1	
OL (e	n->1	
OL), 	m->1	
OLAF 	g->1	i->2	k->2	
OLAF,	 ->7	
OLAF.	A->1	F->1	H->1	M->1	
OLAF:	s->1	
OLAS 	(->1	
OLFAF	,->1	
OM AK	T->1	
OM(19	9->8	
OM(98	)->1	
OM(99	)->1	
OMRÖS	T->2	
OP).V	i->1	
ORNäs	t->1	
OS)].	H->2	
OSSE 	t->1	
Oavse	t->2	
Oberb	a->1	
Obero	e->2	
Och E	u->1	
Och S	i->1	
Och a	b->1	p->1	
Och d	a->1	e->18	r->1	å->1	
Och e	f->1	r->1	
Och g	i->1	
Och h	ä->1	
Och i	 ->1	n->1	
Och j	a->10	
Och k	o->1	
Och m	e->1	
Och n	i->1	u->2	ä->2	
Och o	m->2	
Och s	k->1	l->3	o->2	å->1	
Och t	i->1	
Och v	a->3	e->1	i->3	å->1	
Och ä	v->1	
Och: 	V->1	
Också	 ->2	
Offen	t->3	
Offic	e->1	
Ofta 	h->1	
Oil P	o->1	
Oil-p	r->1	
Olika	 ->1	
Olivi	e->1	
Oljeb	ä->2	
Oljet	a->1	
Olymp	i->1	
Om 50	 ->1	
Om EU	:->1	
Om Eu	r->1	
Om Sc	h->1	
Om Sy	r->1	
Om al	l->3	
Om be	f->1	
Om de	 ->2	n->2	r->1	s->3	t->13	
Om do	m->1	
Om du	 ->1	
Om en	 ->2	
Om er	t->1	
Om et	t->2	
Om fo	r->1	
Om ge	m->1	
Om gi	l->1	
Om in	n->1	t->3	
Om ja	g->2	
Om ka	m->1	
Om ko	a->1	m->2	n->1	
Om la	g->1	
Om ma	n->11	
Om ni	 ->7	
Om nå	g->1	
Om om	r->1	
Om pa	r->2	
Om re	f->1	
Om rå	d->1	
Om sl	u->1	
Om sy	s->1	
Om tr	e->1	
Om tv	å->1	
Om up	p->1	
Om vi	 ->23	
Omagh	 ->1	
Omrös	t->15	
Onest	a->1	
Onödi	g->1	
Orani	n->1	
Ord s	o->1	
Orden	 ->1	
Order	i->1	
Ordet	 ->1	
Ordfö	r->7	
Orkan	e->2	
Oron 	a->1	
Orovä	c->1	
Orsak	e->2	
Oslo 	o->1	
Oslo,	 ->2	
Osman	.->1	
Ouvri	è->1	
Oz dy	k->1	
Oz ha	d->1	
Oz, b	e->1	
P ("d	i->1	
P (Ös	t->2	
P att	 ->2	
P jäm	f->1	
P min	s->1	
P mis	s->1	
P mås	t->1	
P och	 ->1	
P per	 ->3	
P på 	m->1	
P rep	r->1	
P år 	1->1	
P) oc	h->1	
P).Vi	d->1	
P, ef	t->1	
P, i 	v->1	
P, me	d->1	
PA-in	s->1	
PE ha	r->1	
PE är	 ->1	
PE-DE	)->1	-->7	
PE-gr	u->5	
PM so	m->1	
POL (	e->1	
POL),	 ->1	
PPE h	a->1	
PPE ä	r->1	
PPE-D	E->8	
PPE-g	r->5	
PR-ef	f->1	
PSE)J	a->1	
PSE-g	r->3	
PT) E	f->1	
PT) F	r->1	
PT) H	e->9	
PT) J	a->2	
PT) L	e->1	
PT) N	ä->1	
PT) V	i->1	
PVC, 	a->1	
PVC-l	e->1	
PVC.V	i->1	
Pack 	a->1	h->1	
Packs	 ->1	
Paddi	n->2	
Pakis	t->5	
Palac	i->15	
Paler	m->1	
Pales	t->10	
Papay	a->2	
Parag	r->1	
Paris	 ->1	,->1	f->1	
Parla	m->42	
Patte	n->23	
Pays 	d->1	
Pays-	d->1	
Peake	,->1	
Peijs	 ->1	.->1	
Pekin	g->1	
Perso	n->4	
Peter	s->1	
Petro	l->1	
Plane	r->1	
Plant	a->1	
Plast	-->1	i->1	
Plath	 ->3	,->1	
Plato	n->1	
Plooi	j->1	
Pläde	r->1	
Poett	e->5	
Pohja	m->1	
Polen	 ->1	
Pollu	t->1	
Pomés	 ->1	
Ponna	m->1	
Poos 	a->1	
Portu	g->27	
Power	 ->1	,->2	
Preci	s->6	
Prese	n->1	
Preus	s->1	
Prior	i->1	
Probl	e->9	
Proce	n->1	s->2	
Prodi	 ->17	,->1	.->2	;->1	s->7	
Produ	c->2	
Progr	a->1	
Proje	k->2	
Proto	k->2	
Prova	n->3	
Prínc	i->1	
Punkt	 ->2	
Purvi	s->1	
PÖ (Ö	s->2	
PÖ fö	r->1	
PÖ hä	v->1	
PÖ in	o->1	
PÖ mi	n->1	
PÖ oc	h->3	
PÖ om	 ->1	
PÖ so	m->1	
PÖ vi	d->1	
PÖ är	 ->1	
PÖ) s	i->1	
PÖ).J	a->1	
PÖ-le	d->1	
PÖ-me	d->1	
PÖ:s 	a->1	d->1	f->1	s->1	
På al	l->1	
På de	n->12	t->10	
På et	t->1	
På gr	u->2	
På la	n->1	
På ma	r->1	
På mi	l->1	
På må	n->1	
På om	r->2	
På pa	p->1	
På sa	m->4	
På si	n->3	
På så	 ->4	
På up	p->1	
På vi	l->3	
Påstå	e->1	
Pétai	n->1	
Quece	d->1	
R - o	m->1	
R ans	e->1	
R) "T	y->1	
R) De	n->2	t->2	
R) Ef	t->1	
R) Fr	u->1	
R) He	r->1	
R) I 	d->1	s->1	
R) Ja	g->3	
R) Jö	r->1	
R) Ne	j->1	
R) Nä	r->2	
R) Th	y->1	
R) oc	h->1	
R-eff	e->1	
R-gru	p->1	
R.Sed	a->1	
R:s u	p->1	
RA ha	r->1	
REG, 	o->1	
REG-i	n->1	
REG?,	 ->1	
REP (	"->1	
REP r	e->1	
RINA 	h->1	v->1	
RINA,	 ->1	
RN) i	 ->1	
RNäst	a->1	
RPOL 	(->1	
RREG,	 ->1	
RREG-	i->1	
RREG?	,->1	
Rack 	o->1	
Rack,	 ->1	
Rafae	l->3	
Randz	i->4	
Rapka	y->11	
Rappo	r->3	
Rasch	h->1	
Rasis	m->1	
Readi	n->1	
Reakt	i->1	
Redan	 ->3	
Redin	g->8	
Refor	m->7	
Reger	i->6	
Regio	n->1	
Rent 	a->1	t->1	
Repub	l->1	
Reste	r->2	
Resul	t->5	
Retro	a->1	
Revid	e->1	
Revis	i->3	
Rhône	-->1	
Richa	r->1	
Richt	e->2	
Riis-	J->2	
Rika 	v->1	
Riktl	i->4	
Riofö	r->1	
Riske	n->1	
Rober	t->1	
Roble	s->1	
Roiss	y->1	
Rojos	 ->1	
Rom- 	o->1	
Romag	n->1	
Roman	o->2	
Román	,->1	
Roo f	r->1	
Ropet	 ->1	
Roth-	B->7	
Rotte	r->2	
Rover	 ->1	,->1	
Royal	 ->1	
Ruiz 	s->1	
Rumän	i->1	
Rush 	P->1	
Ryssl	a->4	
RÅDSK	A->1	
RÅGOR	N->1	
RÖSTN	I->2	
Räkna	 ->1	
Rätts	s->1	t->1	
Råder	 ->1	
Rådet	 ->14	,->2	s->4	
Rådso	r->1	
Réuni	o->2	
Rösta	 ->1	
S (In	t->1	
S och	 ->1	
S) - 	H->1	
S) är	 ->1	
S)) (	U->1	
S))(G	e->1	
S))(P	a->3	
S))..	(->1	
S)).J	a->1	
S))Fr	u->1	
S))oc	h->1	
S)].H	e->2	
S-zon	 ->1	e->2	
S:s p	a->1	
SA - 	o->1	
SA at	t->1	
SA el	l->1	
SA ha	r->1	
SA på	 ->1	
SA, K	a->1	
SA, s	o->1	
SA.Ja	g->1	
SA.Vi	 ->1	
SA:s.	L->1	
SD fö	r->1	
SE oc	h->2	
SE ti	l->1	
SE)Ja	g->1	
SE-gr	u->3	
SE-kr	i->3	
SE-te	s->1	
SEK (	d->1	
SEK(1	9->3	
SEK(9	9->1	
SEM-2	0->1	
SG, E	E->2	
SG-fö	r->6	
SKAND	E->1	
SOLAS	 ->1	
SP må	s->1	
SP oc	h->1	
SPA-i	n->1	
SPÖ o	c->1	
SPÖ) 	s->1	
SR - 	o->1	
SS oc	h->1	
SS:s 	p->1	
SSE t	i->1	
STNIN	G->2	
SU-gr	u->1	
SU:s 	E->1	e->1	
SYN))	.->1	
Sages	-->1	
Saint	-->1	
Salaf	r->1	
Samhä	l->2	
Samma	 ->4	n->22	
Samor	d->1	
Samti	d->14	
San S	e->1	
Sanni	n->5	
Sanno	l->1	
Santa	 ->1	
Sante	r->2	
Save 	(->2	m->1	ä->1	
Save,	 ->1	
Save-	 ->1	p->2	
SaveN	ä->1	
Schen	g->10	
Schre	y->3	
Schro	e->14	
Schrö	d->1	
Schul	z->3	
Schwa	r->1	
Schwe	i->1	
Schör	l->1	
Schüs	s->4	
Seatt	l->4	
Sebas	t->1	
Sedan	 ->19	,->1	
Segni	,->1	
Segur	o->1	
Seixa	s->5	
Seriö	s->1	
Sett 	u->1	
Shara	s->1	
Sharm	 ->4	-->1	
Sheik	.->1	h->4	
Shell	 ->2	
Sheph	e->3	
Simps	o->1	
Sist 	m->2	
Situa	t->3	
Sju ä	n->1	
Sjukh	u->1	
Själv	 ->1	k->1	
Sjätt	e->1	
Sjöst	e->4	
Skado	r->1	
Skall	 ->4	
Skogs	v->1	
Skott	l->5	
Skull	e->8	
Skydd	e->1	
Skäle	t->1	
Slova	k->1	
Slutl	i->34	
Slutr	e->1	
Sluts	a->3	
Små o	c->1	
Småfö	r->1	
Snabb	 ->1	
Snara	r->1	
Soare	s->1	
Socia	l->4	
Sokra	t->1	
Solan	a->4	
Solbe	s->2	
Som E	u->1	
Som T	h->1	
Som a	r->1	v->1	
Som b	e->1	
Som e	n->5	t->3	x->1	
Som f	ö->3	
Som h	ä->1	
Som j	a->8	
Som k	l->1	o->2	
Som l	e->1	ö->1	
Som m	e->1	
Som n	i->9	
Som p	a->1	o->2	
Som s	v->2	å->2	
Som t	i->1	
Som u	t->1	
Som v	i->2	o->1	
Somli	g->3	
Soula	d->1	
Spani	e->7	
Spenc	e->1	
Spero	n->1	
Sri L	a->3	
St.Va	l->1	
Stabi	l->1	
Stadg	a->1	
State	r->6	
Stati	s->1	
Statl	i->2	
Stock	h->3	
Stora	 ->2	
Storb	r->14	
Storm	a->2	
Straf	f->1	
Stras	b->5	
Strax	 ->1	
Struk	t->1	
Sträv	a->1	
Stämm	e->1	
Ståls	e->1	
Stöd 	m->1	s->1	t->1	
Stöde	n->1	r->2	
Stöds	y->1	
Störr	e->2	
Störs	t->2	
Suanz	e->1	
Subve	n->2	
Sudre	 ->1	,->1	
Svare	t->1	
Svepe	s->1	
Sveri	g->7	
Swobo	d->3	
Sydaf	r->2	
Sydko	r->1	
Sydos	t->2	
Syfte	t->6	
Syrie	n->22	r->2	
Sánch	e->1	
São T	o->2	
Säg m	i->1	
Säker	h->2	
Särsk	i->2	
Så bl	e->1	
Så de	t->3	
Så en	l->1	
Så er	a->1	
Så fr	å->1	
Så hä	r->1	
Så ja	g->3	
Så ka	n->1	
Så ko	m->1	
Så lä	n->3	
Så lå	n->1	t->1	
Så nå	g->1	
Så ri	k->1	
Så se	n->1	
Så so	m->2	
Så sä	g->1	
Så ti	d->1	
Så va	d->1	
Så vi	 ->2	l->1	s->1	
Så vå	r->1	
Så är	 ->1	
Så äv	e->2	
Sådan	 ->1	a->1	
Såled	e->4	
Sånge	n->1	
Såsom	 ->2	
Såväl	 ->1	
Söder	m->2	
T OM 	A->1	
T) De	n->1	
T) Ef	t->1	
T) Fr	å->1	
T) He	r->10	
T) Ja	g->2	
T) Le	d->1	
T) Nä	r->1	
T) Om	 ->1	
T) Vi	 ->1	
TCM.A	t->1	
TE ha	r->1	
TERRE	G->3	
TNING	(->1	.->1	
TO?En	d->1	
TT OM	 ->1	
TUELL	A->1	
TV an	k->1	
TV-bi	l->1	
TV-ka	n->1	
TV-pr	o->1	
TV-sä	n->1	
Ta dä	r->1	
Tacis	 ->1	-->1	
Tack 	f->9	s->15	
Tack,	 ->13	
Tack.	F->1	
Tadzj	i->5	
Taiwa	n->1	
Talar	 ->1	
Talma	n->9	
Tamme	r->22	
Tang 	o->1	
Tanio	;->1	
Tanke	n->3	
Tauer	n->1	
Terro	r->1	
Terró	n->3	
Tesau	r->1	
Texas	 ->2	
Theat	o->21	
Thyss	e->5	
Tibet	 ->12	"->2	,->3	-->1	.->2	?->1	
Tidig	a->1	
Tidni	n->1	
Till 	a->5	d->3	e->8	m->1	o->1	s->13	
Tills	a->2	
Tillv	e->2	ä->1	
Tillä	m->3	
Tillå	t->10	
Titta	 ->1	
Todin	s->1	
Tom S	p->1	
Tomé 	o->1	p->1	
Tongi	v->1	
Toppm	ö->2	
Torre	y->3	
Torv 	f->1	
Torve	n->1	
Total	 ->1	,->1	-->3	F->1	
Trans	i->1	p->2	
Tre ä	n->1	
Tredj	e->1	
Tritt	i->1	
Tror 	n->1	v->1	
Trots	 ->17	
Trovä	r->1	
Träd 	h->1	
Tsats	o->3	
Turki	e->35	
Turkm	e->2	
Tusen	 ->1	
Tvärt	 ->1	o->3	
Två v	i->1	
Två ä	n->1	
Ty en	l->1	
Ty ha	n->1	
Ty in	g->1	
Ty so	m->1	
Ty un	d->1	
Ty va	r->1	
Ty vi	 ->2	
Tycke	r->1	
Tydli	g->1	
Tyskl	a->20	
Tyvär	r->9	
Tänk 	b->1	p->1	
Tågkr	a->1	
U "co	u->1	
U I e	n->1	
U age	r->1	
U att	 ->2	
U bla	n->1	
U bör	 ->1	
U där	 ->1	
U fra	m->1	
U ger	 ->1	
U gör	 ->1	
U har	 ->2	
U i d	e->1	
U inf	ö->2	
U int	e->1	
U kan	 ->3	
U mer	 ->1	
U myc	k->1	
U mås	t->1	
U och	 ->4	
U på 	e->1	
U red	a->1	
U ska	l->1	
U som	 ->4	
U sys	s->1	
U uts	ä->1	
U utv	e->1	
U är 	r->1	v->1	
U, fö	r->1	
U, lå	t->1	
U, me	d->1	
U, nä	r->1	
U, på	 ->1	
U, ty	 ->1	
U, vi	l->1	
U-anp	a->1	
U-bis	t->1	
U-bud	g->1	
U-enh	e->1	
U-fon	d->1	
U-för	d->4	e->1	
U-gen	o->1	
U-gru	p->1	
U-ini	t->1	
U-ins	t->4	
U-kom	m->2	
U-kor	t->4	
U-kri	t->1	
U-lag	s->1	
U-lan	d->1	
U-län	d->3	
U-man	t->1	
U-med	b->4	e->1	
U-niv	å->1	
U-ord	f->1	
U-pro	g->2	
U-ram	p->1	
U-reg	e->1	
U-rät	t->1	
U-str	u->1	
U-sän	d->2	
U-tex	t->1	
U-utv	i->1	
U-vär	l->1	
U.. (	F->1	
U.All	a->1	
U.Dag	e->1	
U.De 	t->1	
U.Det	 ->1	
U.Frå	g->1	
U.Nu 	h->1	
U.Rop	e->1	
U.Vi 	g->1	s->1	v->1	
U:s B	a->1	
U:s E	u->1	
U:s b	e->1	i->2	u->2	y->1	
U:s d	o->1	
U:s e	g->1	u->1	
U:s f	r->1	ö->2	
U:s g	e->1	
U:s h	a->1	e->1	
U:s i	n->6	
U:s k	o->1	u->1	
U:s l	i->2	
U:s m	e->3	i->1	
U:s n	ä->1	
U:s o	c->3	m->1	r->2	
U:s p	o->3	
U:s r	e->1	
U:s s	t->4	
U:s t	e->1	j->1	
U:s u	r->1	
U?Her	r->1	
UCK n	u->1	
UCLAF	 ->1	
UE/NG	L->2	
UELLA	 ->1	
UEN-g	r->1	
UF) ä	r->1	
UGFJ)	 ->1	,->1	
UGFJ:	s->1	
UNIFI	L->1	
UNMIK	,->1	.->2	
USA -	 ->1	
USA a	t->1	
USA e	l->1	
USA h	a->1	
USA p	å->1	
USA, 	K->1	s->1	
USA.J	a->1	
USA.V	i->1	
USA:s	.->1	
USD f	ö->1	
USP o	c->1	
Ulste	r->1	
Undan	t->3	
Under	 ->34	
Ungdo	m->1	
Ungef	ä->2	
Union	e->8	
Uppda	t->1	
Uppen	b->1	
Uppfö	l->1	
Uppgi	f->3	
Upprä	t->1	
Ur de	n->2	
Ur en	 ->1	
Ur pa	r->1	
Urba-	,->1	
Urban	"->1	
Urqui	o->1	
Ursäk	t->1	
Utan 	e->1	t->1	v->1	
Utbil	d->2	
Utdel	n->1	
Utest	å->1	
Utfor	m->2	
Utför	a->1	
Utgif	t->2	
Utifr	å->1	
Utman	i->2	
Utnäm	n->2	
Utsko	t->6	
Uttjä	n->1	
Utvec	k->1	
Utvid	g->1	
Utvär	d->1	
Uzbek	i->2	
V - D	o->1	
V - R	e->1	
V ank	l->1	
V i E	G->1	
V i f	ö->1	
V-bil	d->1	
V-kan	a->1	
V-pro	g->1	
V-sän	d->1	
VC, a	t->1	
VC-le	k->1	
VC.Vi	 ->1	
VD bö	r->1	
VI i 	E->1	
VII:e	 ->1	
VIII 	h->1	k->1	
VIII:	e->1	
VP (Ö	s->2	
VP at	t->2	
VP mi	s->1	
VP) o	c->1	
Vad a	n->2	
Vad b	e->11	i->1	l->1	
Vad d	e->1	
Vad e	u->1	
Vad f	i->1	ö->1	
Vad g	ä->15	ö->1	
Vad h	ä->1	
Vad j	a->5	
Vad k	a->2	o->5	
Vad m	å->1	
Vad s	k->4	m->1	o->2	ä->2	
Vad t	r->1	ä->2	
Vad u	t->1	
Vad v	i->7	
Vad ä	r->6	
Vadan	 ->1	
Valde	z->3	
Valen	 ->1	t->1	
Valet	 ->1	
Valle	l->3	
Van H	u->3	
Vanda	m->1	
Vanli	g->1	
Vapen	 ->1	
Var d	e->1	
Var f	i->1	ö->1	
Var h	a->1	
Var o	c->2	
Var s	k->1	
Vare 	s->2	
Varel	a->1	
Varfö	r->12	
Varje	 ->7	
Varke	n->1	
Vatan	e->3	
Velze	n->1	
Vem b	e->2	
Vem d	i->1	
Vem k	o->1	
Vem s	k->2	
Vem v	i->1	
Vems 	a->1	t->1	
Vendé	e->1	
Venez	u->1	
Venst	r->2	
Verhe	u->2	
Verks	a->1	
Versa	i->1	
Veten	s->1	
Veter	a->1	
Vetsk	a->1	
Vi ac	c->1	
Vi al	l->1	
Vi an	s->16	v->1	
Vi ar	b->1	
Vi av	g->2	h->1	s->1	v->1	
Vi be	f->1	g->1	h->24	t->1	
Vi bi	d->1	
Vi bo	r->1	
Vi bö	r->11	
Vi de	l->2	
Vi di	s->5	
Vi dr	i->1	
Vi er	b->1	
Vi eu	r->1	
Vi fa	s->1	
Vi fi	c->2	n->1	
Vi fo	r->2	
Vi fä	s->1	
Vi få	r->14	
Vi fö	r->13	
Vi ge	r->1	
Vi gj	o->1	
Vi go	d->2	
Vi gr	a->1	
Vi gö	r->3	
Vi ha	d->4	r->87	
Vi ho	p->6	
Vi hy	s->1	
Vi hä	n->1	r->1	
Vi hå	l->2	
Vi i 	G->2	S->1	p->2	t->1	
Vi in	s->7	
Vi ja	g->1	
Vi ka	n->26	
Vi ko	m->21	
Vi kr	i->1	ä->7	
Vi ku	n->1	
Vi kä	n->4	
Vi la	d->2	
Vi li	t->1	
Vi lö	p->1	
Vi me	n->4	
Vi mi	n->1	
Vi mo	t->1	
Vi må	s->77	
Vi or	o->1	
Vi pa	r->1	
Vi pl	a->1	
Vi ra	d->1	
Vi re	s->1	
Vi ri	s->1	
Vi rä	k->2	
Vi rö	s->1	
Vi sa	t->1	
Vi se	r->6	
Vi si	k->1	
Vi sk	a->13	u->9	
Vi so	c->1	
Vi st	ä->2	å->2	ö->5	
Vi sv	a->2	e->1	
Vi sä	g->1	t->2	
Vi ta	c->1	l->3	r->1	
Vi ti	l->2	
Vi tr	o->3	
Vi tv	e->1	i->1	
Vi ty	c->3	s->1	
Vi tä	n->2	
Vi un	d->1	
Vi up	p->6	
Vi ut	e->1	g->1	
Vi va	r->5	
Vi ve	t->15	
Vi vi	d->1	l->29	s->1	
Vi vä	l->3	n->6	
Vi än	d->1	
Vi är	 ->34	
Vi ön	s->1	
Vi, d	e->1	
Via s	t->1	
Vichy	r->1	
Vid E	u->1	
Vid b	e->1	
Vid d	e->4	
Vid e	l->1	n->1	t->1	
Vid l	u->1	
Vid m	i->1	ö->1	
Vid s	i->2	
Vidar	e->7	
Vikte	n->1	
Vilja	n->1	
Vilka	 ->16	
Vilke	n->6	t->2	
Vill 	m->1	n->3	
Villk	o->1	
Vinde	n->1	
Vissa	 ->13	
Visse	r->2	
Visst	 ->1	
Vitbo	k->3	
Vitor	i->7	
Vivie	n->1	
Vlaam	s->1	
Vodaf	o->1	
Volks	w->1	
Von W	o->1	
Värde	n->1	
Värld	s->3	
Västb	a->4	
Västm	a->1	
Västr	a->1	
Vår d	j->1	
Vår e	g->1	
Vår g	e->1	r->4	
Vår i	d->1	n->1	
Vår o	r->1	
Vår r	o->1	ö->1	
Vår u	n->2	p->1	
Vår ö	n->1	
Våra 	e->1	f->2	l->1	m->2	r->1	ä->1	
Vårt 	f->1	m->2	p->2	s->1	u->1	
WTO?E	n->1	
Waffe	n->2	
Wales	 ->8	.->2	;->1	
Walls	t->4	
Washi	n->3	
Web, 	s->1	
West 	M->1	
Wide 	W->1	
Wiebe	n->1	
Wiela	n->4	
Wien 	f->1	o->2	
Wien,	 ->1	
Wilhe	l->1	
Wogau	 ->7	,->5	.->1	M->1	b->1	s->3	
World	 ->1	
Wulf-	M->2	
Wurtz	 ->2	,->1	
Wye P	l->1	
Wye-a	v->2	
Wynn,	 ->1	
X och	 ->2	
X, fa	s->1	
XVII:	e->1	
XVIII	:->1	
XXVII	:->1	I->1	
YN)).	 ->1	
Yasse	r->1	
York 	v->1	
Ytter	l->2	s->1	
Zeela	n->2	
Zimer	a->1	
[KOM(	1->2	
[SEK(	9->1	
].) H	e->1	
].Her	r->2	
a "Am	s->1	
a "ba	n->1	
a "ir	r->1	
a "lä	n->1	
a "sh	a->1	
a "ut	å->1	
a (KO	M->1	
a (ar	t->1	
a - a	t->1	v->2	
a - b	l->1	
a - d	e->7	
a - e	l->1	
a - f	i->1	r->2	ö->4	
a - g	ä->1	
a - h	a->1	u->1	
a - i	 ->2	n->1	
a - j	a->2	u->1	
a - k	a->1	o->1	
a - l	y->1	å->1	
a - m	a->1	e->3	i->1	å->1	
a - o	c->6	m->1	
a - p	a->1	å->2	
a - r	a->1	e->2	ö->1	
a - s	a->1	k->1	o->1	t->1	å->1	
a - t	a->1	
a - u	t->1	
a - v	i->1	
a - ä	r->2	
a -, 	f->1	
a 1 o	c->2	
a 1 p	r->1	
a 10 	p->1	ä->1	
a 100	 ->1	
a 123	 ->1	
a 125	 ->1	
a 133	.->1	
a 15 	å->1	
a 16 	o->1	p->1	
a 167	 ->1	
a 170	 ->1	
a 2 p	r->1	u->1	
a 200	0->1	
a 25 	p->4	
a 250	 ->1	
a 30 	m->1	
a 33 	o->1	
a 35 	m->1	
a 370	 ->1	
a 40 	p->1	
a 5 m	i->1	
a 55 	p->1	
a 6 o	c->1	
a 60 	0->1	
a 70 	a->1	
a 81 	o->4	
a 81.	1->1	
a 85 	o->2	t->1	
a 87,	 ->1	
a 90-	t->1	
a Ahe	r->1	
a Ale	x->1	
a Ali	c->1	
a Alt	e->1	
a Ams	t->1	
a Atl	a->1	
a Azo	r->1	
a B o	c->1	
a Bal	k->1	
a Bar	a->1	c->1	
a Ber	e->1	n->1	
a Bow	i->1	
a Bry	s->2	
a Col	a->1	
a Cos	t->8	
a Dal	a->1	
a Dan	m->1	
a EEG	 ->1	
a EG-	d->1	k->4	
a EU 	b->1	i->2	m->1	
a EU-	f->1	i->2	m->1	p->1	r->1	s->1	
a EU:	s->4	
a Eli	s->1	
a Ell	e->1	
a Eri	k->2	
a Eur	o->56	
a Eva	n->1	
a FN:	s->2	
a FPÖ	 ->2	
a Fei	r->1	
a Fis	c->1	
a Fla	u->1	
a Flo	r->2	
a Flé	c->1	
a Fra	n->4	
a För	i->1	
a Gol	a->1	
a Gra	ç->1	
a Gro	s->1	
a Hai	d->5	
a Han	s->1	
a Hic	k->1	
a Hul	t->1	
a IX 	o->1	
a Int	e->1	
a Isr	a->2	
a Izq	u->1	
a Jan	-->1	
a Jea	n->1	
a Jer	u->1	
a Jon	c->1	
a Jör	g->2	
a Kar	l->1	
a Koc	h->2	
a Kos	o->1	
a Kou	c->1	
a Kun	g->1	
a Lan	g->1	
a Lib	a->3	
a Lii	k->1	
a Loi	r->1	
a Lou	s->1	
a Maa	s->1	
a Mal	t->1	
a Mar	i->1	
a Mel	l->1	
a Mou	r->8	s->1	
a Mul	d->1	
a Nan	a->1	
a Nat	i->1	
a Nie	l->1	
a OLA	F->1	
a PPE	-->1	
a PVC	-->1	
a Pak	i->1	
a Pal	a->1	e->2	
a Poe	t->2	
a Pro	d->1	
a Rac	k->1	
a Rii	s->1	
a Rob	e->1	
a Rom	á->1	
a Rot	t->1	
a Rys	s->1	
a Réu	n->2	
a Sal	a->1	
a Sav	e->1	
a Sch	r->1	
a She	l->1	
a Sta	t->1	
a Sua	n->1	
a Sve	r->1	
a TV-	s->1	
a Ter	r->1	
a Tex	a->1	
a Tur	k->2	
a Tys	k->2	
a UCK	 ->1	
a Wal	e->1	
a Zee	l->2	
a abs	o->3	
a adj	e->1	
a adm	i->4	
a aff	ä->3	
a age	r->5	
a agg	r->1	
a akt	 ->1	i->7	ö->5	
a ald	r->1	
a alk	e->1	
a all	 ->2	a->22	i->2	m->15	t->22	v->3	
a alt	e->5	
a amb	i->8	
a an 	t->1	
a ana	l->3	
a anb	l->1	
a and	a->2	r->34	
a anf	ö->2	
a ang	e->3	r->1	å->2	
a anh	ä->2	
a ank	l->1	
a anl	e->2	ä->1	
a anm	ä->4	
a ann	a->2	
a ano	r->2	
a anp	a->1	
a ans	a->1	e->5	j->1	l->4	t->21	v->39	å->1	ö->2	
a ant	a->6	i->3	y->1	
a anv	ä->28	
a app	l->2	
a ara	b->1	
a arb	e->75	
a arg	u->7	
a arm	é->2	
a arr	a->2	o->1	
a art	i->11	
a arv	.->1	e->2	
a asp	e->17	
a asy	l->2	
a atl	a->1	
a ato	m->4	
a att	 ->470	,->2	.->1	i->3	
a auk	t->1	
a aut	o->1	
a av 	E->5	F->2	K->1	T->1	a->10	b->7	d->59	e->11	f->9	g->3	h->4	i->3	k->4	l->1	m->9	n->1	o->6	p->4	r->1	s->9	t->4	u->6	v->10	y->1	ä->3	å->1	ö->1	
a av,	 ->2	
a av.	D->1	
a ava	n->1	
a avd	e->2	
a avf	a->1	
a avg	ö->2	
a avl	ä->1	
a avs	a->1	e->19	i->6	k->1	l->4	n->2	t->7	
a avt	a->15	
a avv	i->1	
a bak	g->9	o->1	
a bal	a->2	
a ban	k->1	n->1	o->2	
a bar	a->5	n->3	r->1	
a bas	 ->1	,->1	e->2	k->1	
a be 	e->3	h->1	k->1	p->1	
a bea	k->1	
a beb	y->1	
a bed	r->9	ö->5	
a bef	i->1	o->21	r->2	ä->1	
a beg	r->11	ä->8	å->2	
a beh	a->14	o->9	å->1	ö->7	
a bek	l->4	r->2	v->3	y->4	ä->1	
a bel	g->1	o->5	y->1	ä->1	
a bem	a->1	ä->2	
a ber	e->2	i->1	o->2	ä->1	ö->3	
a bes	i->1	l->44	t->52	v->2	ä->1	ö->2	
a bet	a->4	e->1	o->8	r->8	u->1	y->20	ä->70	
a beu	n->1	
a bev	a->1	i->17	
a bib	e->1	l->2	
a bid	r->18	
a bie	f->2	
a bil	a->37	b->1	d->3	e->1	i->7	k->3	p->2	s->3	t->5	v->2	
a bin	d->2	
a bis	t->2	
a bit	 ->1	
a bju	d->1	
a bl.	a->1	
a bla	n->3	
a bli	 ->8	r->15	v->2	
a bo 	k->1	
a bol	a->3	
a bom	b->1	
a bor	d->11	t->7	
a bos	t->2	
a bot	 ->2	
a bra	 ->3	.->1	n->1	
a bri	s->8	t->1	
a bro	a->1	m->1	t->8	
a bru	t->2	
a brä	n->3	
a brå	d->2	
a bud	g->19	o->1	s->4	
a byg	g->7	
a byr	å->4	
a bär	 ->1	a->2	s->1	
a bäs	t->2	
a bät	t->7	
a båd	a->4	e->2	
a båt	a->2	e->1	
a bör	 ->14	d->3	j->8	s->1	
a can	c->1	
a cen	t->10	
a cer	t->4	
a cha	n->4	r->1	
a cit	e->1	
a civ	i->1	
a da 	F->1	
a dag	 ->3	.->1	a->6	e->3	o->7	
a dam	e->38	
a dan	s->1	
a dat	a->2	o->1	u->1	
a de 	8->1	P->2	a->8	b->7	d->4	e->13	f->18	g->6	h->7	i->5	j->1	k->4	l->6	m->15	n->11	o->8	p->6	r->10	s->22	t->6	u->5	v->3	y->2	ä->5	å->4	ö->5	
a deb	a->42	
a dec	e->2	
a def	i->3	
a del	 ->19	,->1	a->22	e->23	f->1	r->1	s->1	t->3	u->2	
a dem	 ->47	,->2	.->8	:->1	a->2	o->22	
a den	 ->132	)->1	,->2	.->9	;->1	n->63	s->1	
a dep	a->1	
a der	a->8	
a des	a->2	s->66	
a det	 ->140	!->1	,->9	.->9	a->4	s->1	t->73	
a dia	l->9	
a die	k->1	
a dif	f->3	
a dig	 ->2	
a dik	e->1	t->1	
a dil	e->1	
a dim	e->9	
a dip	l->4	
a dir	e->48	
a dis	c->2	k->16	p->1	t->1	
a dju	p->2	r->5	
a dog	.->1	
a dok	u->16	
a dom	a->3	i->1	s->11	
a dra	 ->1	b->4	g->6	s->1	
a dri	f->1	v->4	
a dro	g->1	
a dru	c->1	
a drö	m->1	
a dub	b->2	
a dum	p->1	t->1	
a dyn	a->1	
a dyr	 ->1	a->2	
a där	 ->10	,->1	.->3	f->4	m->2	
a då 	b->1	d->2	i->1	o->1	
a dål	i->1	
a död	a->1	s->1	
a döm	a->1	
a dör	r->2	
a döt	t->1	
a eff	e->26	
a eft	e->23	
a ege	t->1	
a egn	a->26	
a ego	i->1	
a eko	l->1	n->33	
a ekv	a->1	
a ele	m->4	
a eli	m->1	
a ell	e->48	
a elv	a->1	
a eme	l->5	
a emo	t->12	
a en 	"->1	a->16	b->18	c->4	d->16	e->29	f->21	g->20	h->14	i->8	j->3	k->29	l->9	m->21	n->10	o->7	p->10	r->20	s->41	t->15	u->13	v->14	ä->1	å->3	ö->6	
a en,	 ->1	
a ena	d->2	
a enb	a->1	
a end	a->4	
a ene	r->44	
a eng	e->2	
a enh	e->9	ä->3	
a eni	g->1	
a enk	e->2	l->1	
a enl	i->7	
a eno	r->2	
a ens	 ->1	e->1	k->2	
a env	i->2	
a er 	-->1	a->7	e->3	f->4	h->1	i->1	k->2	m->1	o->10	p->1	t->2	u->6	
a er,	 ->4	
a era	 ->5	
a erb	j->4	
a erf	a->10	o->2	
a eri	n->2	
a erk	ä->2	
a ers	ä->2	
a ert	 ->1	
a eta	b->2	p->1	
a etc	.->1	?->1	
a etn	i->3	
a ett	 ->178	
a eur	o->35	
a eve	n->3	
a exa	k->2	
a exe	m->10	
a exi	l->1	s->1	
a exp	e->1	l->1	o->2	
a ext	e->1	r->6	
a fak	t->11	
a fal	l->54	
a fam	i->4	
a fan	n->1	t->2	
a far	h->1	l->3	o->2	s->1	t->20	v->5	
a fas	,->1	t->13	
a fat	t->8	
a fel	 ->1	a->2	
a fem	 ->4	t->1	å->2	
a fen	o->1	
a fil	m->1	o->1	
a fin	a->11	n->9	s->1	
a fis	k->8	
a fla	g->1	
a fle	r->10	s->1	x->3	
a fli	c->1	
a flo	t->1	
a fly	k->2	
a flö	d->1	
a fog	a->1	
a fol	k->32	
a fon	d->10	
a for	a->1	d->38	m->14	s->7	t->13	u->1	
a fos	s->1	
a fot	b->1	
a fra	m->114	n->2	s->1	
a fre	d->5	
a fri	 ->1	-->2	a->2	g->1	h->6	s->2	v->4	
a fro	n->1	
a fru	 ->3	k->4	
a frä	m->2	
a frå	g->235	n->52	
a ful	l->7	
a fun	d->2	g->5	k->3	n->1	
a fus	i->2	
a fyr	a->1	
a fär	d->1	
a fäs	t->1	
a få 	b->1	d->1	e->2	f->1	h->1	l->1	m->2	o->1	p->1	s->3	v->1	
a fåg	e->1	l->2	
a fån	g->2	
a får	 ->18	
a föd	d->1	e->1	o->1	
a föl	j->30	
a för	 ->345	,->5	.->1	b->28	d->17	e->159	f->20	h->31	i->1	k->4	l->13	m->3	n->10	o->5	p->9	r->4	s->139	t->15	u->13	v->21	ä->21	å->1	ö->1	
a gal	e->1	l->1	
a gam	l->3	m->2	
a gan	s->2	
a gar	a->11	
a gav	 ->1	
a ge 	b->2	e->4	g->1	o->1	s->1	
a gem	e->65	
a gen	a->1	e->4	o->44	t->3	u->1	
a geo	s->1	
a ger	 ->2	
a ges	 ->1	
a gic	k->1	
a gif	t->1	
a gig	a->1	
a gil	t->4	
a giv	a->10	e->1	
a gjo	r->6	
a gla	d->1	
a glä	d->3	
a glö	m->2	
a gnä	l->1	
a god	 ->1	a->10	k->2	t->2	
a gra	d->5	n->4	t->11	
a gre	k->2	
a gro	g->1	
a gru	n->34	p->57	
a gry	m->1	
a grä	n->17	
a grö	n->1	
a gäc	k->1	
a gäl	l->27	
a gär	n->2	
a gå 	f->1	u->1	
a gån	g->40	
a går	 ->5	
a gör	 ->6	.->1	a->27	s->1	
a ha 	e->5	h->1	n->1	r->1	s->1	y->1	
a had	e->8	
a haf	t->1	
a hal	v->2	
a ham	n->8	
a han	d->65	s->3	t->4	
a hap	p->1	
a har	 ->108	,->1	m->2	
a hat	e->1	
a hav	e->2	s->2	
a hel	a->10	h->2	s->1	t->15	
a hem	l->3	m->1	
a hen	n->7	
a her	r->6	
a het	e->1	
a hin	d->14	
a his	t->7	
a hit	 ->1	,->1	t->3	
a hjä	l->4	r->2	
a hom	o->1	
a hon	o->12	
a hop	p->4	
a hor	i->1	
a hos	 ->6	
a hot	 ->2	e->1	
a hum	ö->1	
a hun	d->2	
a hur	 ->29	.->2	u->3	
a hus	 ->1	,->1	
a huv	u->5	
a hyl	l->1	
a hyp	o->1	
a hys	a->1	
a häf	t->1	
a häl	f->1	s->3	
a hän	d->15	s->33	v->4	
a här	 ->9	,->2	
a häv	d->3	
a hål	l->19	
a hår	d->1	k->1	t->1	
a håv	a->1	
a hög	 ->1	a->3	e->3	r->1	s->9	t->2	
a höj	d->1	
a höl	l->1	
a hör	 ->1	a->4	t->2	
a i A	m->2	
a i B	r->1	
a i C	a->1	e->3	
a i D	a->3	
a i E	C->1	G->1	U->1	u->47	
a i F	a->1	i->1	ö->1	
a i G	o->1	
a i I	r->2	
a i K	o->5	
a i L	i->1	o->2	u->1	
a i M	a->1	
a i P	P->1	o->2	
a i R	o->1	y->1	
a i S	t->1	
a i T	a->1	h->1	i->2	u->1	
a i U	E->1	
a i W	a->1	
a i a	l->5	n->1	r->4	t->2	
a i b	e->3	i->1	r->1	
a i d	a->7	e->81	i->2	
a i e	k->1	n->19	r->2	t->11	x->1	
a i f	a->1	l->1	o->1	r->19	u->1	ö->7	
a i g	e->5	o->2	r->1	å->1	
a i h	a->3	e->3	u->1	
a i i	n->3	
a i j	u->1	
a i k	o->11	r->6	v->1	
a i l	a->4	i->2	
a i m	a->1	e->4	i->9	o->2	å->2	ö->1	
a i n	i->1	ä->2	
a i o	c->2	l->1	m->4	
a i p	a->2	e->1	o->1	r->3	
a i r	a->1	e->1	ä->1	å->2	
a i s	a->5	e->1	i->4	j->1	k->1	l->2	o->1	t->5	y->3	ä->1	å->2	
a i t	.->1	a->1	e->1	i->1	v->1	
a i u	n->7	t->3	
a i v	a->4	e->2	i->4	ä->2	å->8	
a i y	r->1	t->1	
a i Ö	s->6	
a i ä	n->1	
a i å	t->1	
a i ö	s->1	v->2	
a i.D	e->1	
a i.N	ä->1	
a i.S	e->1	
a iak	t->2	
a ibl	a->1	
a ick	e->2	
a ide	a->2	n->3	o->1	
a idé	 ->4	e->3	n->3	
a ifa	l->1	
a ifr	å->4	
a ige	n->9	
a ign	o->1	
a igå	n->3	
a ihj	ä->1	
a iho	p->3	
a ihå	g->14	
a ika	p->1	
a ill	a->1	e->1	
a ima	g->1	
a imm	i->1	
a imp	o->1	u->2	
a in 	a->1	b->2	d->4	f->1	h->1	i->4	k->1	l->1	m->1	o->2	p->3	r->2	s->3	u->2	v->4	y->1	
a in,	 ->1	
a inb	j->1	l->2	
a inc	i->3	
a ind	i->6	u->9	
a inf	e->1	l->1	o->12	r->3	ö->10	
a ing	r->2	
a inh	e->1	
a ini	t->24	
a ink	l->2	o->2	ö->1	
a inl	e->3	ä->10	
a inn	a->2	e->23	o->1	
a ino	m->25	
a inr	i->3	ä->3	
a ins	a->21	i->1	l->2	p->1	t->70	y->2	
a int	e->78	o->1	r->53	
a inv	a->4	e->6	i->1	ä->3	å->1	
a irr	a->1	
a iso	l->1	
a isä	r->2	
a itu	 ->14	
a ive	r->1	
a ja,	 ->1	
a jag	 ->5	
a job	b->3	
a jor	d->14	
a jul	k->1	
a jur	i->6	
a jus	t->2	
a jäm	f->2	n->1	s->4	v->1	
a jär	n->1	
a kal	l->1	
a kam	m->24	p->7	
a kan	 ->51	a->1	d->1	s->3	
a kap	a->1	i->3	
a kar	a->5	t->3	
a kat	a->16	o->2	
a ked	j->2	
a kil	o->1	
a kin	e->1	
a kl.	 ->1	
a kla	p->1	r->17	s->2	u->1	
a kli	b->1	e->1	m->5	
a klo	c->1	
a kly	f->3	
a kna	p->1	
a kno	w->1	
a knu	t->1	
a kny	t->2	
a koa	l->1	
a kod	 ->2	e->1	
a kok	o->1	
a kol	-->1	l->101	
a kom	 ->1	m->217	p->12	
a kon	c->3	f->13	k->79	s->47	t->44	v->3	
a kop	p->1	
a kor	,->1	r->7	t->7	
a kos	t->24	
a kra	f->10	v->24	
a kre	a->2	t->3	
a kri	g->5	n->1	s->10	t->13	
a kro	p->1	
a krä	n->2	v->5	
a krå	n->1	
a kul	t->14	
a kun	d->3	n->7	s->3	
a kur	s->1	
a kus	t->14	
a kva	l->11	r->8	
a kvi	n->14	
a kvo	t->3	
a kvä	l->1	
a kyl	a->1	
a käl	l->3	
a kän	d->1	n->7	s->5	
a kär	a->4	l->2	n->11	
a köl	a->1	
a köp	 ->1	
a lab	o->2	
a lad	e->1	
a lag	 ->1	a->5	f->1	l->1	o->1	s->17	t->1	
a lan	d->20	
a lar	m->1	v->1	
a led	a->25	d->1	e->2	n->4	
a leg	i->1	
a lek	e->1	
a lev	a->4	n->1	
a lib	e->9	
a lig	g->9	
a lik	a->12	g->1	n->1	s->1	
a lin	j->3	
a lis	t->2	
a lit	a->1	e->7	
a liv	,->3	e->7	s->17	
a lju	g->1	s->1	
a lob	b->1	
a lok	a->10	
a lov	y->1	
a luc	k->2	
a lug	n->1	
a lyc	k->1	
a lyf	t->1	
a lys	s->3	
a läg	e->4	g->6	r->1	
a läk	a->1	
a läm	n->6	p->6	
a län	d->67	g->3	
a lär	d->5	
a läs	t->1	
a lät	t->3	
a lån	g->4	
a låt	e->1	
a löf	t->6	
a lön	 ->1	t->2	
a löp	t->1	
a lös	a->4	n->16	
a maj	o->6	
a mak	r->1	t->4	
a man	 ->5	d->7	
a mar	g->1	i->1	k->26	
a mas	k->2	s->2	
a mat	e->8	
a max	i->1	
a med	 ->223	,->3	.->1	b->59	d->13	e->30	f->4	g->2	i->4	l->80	v->11	
a meg	a->1	
a mek	a->3	
a mel	l->21	
a men	 ->10	i->6	
a mer	 ->14	,->1	.->2	a->1	
a mes	t->3	
a met	a->1	o->7	
a mig	 ->19	,->1	.->1	?->1	r->1	
a mik	r->1	
a mil	j->29	l->1	
a min	 ->14	,->1	a->11	d->5	i->11	n->6	o->5	s->2	u->1	
a mis	s->12	t->1	ä->1	
a mit	t->23	
a mob	i->2	
a mod	 ->1	e->11	i->2	
a mom	s->1	
a mon	o->8	
a mor	d->1	
a mot	 ->19	,->1	i->2	p->2	s->5	t->1	å->2	
a mun	t->2	
a mur	a->1	
a mus	i->1	
a myc	k->46	
a myg	g->1	
a myn	d->55	
a mäk	t->1	
a män	g->3	n->21	s->2	
a mär	k->2	
a mät	t->1	
a mål	 ->20	,->5	.->7	e->15	s->8	
a mån	a->15	d->1	g->8	
a mås	t->62	
a måt	t->2	
a möd	r->1	
a möj	l->57	
a mör	d->1	
a möt	a->1	e->6	
a nai	v->1	
a nam	n->2	
a nar	k->1	
a nat	i->39	u->4	
a ned	 ->5	l->1	s->2	
a neg	a->2	
a nej	 ->1	
a neo	n->1	
a ner	e->1	
a ni 	g->1	h->2	ä->1	
a nim	b->1	
a nio	 ->2	
a niv	å->14	
a nog	 ->1	.->1	a->1	g->1	
a non	 ->2	
a nor	m->8	
a not	a->1	
a nr 	1->2	2->2	3->10	4->7	5->1	6->1	7->1	8->1	9->1	
a nu 	n->1	
a nu?	J->1	
a nul	l->1	
a nun	n->1	
a nuv	a->1	
a ny 	o->1	
a nya	 ->29	,->1	
a nyc	k->3	
a nyh	e->5	
a nyl	i->1	
a nyt	t->5	
a nyå	r->1	
a näm	n->13	
a när	 ->26	a->1	i->2	m->3	v->3	
a näs	t->4	
a nät	 ->2	v->8	
a nå 	f->1	ä->1	
a någ	o->47	r->31	
a nåt	t->1	
a nöd	b->1	v->8	
a nöj	a->2	d->1	
a nöt	t->1	
a oav	s->1	
a oba	l->4	
a obe	f->1	g->1	r->4	s->1	
a obl	i->3	
a och	 ->537	,->2	
a ock	s->20	
a odd	s->1	
a odu	g->1	
a oeg	e->2	
a oen	i->1	
a ofe	l->1	
a off	e->7	i->1	r->5	
a ofr	å->1	
a oft	a->2	
a ofö	r->2	
a oge	n->1	
a oin	t->1	
a ojä	m->2	
a okl	a->3	
a oko	n->1	
a oli	k->15	
a olj	a->1	e->7	
a oly	c->10	
a olö	s->1	
a om 	-->2	2->1	3->1	B->1	E->1	F->1	G->1	I->2	K->1	L->1	S->1	T->3	a->46	b->7	d->49	e->15	f->22	g->3	h->8	i->8	j->3	k->19	l->5	m->14	n->5	o->5	p->4	r->6	s->11	t->2	u->7	v->14	ä->1	å->2	ö->2	
a om,	 ->6	
a om.	D->2	J->2	
a omb	u->5	
a ome	d->2	
a omf	a->9	
a omg	å->2	
a omr	å->89	ö->4	
a oms	t->31	
a omv	ä->3	
a omö	j->1	
a ond	a->1	
a onö	d->2	
a opa	r->1	
a ope	r->4	
a opi	n->1	
a opp	o->1	
a opt	i->2	
a ord	 ->20	,->2	a->2	e->9	f->82	n->6	
a ore	a->1	
a org	a->32	
a ori	e->1	k->1	m->1	
a oro	 ->1	,->1	.->3	l->1	n->1	s->2	
a ors	a->8	
a ort	.->1	
a orä	t->1	
a oss	 ->61	,->2	.->1	
a osä	k->1	
a oti	l->1	
a pak	e->1	
a pal	e->1	
a par	a->5	l->84	t->41	
a pas	s->1	
a pat	i->1	
a ped	a->1	
a pek	a->1	
a pel	a->2	
a pen	g->18	n->3	s->1	
a per	i->6	s->17	
a pes	t->1	
a pht	a->1	
a pir	a->1	
a pla	n->21	s->1	t->5	
a ple	n->1	
a plä	d->1	
a pol	i->82	
a pop	u->1	
a por	t->1	
a pos	i->6	
a pra	k->3	t->1	x->5	
a pre	c->3	f->3	j->1	m->1	s->10	
a pri	c->1	n->30	o->9	s->3	v->3	
a pro	b->58	c->19	d->6	f->2	g->61	j->22	p->2	t->4	v->5	
a prö	v->1	
a pub	l->1	
a pum	p->1	
a pun	d->2	k->76	
a på 	A->1	B->2	E->2	G->1	a->26	b->5	d->31	e->25	f->6	g->13	h->3	k->3	l->4	m->9	n->8	o->3	p->3	r->5	s->16	t->9	u->2	v->16	ä->4	
a på,	 ->4	
a på.	U->1	Ä->2	
a på:	 ->1	
a påf	ö->1	
a påg	å->2	
a påm	i->5	
a påp	e->9	
a pås	t->4	
a påt	r->1	
a påv	e->1	
a rad	i->5	
a ram	 ->2	e->6	p->3	v->2	
a ran	d->12	
a rap	p->38	
a rea	k->9	l->2	
a red	a->9	o->4	u->2	
a ref	l->1	o->32	
a reg	e->94	i->65	l->32	
a rek	o->8	
a rel	a->5	e->1	
a ren	o->2	s->3	t->2	
a rep	r->4	u->4	
a res	e->2	o->28	p->10	t->2	u->50	
a ret	o->1	
a rev	i->5	
a rig	o->1	
a rik	a->1	e->2	t->37	
a rim	l->1	
a ris	k->18	
a ro,	 ->1	
a rol	l->6	
a rom	e->1	
a rub	r->1	
a rum	 ->17	.->2	
a run	d->2	t->1	
a rut	i->4	
a ryg	g->1	
a räc	k->1	
a räd	d->5	s->1	
a räk	e->1	n->3	
a rät	t->87	
a råd	 ->5	.->1	a->1	e->30	g->3	s->4	
a råo	l->1	
a råt	t->1	
a rör	 ->4	a->3	d->1	e->2	l->10	
a rös	t->11	
a röt	t->2	
a s.k	.->1	
a sad	e->4	
a sag	t->1	
a sak	 ->13	.->1	e->14	f->1	n->2	o->1	
a sam	a->14	f->5	h->12	m->66	o->7	r->2	s->1	t->13	v->2	
a san	k->2	n->2	t->1	
a sat	s->3	t->1	
a sce	n->4	
a se 	a->3	d->2	m->1	t->1	
a sed	a->6	
a seg	e->1	
a sei	s->1	
a sek	e->2	r->3	t->28	u->2	
a sen	a->5	
a ser	 ->4	
a ses	s->2	
a set	t->4	
a sex	 ->2	
a sid	a->35	o->6	
a sif	f->8	
a sig	 ->109	,->3	.->6	n->2	
a sim	u->1	
a sin	 ->29	a->46	
a sit	t->19	u->40	
a sju	k->1	n->3	
a sjä	l->10	t->4	
a sjö	f->4	m->2	n->2	
a ska	d->10	l->54	m->1	n->2	p->9	t->12	
a ske	 ->1	d->2	p->3	r->2	t->2	
a ski	c->1	l->26	p->1	s->2	
a skj	u->1	
a sko	g->4	l->5	
a skr	a->1	i->3	o->5	ä->2	
a sku	l->31	t->1	
a sky	d->7	l->3	
a skä	l->20	r->1	
a skö	t->1	v->1	
a sla	g->17	
a slu	t->25	
a slä	k->1	
a slå	 ->2	r->1	
a smu	s->1	t->1	
a små	 ->8	f->1	g->1	s->1	
a sna	b->8	r->2	
a sne	d->2	
a snä	l->1	
a soc	i->37	
a sol	i->4	
a som	 ->215	,->3	m->1	
a sor	t->1	
a spa	r->1	
a spe	c->17	g->1	k->3	l->10	
a spo	n->1	
a spr	å->2	
a spä	n->3	r->1	
a spå	r->1	
a spö	k->2	
a sta	b->1	c->1	d->7	n->8	t->53	
a ste	g->9	n->1	
a sti	c->2	m->2	
a sto	l->3	p->6	r->24	
a str	a->16	i->4	u->23	y->1	ä->5	å->1	ö->5	
a stu	d->9	n->1	
a sty	c->1	r->5	
a stä	l->25	m->1	
a stå	 ->1	l->6	n->58	r->6	
a stö	d->86	r->14	t->1	
a sub	j->1	s->4	v->2	
a sum	m->7	
a sut	t->1	
a suv	e->1	
a sva	g->1	r->9	
a svå	n->1	r->20	
a syd	e->1	
a syf	t->8	
a sym	b->2	p->1	
a syn	 ->2	d->1	e->1	n->1	o->1	p->10	s->3	v->2	
a sys	s->17	t->32	
a säg	a->25	e->8	s->1	
a säk	e->16	r->2	
a säm	r->1	
a sän	d->4	
a sär	s->8	
a säs	o->1	
a sät	t->65	
a så 	a->13	b->2	f->2	h->3	k->2	l->1	m->3	n->1	o->1	s->1	t->1	v->4	
a så.	I->1	O->1	
a såd	a->11	
a såg	 ->1	
a sån	g->2	
a sås	o->2	
a såv	ä->1	
a sön	e->1	
a sör	j->1	
a t.o	.->2	
a ta 	d->2	f->1	h->2	m->1	s->1	t->1	u->10	
a tac	k->15	
a tag	 ->2	i->3	
a tak	e->1	
a tal	 ->3	.->1	a->12	e->3	
a tan	k->13	
a tar	 ->5	v->1	
a tas	 ->4	
a tax	e->1	
a tea	t->1	
a tec	k->3	
a tek	n->9	
a tel	e->1	
a tem	a->1	p->1	
a ten	d->6	
a ter	m->3	r->8	
a tex	t->18	
a tid	.->2	e->16	i->3	n->1	p->1	s->8	t->1	
a tig	e->1	
a til	l->328	
a tim	m->2	
a tin	g->1	
a tio	t->1	
a tit	t->1	
a tjä	n->26	r->1	
a tog	 ->3	s->3	
a tol	e->3	k->2	
a tom	m->1	
a ton	 ->1	g->1	v->2	
a tor	s->1	v->2	
a tot	a->4	
a tox	i->1	
a tra	d->8	f->1	g->2	n->14	v->1	
a tre	 ->15	d->1	t->1	
a tri	o->1	
a tro	 ->1	j->1	l->1	r->1	t->1	v->2	
a tru	p->1	s->2	
a try	c->1	g->2	
a trä	d->3	n->1	s->1	t->1	
a trå	d->2	
a trö	s->1	
a tun	g->2	n->1	
a tur	e->1	
a tus	e->2	
a tvi	n->3	s->3	v->2	
a två	 ->25	n->1	
a tyc	k->6	
a tyd	e->1	l->8	
a tyn	g->4	
a typ	 ->11	.->2	e->4	g->1	
a tys	k->2	
a täc	k->1	
a tän	k->4	
a täv	l->1	
a tåg	k->1	
a tål	a->1	
a ult	r->1	
a umg	ä->1	
a und	a->15	e->45	g->1	v->3	
a ung	a->1	d->1	e->2	
a uni	l->1	o->268	v->1	
a upp	 ->108	.->4	b->1	d->3	e->1	f->14	g->25	h->3	l->2	m->18	n->2	r->5	s->6	t->5	v->1	
a ur 	b->1	d->1	e->3	m->3	t->1	
a ura	n->1	
a urh	o->1	
a urs	k->2	ä->2	
a urv	a->1	
a ut 	b->1	d->4	e->4	f->1	h->2	i->2	m->2	n->1	o->1	p->2	r->1	t->1	u->1	ö->1	
a ut.	J->2	
a ut:	 ->1	
a uta	n->19	r->1	
a utb	a->1	i->5	u->1	y->2	
a ute	s->2	
a utf	l->1	o->6	ö->3	
a utg	i->5	j->1	å->4	ö->3	
a uth	ä->1	
a uti	f->1	
a utk	a->13	
a utl	ä->3	
a utm	a->6	ä->4	
a utn	y->4	
a utr	e->2	i->1	u->1	
a uts	e->1	k->9	l->5	t->3	ä->2	
a utt	a->8	j->3	o->1	r->7	
a utv	e->54	i->10	ä->7	
a utö	v->1	
a vac	k->2	
a vad	 ->28	
a vag	n->1	
a vak	s->2	
a val	 ->5	,->1	.->2	;->1	d->2	e->3	f->1	k->1	r->1	u->6	
a van	 ->6	o->1	
a vap	e->6	n->2	
a var	 ->27	.->1	a->13	d->1	f->2	i->11	j->6	k->1	m->1	n->4	s->1	t->2	
a vat	t->1	
a vec	k->21	
a ved	e->1	
a vel	a->1	
a vem	 ->1	
a ven	t->1	
a ver	b->1	k->61	s->7	
a vet	 ->5	a->5	e->3	
a vi 	d->1	g->1	k->2	n->1	s->1	t->2	ä->1	ö->1	
a vic	e->3	
a vid	 ->17	a->7	d->2	g->1	h->1	
a vik	t->38	
a vil	d->1	j->18	k->13	l->41	
a vin	d->2	s->4	
a vir	k->1	
a vis	 ->1	a->11	d->1	e->1	i->1	s->19	
a vit	b->5	
a von	 ->2	
a vor	e->2	
a vot	e->2	
a vra	k->2	
a väd	e->1	j->2	
a väg	.->1	a->3	e->5	l->3	r->3	
a väk	t->1	
a väl	 ->4	.->1	d->2	f->1	g->1	j->5	k->3	
a vän	n->2	s->3	
a vär	d->19	l->21	s->2	
a väs	e->5	
a väv	n->2	t->1	
a väx	e->4	t->1	
a våg	 ->1	l->1	
a vål	d->4	
a vår	 ->17	,->1	a->15	t->13	
a yrk	e->3	
a ytl	i->1	
a ytt	e->11	r->4	
a Öst	e->6	
a äga	r->6	
a ägd	e->1	
a äge	r->1	
a ägn	a->1	
a ägt	 ->1	
a ämb	e->3	
a ämn	a->1	e->16	
a än 	i->3	s->1	
a änd	a->6	p->1	r->88	
a änn	u->7	
a änt	l->3	
a är 	E->1	a->28	b->4	d->30	e->78	f->17	g->3	h->4	i->18	j->2	k->3	l->6	m->16	n->15	o->11	p->3	r->4	s->17	t->11	u->3	v->14	ä->1	å->1	ö->2	
a är,	 ->3	
a är.	D->1	E->1	F->1	
a är:	 ->2	
a ära	d->1	
a äre	n->4	
a ärl	i->2	
a äve	n->10	
a å m	i->2	
a åkl	a->8	
a år 	2->1	a->2	f->4	i->1	k->1	s->5	t->2	
a år,	 ->7	
a år.	D->1	F->1	J->1	V->2	
a åre	n->2	t->22	
a årh	u->2	
a årl	i->2	
a års	 ->1	b->1	t->1	
a årt	a->1	
a åsa	m->1	
a åsi	k->5	
a åsk	å->1	
a åst	a->2	
a åt 	i->1	s->1	
a åt.	K->1	
a åta	 ->1	g->14	l->7	
a åte	r->22	
a åtf	ö->1	
a åtg	ä->99	
a öar	 ->1	n->2	
a öde	s->2	
a öga	t->1	
a ögo	n->5	
a öka	d->4	n->1	r->2	s->1	
a ökn	i->2	
a öns	k->7	
a öpp	e->4	n->2	
a öre	 ->1	
a öro	n->1	
a öst	e->4	l->1	u->1	
a öve	r->80	
a övr	i->2	
a! De	t->1	
a! Vi	 ->1	
a!Av 	d->1	
a!Den	 ->1	
a!Det	 ->3	
a!Fru	 ->3	
a!För	e->1	
a!Her	r->2	
a!Jag	 ->1	
a!Låt	 ->1	
a!Män	n->1	
a!Om 	n->1	
a!Äve	n->1	
a" bi	l->1	
a" so	m->1	
a" va	r->1	
a", v	i->1	
a".. 	(->1	
a".Ba	r->1	
a".De	s->1	t->1	
a".Hi	s->1	
a".Ju	s->1	
a".Ki	n->1	
a"; ö	v->1	
a"ind	i->1	
a) ad	 ->1	
a) bä	t->1	
a, 16	7->1	
a, 50	 ->1	
a, Br	o->1	
a, Ev	a->1	
a, Ja	p->1	
a, Kv	ä->1	
a, Sa	m->1	
a, Sc	h->1	
a, ad	e->1	
a, al	l->3	
a, an	g->1	s->1	
a, ar	b->2	
a, at	t->24	
a, av	 ->3	s->1	
a, ba	r->1	
a, be	t->1	
a, bi	d->1	l->1	
a, bl	.->3	a->2	
a, bo	r->1	
a, bå	d->1	
a, co	m->1	
a, de	 ->11	m->3	n->7	s->2	t->13	
a, dj	u->2	
a, dv	s->6	
a, dä	r->6	
a, då	 ->3	
a, dö	d->1	
a, ef	t->12	
a, ek	o->1	
a, el	l->4	
a, en	 ->6	e->2	h->1	l->2	
a, er	a->1	
a, et	t->5	
a, eu	r->1	
a, ex	a->1	
a, fo	r->1	
a, fr	a->5	e->1	u->4	ä->2	å->1	
a, fu	l->1	
a, få	r->2	
a, fö	r->38	
a, ga	r->1	
a, ge	d->1	n->2	
a, gö	r->1	
a, ha	d->1	n->1	r->12	
a, he	l->1	r->13	
a, hj	ä->1	
a, hu	m->1	r->2	s->1	v->1	
a, hö	g->2	
a, i 	a->3	b->1	d->3	e->2	f->1	i->1	j->1	m->1	r->1	s->9	
a, ib	l->1	
a, in	g->1	k->1	n->1	o->2	t->10	
a, ja	g->3	
a, jo	r->1	
a, ju	s->2	
a, ka	n->6	t->1	
a, ko	m->5	n->3	o->1	
a, le	m->1	
a, li	k->6	
a, lä	g->1	
a, lå	n->2	t->1	
a, me	d->9	n->38	s->1	
a, mi	l->3	n->1	
a, mo	r->1	
a, må	s->4	
a, na	t->2	
a, ne	d->1	j->1	
a, nu	 ->1	
a, ny	a->1	
a, nä	m->2	r->6	
a, nå	g->4	
a, oa	v->1	
a, ob	e->1	
a, oc	h->86	k->1	
a, om	 ->16	
a, or	g->1	
a, pa	r->1	
a, pe	r->1	
a, pr	e->2	i->2	
a, på	 ->3	p->1	
a, ra	s->2	
a, re	a->1	g->6	
a, ri	k->1	
a, rä	t->2	
a, sa	m->5	
a, se	 ->1	r->1	
a, sk	a->2	u->1	
a, sl	ä->1	
a, sn	a->1	
a, so	c->3	m->43	
a, st	a->1	o->1	r->2	å->1	
a, sv	å->1	
a, sä	g->1	r->3	
a, så	 ->12	d->1	s->6	v->1	
a, sö	k->1	
a, t.	e->1	
a, ta	r->1	
a, te	o->1	
a, ti	l->10	
a, tj	ä->1	
a, to	r->1	
a, tr	e->1	o->4	
a, tu	l->1	
a, ty	 ->1	
a, tö	m->1	
a, un	d->2	i->1	
a, up	p->1	
a, ut	a->18	f->1	g->1	o->1	v->1	
a, va	d->4	r->4	
a, ve	r->2	
a, vi	 ->7	d->1	k->1	l->24	s->2	
a, vo	r->1	
a, vä	g->1	
a, äg	a->1	
a, är	 ->8	
a, äv	e->4	
a, åt	e->1	f->1	g->1	m->1	
a, öp	p->1	
a, öv	e->1	
a-, S	a->1	
a-Isr	a->1	
a-Rom	a->1	
a-oly	c->1	
a. 12	0->1	
a. De	t->2	
a. Dä	r->1	
a. Då	 ->1	
a. En	l->1	
a. Fö	l->1	
a. Hå	l->1	
a. Ja	g->1	
a. Ko	m->1	
a. Kä	r->1	
a. Me	n->3	
a. So	m->1	
a. Va	r->2	
a. ar	t->1	
a. at	t->1	
a. be	t->1	
a. de	s->1	
a. en	 ->1	
a. et	t->1	
a. få	r->1	
a. fö	r->4	
a. ge	n->1	
a. gö	r->1	
a. i 	M->1	p->1	
a. kr	i->1	
a. me	d->1	
a. nä	r->3	
a. ol	j->1	
a. om	 ->1	
a. på	 ->1	
a. sk	a->2	
a. st	o->1	
a. un	d->1	
a. va	d->1	
a. Åt	g->1	
a.(Ih	å->1	
a.(Pa	r->1	
a.(Ta	l->2	
a.)Be	t->1	
a.)Fr	u->1	
a.- (	P->4	
a.. H	e->1	
a.. T	a->1	
a..(E	N->1	
a..(I	T->1	
a..(N	L->1	
a...(	T->1	
a...L	å->1	
a.18 	m->1	
a.All	a->4	t->6	
a.Ams	t->1	
a.Ann	a->2	
a.Ans	e->1	
a.Av 	a->1	d->3	v->1	
a.Bak	o->2	
a.Ber	e->1	o->1	
a.Bes	l->2	
a.Bet	ä->1	
a.Bil	l->1	
a.Bla	n->1	
a.Bor	d->1	
a.Cor	p->1	
a.De 	f->3	g->1	o->1	p->1	s->2	
a.Den	 ->18	n->6	
a.Des	s->9	
a.Det	 ->92	t->22	
a.Doc	k->1	
a.Där	 ->1	e->2	f->11	
a.Då 	h->1	k->1	
a.EG-	d->1	
a.Eft	e->8	
a.Eme	l->3	
a.En 	a->2	f->2	k->2	m->1	s->1	u->1	
a.Enk	e->1	
a.Enl	i->3	
a.Ett	 ->8	
a.Eur	o->4	
a.Fac	k->2	
a.Fra	m->1	
a.Fru	 ->4	
a.Frå	g->3	
a.Föl	j->1	
a.För	 ->19	e->2	l->1	s->3	
a.Gem	e->1	
a.Ger	 ->1	
a.Giv	e->1	
a.Han	d->1	s->1	
a.Hel	t->1	
a.Her	r->33	
a.Hul	t->1	
a.Hur	 ->3	
a.Här	 ->4	
a.I E	u->1	
a.I a	l->1	
a.I b	e->1	
a.I d	a->1	e->5	i->1	
a.I e	n->2	
a.I f	r->3	ö->2	
a.I l	i->4	
a.I m	o->1	
a.I p	a->1	r->2	
a.I r	e->2	
a.I s	l->1	å->1	
a.I t	j->1	
a.I v	ä->1	å->1	
a.I ö	v->1	
a.Ibl	a->2	
a.Ing	e->1	
a.Ino	m->3	
a.Int	e->3	
a.Jag	 ->98	
a.Jus	t->2	
a.Kaf	o->1	
a.Kan	s->1	
a.Kom	m->9	p->1	
a.Kon	k->2	
a.Kär	a->1	n->1	
a.Lik	s->1	
a.Liv	s->1	
a.Läg	g->1	
a.Låt	 ->6	
a.Maj	o->1	
a.Man	 ->3	
a.Med	 ->7	a->1	b->1	l->2	
a.Men	 ->27	
a.Min	 ->3	a->6	n->1	
a.Mån	g->2	
a.Nat	i->1	u->1	
a.Ni 	a->1	b->1	f->1	h->1	k->1	m->1	
a.Nu 	k->1	ä->2	
a.När	 ->10	
a.Och	 ->9	
a.Om 	a->1	d->1	e->1	m->2	n->1	p->1	v->4	
a.Ord	f->1	
a.Ors	a->1	
a.Par	l->1	
a.Per	s->1	
a.Pre	c->2	
a.Pro	g->1	j->1	
a.På 	a->1	d->6	e->1	o->1	s->2	
a.Reg	i->1	
a.Res	u->1	
a.Rum	ä->1	
a.Råd	e->2	
a.Sam	t->1	
a.Sed	a->2	
a.Sit	u->2	
a.Sju	 ->1	
a.Sky	d->1	
a.Slu	t->3	
a.Små	f->1	
a.Som	 ->6	
a.Sta	t->1	
a.Stö	d->1	r->1	
a.Syf	t->1	
a.Säg	 ->1	
a.Så 	e->1	l->1	s->1	
a.Sån	g->1	
a.Tac	k->2	
a.Tad	z->1	
a.Til	l->2	
a.Top	p->1	
a.Tro	t->5	
a.Ty 	v->1	
a.Und	e->3	
a.Ung	d->1	
a.Upp	g->2	
a.Ur 	e->1	
a.Uta	n->1	
a.Utb	i->1	
a.Utd	e->1	
a.Utf	o->1	
a.Utn	ä->1	
a.Vad	 ->10	
a.Var	 ->1	e->1	j->1	
a.Vem	s->1	
a.Ver	k->1	
a.Vi 	a->2	b->9	d->1	f->1	g->1	h->17	i->1	k->7	l->2	m->11	r->1	s->5	t->4	u->4	v->6	
a.Via	 ->1	
a.Vid	 ->1	a->3	
a.Vik	t->1	
a.Vil	l->1	
a.Vis	s->2	
a.Vär	d->1	
a.Väs	t->1	
a.Vår	 ->1	a->2	
a.Än 	e->1	
a.Änd	r->1	
a.Änt	l->1	
a.Är 	d->2	k->1	
a.Äve	n->5	
a.Å a	n->2	
a.År 	1->1	
a.Öve	r->1	
a/Eur	o->1	
a/hal	v->1	
a/sam	m->1	
a: "D	e->1	
a: "i	n->1	
a: De	 ->1	
a: Fö	r->2	
a: I 	b->1	s->1	
a: Ja	g->2	
a: Nä	r->1	
a: Va	d->1	
a: Ve	m->1	
a: an	t->1	
a: at	t->1	
a: de	 ->1	
a: ge	n->1	
a: hu	r->2	
a: ma	n->1	
a: om	 ->1	
a: rä	t->1	
a: sk	a->1	
a: un	d->1	
a: up	p->1	
a: ut	b->1	
a: ve	m->2	
a: vi	 ->2	l->1	
a: Äv	e->1	
a:För	o->1	
a; de	t->1	
a; en	 ->1	
a; fö	r->2	
a; ja	g->2	
a; ko	m->1	
a; lo	j->1	
a; oc	h->1	
a; pu	n->1	
a; vi	 ->2	
a?"Ja	 ->1	
a?. (	E->1	
a?Ans	e->1	
a?Avs	l->1	
a?De 	h->1	
a?Den	 ->1	
a?Det	 ->6	
a?Ett	 ->1	
a?Fru	 ->1	
a?För	 ->1	
a?Har	 ->1	
a?Her	r->1	
a?Hur	 ->1	
a?I F	r->1	
a?I d	a->1	
a?Ini	t->1	
a?Jag	 ->3	
a?Jo,	 ->1	
a?Man	 ->1	
a?Nej	,->1	
a?När	 ->1	
a?Pro	b->1	
a?På 	v->1	
a?Sva	r->1	
a?Vad	 ->3	
a?Vi 	s->2	
a?Vil	k->1	
a?Vis	s->1	
a?Är 	d->1	
aHerr	 ->1	
aNäst	a->2	
aaffä	r->1	
aams 	B->1	
aan f	ö->1	
aan.V	a->1	
aans 	b->4	m->1	
aarde	r->1	
aastr	i->6	
ab sk	a->1	
abaré	b->1	
abase	n->1	
abb h	j->1	
abb o	c->2	
abb v	a->1	
abba 	b->2	f->1	o->2	p->1	r->1	t->1	u->1	v->1	å->1	
abbad	e->27	
abbar	 ->3	e->11	
abbas	 ->7	t->3	
abbat	 ->3	s->9	
abbt 	f->5	g->2	h->1	k->3	l->1	m->2	o->1	p->1	s->14	t->1	u->1	v->2	
abbt,	 ->3	
abbt.	J->1	M->1	O->2	T->1	V->1	
abbva	r->1	
abeha	n->7	
abekä	m->1	
abel 	H->1	P->1	i->1	n->1	r->1	
abel!	M->1	
abel,	 ->3	
abel.	D->1	V->2	Ä->1	
abell	 ->4	.->2	
abelt	 ->11	.->8	;->1	?->1	
aberg	e->1	
abete	r->1	
abeth	 ->1	
abil 	g->1	o->1	
abila	 ->1	r->1	
abili	s->3	t->16	
abilt	 ->2	
abine	t->3	
abise	n->1	
abisk	 ->1	-->1	a->4	
abla 	d->1	e->1	f->1	i->2	s->3	t->1	
abla"	.->1	
abla,	 ->1	
abla.	M->1	N->1	Ö->1	
ablan	c->1	
abler	a->11	i->2	
ablon	m->1	
abock	"->1	a->1	
abon 	f->1	g->1	k->1	m->1	
abon,	 ->1	
abon.	V->1	
abonm	ö->2	
abora	t->3	
abrep	u->1	
abrie	n->3	
abrik	e->1	
absol	u->40	
absor	b->1	
absta	t->2	
abstr	a->1	
absur	d->1	t->2	
abu i	n->1	
abukt	e->2	
abula	r->1	
abvär	l->1	
ac bl	i->1	
ac bö	r->1	
ac os	v->1	
ac", 	f->1	
ac-sy	s->1	
aca M	o->3	
aca s	a->1	
acao 	t->1	
accep	t->88	
ace o	c->1	
ace.D	e->1	
ace.J	a->1	
acera	 ->4	d->5	s->2	t->4	
aceri	n->2	
aceut	i->1	
acill	 ->1	
acio 	V->3	f->1	h->1	s->2	
acio,	 ->3	
acio.	J->1	N->1	
acio:	 ->1	
acios	 ->2	
acis 	f->1	
acis-	p->1	
acite	t->5	
ack a	t->1	
ack f	r->2	ö->9	
ack g	å->2	
ack h	a->1	
ack m	o->1	
ack o	c->4	
ack p	å->1	
ack s	o->1	ä->1	å->15	
ack t	i->11	
ack v	a->7	
ack, 	f->5	h->6	k->4	
ack-p	o->1	
ack.F	r->1	
ack.H	e->1	
ack.J	a->1	
acka 	A->1	G->2	K->2	L->1	P->2	S->1	a->5	d->4	e->4	f->21	h->7	i->1	k->11	l->3	m->4	o->3	p->3	r->3	u->1	v->5	
ackar	 ->20	s->1	
ackat	 ->2	s->1	
ackde	l->8	
acken	 ->1	
acker	t->2	
ackfö	r->7	
ackla	.->1	s->1	
ackni	n->6	
ackor	 ->1	
ackra	 ->5	s->1	
acks 	u->1	
acksa	m->9	
ackso	n->2	
aco-a	f->1	
acob 	S->2	
acque	s->3	
acqui	s->1	
actor	t->1	
acète	 ->1	
ad - 	ä->1	
ad Ad	e->1	
ad BN	I->1	
ad Eu	r->1	
ad FP	Ö->1	
ad Gu	i->1	
ad Ku	l->2	
ad Sy	r->1	
ad al	l->1	
ad an	a->1	s->4	t->1	v->4	
ad ar	g->1	
ad at	t->16	
ad av	 ->18	s->1	
ad be	h->2	s->5	t->24	
ad bi	l->1	n->1	
ad bl	i->1	o->1	
ad bo	m->1	
ad by	g->1	
ad da	g->4	
ad de	 ->7	l->1	m->1	n->5	s->1	t->16	
ad do	k->2	m->1	
ad då	 ->1	
ad ef	t->2	
ad el	e->1	l->4	
ad en	 ->2	e->4	
ad er	 ->1	
ad et	t->1	
ad eu	r->2	
ad fe	d->1	
ad fi	n->1	
ad fl	e->1	
ad fo	r->2	
ad fr	a->1	å->4	
ad fö	r->23	
ad ge	n->1	r->1	
ad gi	l->1	
ad gr	u->2	
ad gä	l->60	
ad gö	r->1	
ad ha	n->4	r->1	
ad ho	c->2	
ad hä	l->1	n->2	
ad i 	L->1	a->1	b->2	d->1	e->2	f->3	h->1	m->1	o->1	å->1	
ad id	é->1	
ad im	p->1	
ad in	f->6	r->1	s->4	t->1	
ad ja	g->12	
ad ju	r->1	
ad jä	m->1	
ad ka	n->5	
ad ko	m->16	n->10	r->1	
ad kr	i->1	
ad kv	a->1	
ad le	d->1	
ad ma	i->1	j->6	n->9	t->1	
ad me	d->4	l->4	n->1	
ad mi	l->2	
ad mo	t->1	
ad må	s->3	
ad na	m->1	t->1	
ad ni	 ->3	,->1	
ad nå	g->1	
ad oc	h->11	
ad ol	i->2	
ad om	 ->21	f->1	
ad or	d->1	
ad pa	r->1	
ad pe	r->1	
ad po	l->4	
ad pr	e->1	i->1	o->1	
ad pu	n->1	
ad på	 ->9	
ad re	a->1	f->1	v->1	
ad ri	k->1	
ad ro	l->2	
ad rä	d->1	t->3	
ad rå	d->1	
ad sa	k->1	m->2	
ad se	d->1	k->1	r->1	
ad si	t->3	
ad sk	a->3	e->1	r->1	u->1	
ad sm	å->2	
ad sn	e->1	
ad so	c->1	m->66	
ad st	a->1	r->1	y->1	å->1	ö->1	
ad su	b->1	
ad sy	s->8	
ad sä	g->2	k->2	
ad ta	g->1	
ad ti	d->1	l->12	
ad tj	ä->1	
ad tr	a->1	o->1	
ad tä	n->2	
ad un	d->1	
ad up	p->1	
ad ur	s->1	
ad ut	v->4	
ad va	n->1	
ad ve	r->2	t->5	
ad vi	 ->24	d->1	l->1	
ad vo	n->1	
ad vå	r->3	
ad yr	k->1	
ad än	 ->1	
ad är	 ->11	e->1	
ad äv	e->1	
ad öp	p->1	
ad öv	e->18	
ad, "	a->1	
ad, a	t->2	
ad, e	f->1	n->1	
ad, f	ö->1	
ad, h	a->1	
ad, i	 ->1	n->1	
ad, m	e->3	
ad, o	c->1	
ad, s	k->1	p->1	
ad, t	r->1	y->1	
ad, u	p->1	
ad, v	i->1	
ad, ä	v->1	
ad-ko	s->1	
ad."M	e->1	
ad.(S	a->1	
ad.De	t->7	
ad.Eu	r->1	
ad.Fr	å->1	
ad.He	r->6	
ad.Ja	g->4	
ad.Ko	m->2	
ad.Me	n->4	
ad.Mä	n->1	
ad.Må	n->1	
ad.Om	r->14	
ad.Pa	r->1	
ad.Re	g->1	
ad.Su	b->1	
ad.Ut	a->1	
ad.Ve	t->1	
ad.Vi	l->1	s->1	
ad: e	n->1	
ad; d	e->1	
ad?Dä	r->1	
ad?He	r->1	
ad?Vi	 ->1	
ada E	u->1	
ada d	e->4	
ada e	r->1	
ada f	i->1	
ada k	o->1	
ada o	c->1	
ada r	i->1	
ada s	o->1	
ada ö	v->2	
ada!D	e->1	
ada, 	J->1	e->1	r->1	
ada.M	e->1	
adade	s->2	
adaga	s->1	
adaki	s->1	
adan 	d->1	
adan.	D->1	
adana	 ->2	
adar 	a->1	d->1	g->1	j->1	m->2	
adat.	F->1	
adats	,->2	.->1	
addad	 ->1	
adde 	j->1	m->1	
adder	 ->1	
addin	g->2	
addit	i->1	
ade "	f->1	l->2	
ade -	 ->3	
ade 1	9->2	
ade 2	0->1	
ade 4	0->1	
ade E	u->4	
ade F	r->1	
ade H	a->1	e->1	o->1	
ade I	r->1	
ade N	a->1	
ade O	i->1	
ade T	u->1	
ade V	a->1	
ade a	d->1	g->1	m->1	n->9	r->8	t->28	v->14	
ade b	e->13	i->4	l->1	r->4	y->1	å->2	
ade d	a->3	e->28	i->2	o->1	ä->1	å->1	ö->1	
ade e	f->2	k->1	l->1	m->2	n->13	t->3	
ade f	a->5	i->2	l->4	r->9	u->3	y->1	å->2	ö->25	
ade g	e->3	j->2	l->1	o->3	r->1	å->2	
ade h	a->7	e->5	o->1	ä->1	å->1	ö->1	
ade i	 ->35	n->18	
ade j	a->13	o->1	
ade k	a->6	i->1	l->1	o->25	r->5	u->23	
ade l	e->6	ä->1	
ade m	a->9	e->13	i->3	o->3	u->1	y->2	ä->6	å->11	ö->1	
ade n	i->3	o->1	y->5	ä->2	å->2	
ade o	c->21	e->1	l->1	m->41	r->2	s->3	v->1	
ade p	a->8	e->7	l->2	o->1	r->9	å->9	
ade r	a->1	e->20	i->1	ä->3	å->3	
ade s	a->5	e->3	i->11	k->5	l->1	n->1	o->3	t->14	u->1	v->3	y->8	ä->3	å->1	
ade t	.->1	a->1	i->25	j->1	r->3	y->1	
ade u	n->5	p->1	r->4	t->6	
ade v	a->10	e->4	i->21	o->1	ä->2	å->2	
ade y	r->1	
ade Ö	s->1	
ade ä	g->1	n->1	r->4	
ade å	t->7	
ade ö	n->2	v->4	
ade, 	a->2	b->1	d->2	e->1	h->2	i->2	k->1	m->3	n->3	o->6	s->2	v->1	ö->1	
ade. 	O->1	V->1	
ade.A	t->1	v->1	
ade.D	e->6	ä->1	
ade.E	n->2	
ade.F	ö->2	
ade.H	e->2	u->1	
ade.J	a->2	
ade.M	e->1	
ade.P	r->1	
ade.S	l->2	o->2	å->1	
ade.T	V->1	o->1	r->1	
ade.V	i->2	
ade: 	k->1	
ade?J	a->1	
adeer	s->2	
adefo	n->1	
adeir	a->2	
adekv	a->5	
adels	 ->2	
ademi	,->1	n->1	
ademo	k->2	
aden 	-->2	a->16	b->2	d->1	e->1	f->11	g->2	h->2	i->6	l->1	m->6	o->13	p->3	r->1	s->7	t->1	u->1	v->1	ä->8	
aden)	(->2	.->1	
aden,	 ->29	
aden.	 ->1	.->2	A->2	D->6	E->1	F->2	I->2	J->3	K->1	M->2	O->1	P->1	S->2	U->1	V->4	
adens	 ->17	i->2	
ader 	-->1	I->2	a->2	d->1	e->5	f->5	i->3	k->4	l->3	m->5	o->11	p->7	r->1	s->11	u->2	v->1	
ader,	 ->12	
ader-	p->1	
ader.	 ->1	A->1	D->7	I->1	J->3	N->1	O->1	U->2	V->1	
ader;	 ->1	
adera	 ->2	.->1	s->1	
adern	a->81	
aders	 ->1	p->2	
ades 	-->1	1->2	2->1	S->1	V->1	a->16	d->5	e->3	f->13	g->1	h->4	i->18	k->4	m->5	n->1	o->9	p->1	s->5	t->9	u->4	v->3	
ades,	 ->5	
ades.	)->1	D->1	J->1	M->2	U->1	
adest	å->1	
adet 	s->1	u->1	
adet.	D->1	
adga 	f->4	k->1	m->1	o->2	p->1	s->2	ä->2	ö->1	
adga,	 ->1	
adgad	e->1	
adgan	 ->9	.->1	
adgar	 ->1	.->1	
adgor	 ->1	
adiet	 ->3	.->1	
adika	l->16	
ading	 ->1	
adins	t->1	
adiol	o->2	
aditi	o->19	
adium	 ->3	.->1	
adiz 	e->1	f->2	
adiz,	 ->1	
adiz-	k->1	
adjek	t->2	
adkom	m->24	
adlig	 ->2	a->5	t->3	
adlin	e->1	
admin	i->25	
admiu	m->3	
ado, 	a->1	
ador 	d->1	f->1	o->1	p->2	s->5	u->1	v->1	
ador,	 ->4	
ador.	H->1	M->1	
adorn	a->8	
adou 	f->1	
adox,	 ->1	
adoxa	l->5	
adrag	a->3	
adria	t->1	
adrid	 ->1	,->1	.->1	
ads b	e->1	
ads- 	o->1	
ads-i	n->2	
ads-n	y->1	
ads/i	n->1	
adsak	t->1	
adsan	d->3	
adsar	b->1	
adsbe	f->5	
adsce	n->1	
adsdo	m->1	
adsef	f->4	
adsek	o->14	
adsfr	i->4	
adsfö	r->1	
adsin	s->1	t->2	
adskr	a->1	
adsli	b->1	
adslå	n->1	
adsmy	n->1	
adsmö	j->1	
adsni	v->1	
adsom	r->1	
adsor	g->1	
adspr	i->1	o->5	
adsst	a->3	
adsti	l->1	
adsup	p->1	
adsve	r->1	
adsvi	l->2	
adt, 	O->1	
advis	 ->3	
advok	a->5	
adzji	k->5	
adör 	M->1	
ael -	 ->1	
ael a	t->3	v->1	
ael b	e->1	
ael d	r->1	
ael f	å->1	ö->1	
ael h	i->1	
ael i	n->1	
ael l	ö->1	
ael m	å->1	
ael o	c->10	
ael v	e->1	
ael, 	k->1	m->1	n->1	ö->1	
ael-S	y->1	
ael.D	e->1	ä->1	
ael.N	ä->1	
ael.S	a->1	
ael?E	l->1	
aeler	 ->1	n->4	
aelis	k->15	
aelkr	i->1	
aels 	e->1	p->2	s->1	v->1	å->1	
af om	 ->1	
afael	 ->2	.->1	
afats	 ->1	
afety	-->1	
aff o	c->2	
aff, 	p->1	
aff- 	o->2	
affa 	a->3	b->1	d->1	e->4	f->3	k->3	m->1	r->1	s->2	u->1	
affad	e->3	
affan	d->1	
affar	 ->1	
affas	 ->3	
affat	.->1	
affbe	s->1	
affen	 ->1	-->1	s->1	
affla	g->1	
affpr	o->2	
affrä	t->28	
affär	e->11	s->1	
afi p	å->1	
afi.D	e->1	
afi.V	i->1	
afik 	s->1	ä->1	
afik-	 ->1	
afik.	B->1	D->1	
afike	n->3	
afikl	e->1	
afin.	V->1	
afisk	 ->2	a->6	t->2	
aflyk	t->1	
afone	-->1	
afor 	o->1	
afran	c->1	
afrik	a->2	
afryt	t->2	
afråg	a->2	o->10	
aft 2	0->1	
aft a	l->1	t->2	v->3	
aft b	e->2	
aft d	e->3	ä->1	
aft e	n->1	t->2	x->1	
aft f	a->1	l->1	r->1	ö->6	
aft h	a->1	
aft i	 ->3	n->1	
aft k	a->1	
aft m	e->2	y->1	å->1	ö->1	
aft n	ä->2	å->2	
aft o	c->3	m->1	
aft p	r->2	å->2	
aft s	a->1	e->1	i->1	k->2	o->2	t->3	v->1	å->2	
aft t	a->1	i->3	
aft u	n->1	t->1	
aft v	i->1	ä->1	å->1	
aft ä	r->1	
aft, 	S->1	f->1	m->3	o->1	s->2	u->1	v->2	
aft.D	e->1	ä->1	
aft.H	e->1	
aft.M	e->1	
aft.V	i->2	
aft? 	M->1	
aft?N	e->1	
aften	 ->13	,->1	.->3	
after	 ->4	,->2	.->2	n->1	
aftfu	l->12	
aftig	 ->9	,->1	a->14	t->10	
afton	e->1	
aftsa	n->4	
aftso	l->1	
aftsp	l->1	r->1	
aftsr	e->1	
aftss	ä->1	
aftsv	e->1	
aftta	g->1	
afttr	ä->4	
aftve	r->8	
ag - 	d->2	j->1	m->1	o->4	s->1	t->1	ä->1	
ag 1 	m->1	o->1	
ag 1,	 ->1	2->1	
ag 10	 ->4	.->1	
ag 11	,->1	
ag 12	 ->1	
ag 13	 ->1	
ag 15	 ->1	
ag 17	 ->1	
ag 18	 ->2	
ag 19	 ->2	9->1	
ag 2,	 ->2	
ag 22	 ->1	,->2	
ag 23	 ->1	
ag 26	 ->1	
ag 3 	o->1	
ag 34	 ->1	
ag 38	 ->2	:->1	
ag 4 	o->1	
ag 4.	I->2	
ag 43	 ->1	
ag 44	 ->1	
ag 45	.->3	
ag 5,	 ->2	
ag 6 	o->2	
ag Ga	z->1	
ag IN	T->1	
ag ab	s->1	
ag ac	c->2	
ag al	l->3	
ag an	s->89	t->4	v->1	
ag at	t->87	
ag av	 ->12	r->2	s->5	t->1	v->2	
ag ba	d->2	r->7	
ag be	 ->3	a->1	f->4	g->3	h->2	k->14	r->22	t->8	u->1	
ag bi	d->1	
ag bl	e->5	i->3	
ag bo	r->1	
ag bö	r->4	
ag ci	t->2	
ag de	 ->3	l->7	n->4	t->4	
ag do	c->3	
ag dr	a->2	o->1	
ag dä	r->5	
ag då	 ->1	
ag dö	r->1	
ag ef	t->2	
ag el	l->1	
ag em	e->3	o->3	
ag en	 ->10	b->1	d->1	
ag er	 ->7	,->1	h->1	i->2	k->2	
ag et	t->3	
ag fa	s->1	
ag fi	c->2	n->3	
ag fo	r->5	
ag fr	a->14	å->37	
ag fu	l->1	n->1	
ag få	r->8	t->3	
ag fö	r->109	
ag ga	n->1	r->1	v->1	
ag ge	 ->2	n->2	r->5	
ag gi	c->1	
ag gj	o->2	
ag gl	a->2	ä->8	
ag go	d->1	
ag gr	a->9	u->1	
ag gä	l->3	r->7	
ag gå	r->1	
ag gö	r->2	
ag ha	 ->1	d->3	n->1	r->110	
ag he	d->1	l->7	n->1	
ag hi	n->1	
ag ho	p->54	t->1	
ag hu	r->1	
ag hä	l->2	n->1	r->9	v->4	
ag hå	l->14	
ag hö	l->1	r->6	
ag i 	B->1	E->2	F->1	I->1	K->2	S->2	T->2	a->3	b->1	d->13	e->6	f->6	m->1	p->1	s->3	u->2	v->3	
ag i,	 ->1	
ag in	 ->1	d->1	f->4	g->5	k->1	n->3	o->3	s->14	t->55	v->1	
ag ja	g->1	
ag ju	 ->1	s->1	
ag jä	m->1	
ag ka	m->1	n->64	
ag kl	.->2	a->2	
ag ko	l->1	m->39	n->3	
ag kr	a->1	
ag ku	n->2	
ag kä	n->10	
ag kö	p->1	
ag la	d->1	g->2	n->1	
ag le	d->2	g->1	
ag li	k->1	t->2	
ag ly	f->2	s->5	
ag lä	g->3	m->1	s->2	
ag lå	t->1	
ag lö	s->1	
ag ma	n->1	
ag me	d->20	n->7	r->3	
ag mi	g->14	n->6	s->1	
ag mo	t->4	
ag my	c->4	
ag mä	r->1	
ag må	h->1	s->22	
ag na	t->5	
ag ni	 ->2	
ag no	g->1	l->1	t->3	
ag nu	 ->5	m->1	
ag ny	s->1	t->1	
ag nä	m->7	r->4	s->2	
ag nö	d->1	
ag oc	h->33	k->19	
ag of	t->1	
ag om	 ->27	b->1	
ag or	d->2	
ag os	v->1	
ag pe	r->5	
ag pl	ä->1	
ag po	l->1	s->2	ä->2	
ag pr	i->1	o->1	
ag på	 ->14	g->1	m->3	p->1	
ag re	d->13	f->1	g->1	k->4	s->1	
ag ri	k->2	s->1	
ag rä	d->1	k->5	
ag rå	d->2	
ag rö	r->3	s->10	
ag sa	d->10	k->1	m->1	
ag se	 ->1	d->3	r->11	t->1	
ag sj	ä->14	
ag sk	a->42	e->1	i->1	r->1	u->112	y->1	ä->1	
ag so	c->1	m->84	
ag sp	e->1	r->1	
ag st	o->1	ä->6	å->4	ö->10	
ag sv	a->2	
ag sy	f->4	m->2	
ag sä	g->32	k->3	r->2	
ag så	 ->1	g->2	l->1	
ag ta	 ->4	c->26	g->1	l->15	r->5	s->1	
ag ti	d->2	l->84	
ag to	g->2	
ag tr	o->115	
ag tv	i->2	u->1	å->1	
ag ty	c->42	d->3	v->1	
ag tä	n->16	v->1	
ag un	d->11	
ag up	p->38	
ag ut	 ->1	a->5	g->4	t->9	
ag va	d->2	l->1	r->9	
ag ve	r->8	t->23	
ag vi	d->5	l->262	s->3	
ag vä	d->2	g->1	l->16	n->7	x->1	
ag vå	g->2	
ag Ös	t->1	
ag äg	n->1	
ag äl	s->1	
ag än	d->4	n->1	
ag är	 ->110	,->2	l->1	
ag äv	e->2	
ag å 	e->1	u->1	
ag åt	 ->2	e->2	g->1	
ag ön	s->6	
ag öv	e->7	
ag, a	t->3	v->1	
ag, b	å->1	ö->1	
ag, d	e->3	v->1	ä->1	
ag, e	f->5	l->2	n->2	t->1	
ag, f	o->1	r->3	ö->7	
ag, g	e->2	
ag, h	a->1	e->3	
ag, i	 ->2	n->3	
ag, l	e->1	i->2	
ag, m	e->8	i->2	
ag, n	y->1	ä->2	
ag, o	a->1	c->9	
ag, p	å->1	
ag, s	o->10	p->1	ä->1	å->4	
ag, t	a->1	j->1	o->1	r->1	ä->1	
ag, u	t->5	
ag, v	a->2	i->4	o->1	
ag, ä	r->4	v->2	
ag. D	e->1	
ag. H	ä->1	
ag. P	å->1	
ag.(A	p->1	
ag.)F	ö->2	
ag.)H	e->1	
ag.. 	F->1	
ag.An	d->1	
ag.Ar	b->1	
ag.Av	 ->1	
ag.Be	k->1	t->1	
ag.De	n->8	s->1	t->10	
ag.Di	s->1	
ag.Dä	r->3	
ag.Ef	f->1	t->1	
ag.Er	i->1	
ag.Fr	a->1	u->1	å->1	
ag.Fö	r->5	
ag.Ge	n->1	
ag.He	r->6	
ag.Hu	r->1	
ag.Hy	c->1	
ag.I 	d->5	s->1	
ag.In	t->1	
ag.Ja	g->13	
ag.Ju	s->1	
ag.Ka	t->1	
ag.Ko	m->3	
ag.Li	v->1	
ag.Lå	t->1	
ag.Me	n->1	
ag.Må	n->2	
ag.Oc	h->1	
ag.Om	 ->1	
ag.Pa	r->1	
ag.Ra	p->1	
ag.Re	t->1	
ag.Sk	a->1	u->1	
ag.Sy	f->1	
ag.Ti	l->1	t->1	
ag.Un	g->1	
ag.Va	d->2	
ag.Vi	 ->5	s->1	
ag.Vå	r->1	
ag: d	e->1	
ag: j	a->1	
ag:De	n->1	
ag; s	l->1	
ag?De	n->1	
ag?Fi	n->1	
ag?Fr	u->1	
ag?Fö	r->1	
aga 2	 ->1	
aga H	a->1	
aga a	t->3	
aga d	e->5	i->2	
aga j	u->1	
aga n	å->1	
aga o	c->1	
aga r	e->2	
aga s	u->1	
aga!F	ö->1	
aga, 	k->1	o->1	
aga.D	e->1	
aga.F	ö->1	
aga.V	i->1	
agade	 ->5	
agan 	s->1	t->1	
agand	a->3	e->221	
agans	v->3	
agar 	a->4	d->6	e->4	f->2	h->2	i->1	j->2	o->3	p->1	s->5	t->3	v->2	ä->3	ö->1	
agar,	 ->5	
agar.	D->1	E->1	O->1	T->1	V->1	
agara	n->2	
agare	 ->40	"->1	,->10	.->7	n->10	s->3	
agarl	a->2	ä->1	
agarm	y->14	
agarn	a->25	
agars	 ->2	
agarv	ä->1	
agarä	m->1	
agas 	e->1	i->1	v->1	
agas,	 ->1	
agas.	P->1	
agask	a->1	
agast	e->2	
agat 	m->1	
agate	l->2	
agats	 ->2	
agav 	K->1	i->1	o->1	
agbar	 ->2	.->1	a->2	t->10	
agd a	t->1	
agd i	n->1	
agd o	c->1	
agd p	å->1	
agd, 	m->1	
agda 	f->1	h->2	o->1	r->1	ä->1	
agda.	V->1	
age p	r->1	
age s	o->1	
agedi	 ->1	.->1	e->2	
agel,	 ->1	
agels	e->5	
agema	n->9	
agen 	-->2	1->6	2->3	3->4	4->2	7->1	a->2	b->3	d->2	e->2	f->15	g->3	h->5	i->12	k->2	m->1	n->1	o->18	p->2	r->2	s->12	t->14	u->4	ä->7	å->1	
agen!	R->1	
agen,	 ->15	
agen.	(->1	B->1	D->4	F->1	H->1	J->6	K->2	M->1	N->1	S->2	V->2	
agen:	 ->2	
agen;	 ->1	
agend	a->1	
agens	 ->55	
agent	u->1	
ager 	t->2	
ager.	T->1	
agera	 ->31	,->3	.->1	d->5	n->12	r->12	t->5	
agerk	r->1	
ages-	 ->1	
aget 	(->2	-->1	A->1	R->1	a->10	b->4	e->5	f->14	g->6	h->4	i->10	k->6	l->4	m->1	n->1	o->19	p->4	r->2	s->17	t->18	u->1	v->1	ä->4	
aget)	 ->1	,->1	.->2	
aget,	 ->19	
aget.	A->1	D->6	E->1	F->4	H->2	I->2	J->5	K->1	L->1	M->3	N->1	O->2	P->1	S->2	T->1	V->1	
aget:	 ->1	
aget;	 ->1	
aget?	V->1	
agets	 ->18	
agett	,->1	
agför	s->5	
agg d	e->1	
agg f	a->1	
agg i	n->1	
agg m	a->1	
agg o	c->1	
agg s	o->1	
agg, 	e->2	i->1	k->1	m->1	t->1	v->1	
agg.D	ä->1	
agg.F	ö->1	
agg.K	o->1	
agg.M	a->1	
agg.N	u->1	
agg; 	f->1	
agga 	f->2	
aggad	e->2	
aggan	 ->1	
aggen	 ->1	s->1	
aggni	n->1	
aggor	n->1	
aggre	s->1	
agh m	e->1	
aghet	 ->4	.->1	e->7	
aginä	r->1	
agisk	a->5	t->1	
agit 	-->1	a->5	b->3	d->7	e->10	f->5	h->8	i->7	k->1	l->2	m->2	n->4	o->2	p->4	s->8	t->8	u->13	v->3	ä->1	å->1	
agit,	 ->2	
agit.	F->2	I->1	M->1	
agita	t->1	
agits	 ->22	,->2	.->3	
agiva	n->2	
agivi	t->1	
aglig	 ->2	.->1	a->10	e->8	h->2	t->12	
agmar	 ->1	
agmat	i->1	
agn f	ö->3	
agna 	d->2	e->1	g->1	i->3	k->1	l->1	m->2	o->1	p->3	r->1	s->1	u->1	v->1	ä->3	å->1	ö->1	
agna,	 ->1	
agna.	D->1	I->1	
agnad	e->4	
agnar	 ->2	
agnat	 ->2	i->1	
agne 	f->1	i->1	o->2	s->3	
agne-	A->1	
agnen	 ->2	
agner	a->1	
agnes	 ->1	
agnin	g->69	
agnis	k->1	
agnit	u->1	
agoge	r->1	
agogi	 ->1	.->2	s->1	
agolf	e->4	
agom 	a->1	
agomå	l->3	
agor 	t->2	
agor?	Ä->1	
agord	n->52	
agorn	a->2	
agosk	r->1	
agraf	 ->1	r->2	
agran	t->1	
agrar	 ->1	a->1	
agren	,->1	
agrot	u->1	
agrup	p->1	
ags a	n->1	t->8	
ags d	a->1	
ags f	a->1	r->1	y->1	ö->5	
ags i	d->1	n->1	
ags m	å->1	
ags o	m->3	
ags p	r->1	å->1	
ags r	a->1	e->1	
ags s	i->1	k->1	t->1	
ags u	n->1	t->1	
ags v	a->1	e->1	
ags, 	1->1	u->1	
ags.F	ö->1	
agsam	h->2	m->1	
agsan	a->1	
agsar	t->1	
agsav	t->1	
agsbe	s->1	
agsbo	r->1	
agsde	l->1	
agsek	o->5	
agsfa	l->1	
agsfä	s->1	
agsfö	r->3	
agsgi	v->8	
agsgr	u->2	
agsin	t->1	
agsju	r->2	
agsko	n->1	
agskr	a->1	
agsli	v->1	
agslä	g->2	
agsmä	s->2	
agsna	r->1	
agsne	d->1	
agsre	f->1	g->4	
agsrå	d->2	
agssi	t->1	
agsst	ö->3	
agsta	d->1	
agste	x->2	
agsti	d->2	f->127	l->2	
agsän	d->3	
agt -	 ->1	
agt 4	8->1	
agt a	l->2	t->12	v->1	
agt b	e->1	å->1	
agt d	e->2	
agt e	d->1	
agt f	l->1	r->27	ö->2	
agt i	 ->3	n->1	
agt j	a->1	
agt m	i->1	ä->1	ö->1	
agt n	e->9	å->1	
agt o	c->1	
agt s	i->2	
agt ä	r->1	
agt, 	h->1	k->1	o->1	s->1	u->1	v->2	ä->2	
agt. 	I->1	
agt.J	a->1	
agtex	t->2	
agts 	-->2	8->1	a->5	b->1	f->17	h->3	i->3	n->1	o->1	t->1	u->1	
agts,	 ->2	
ague,	 ->1	
agång	 ->3	,->1	s->6	
ahand	s->1	
ahus 	u->1	
ahåll	a->36	e->2	i->5	
ai La	m->7	
aider	 ->13	,->3	.->3	s->18	
aids 	i->1	ä->1	
aids-	s->1	
aidsp	a->2	
ail m	e->1	
aille	s->1	
ailur	e->1	
ain",	 ->1	
ain, 	h->1	
aine 	h->1	n->1	
aine,	 ->1	
ainsa	m->2	
ainst	a->22	r->8	
aint-	E->1	
aire.	D->1	
aiva 	o->1	
aivit	e->1	
aiwan	 ->1	
aj 19	9->3	
aj 20	0->1	
aj fö	r->1	
aj, o	c->1	
aj.Ja	g->1	
aj.To	n->1	
ajori	t->42	
ajour	n->1	
ak at	t->4	
ak be	r->1	s->1	
ak fö	r->1	
ak gä	l->3	
ak ha	r->3	
ak ho	p->1	
ak hä	n->1	
ak i 	k->1	
ak in	t->1	
ak ja	g->1	
ak ko	m->1	
ak ku	r->1	
ak lo	v->1	
ak me	d->2	r->1	
ak mo	t->1	
ak må	s->1	
ak nä	r->1	
ak sa	d->1	
ak se	g->1	
ak sj	ä->1	
ak so	m->9	
ak ti	l->3	
ak ut	 ->1	
ak va	d->1	r->1	
ak vi	 ->2	d->1	l->1	
ak är	 ->2	
ak öv	e->1	
ak, a	t->1	
ak, b	e->1	
ak, h	ä->1	
ak, m	e->1	
ak, s	o->1	
ak, v	ä->1	
ak.At	t->1	
ak.De	 ->2	t->1	
ak.Et	t->1	
ak.Ni	 ->1	
ak.Tr	ä->1	
ak.Ty	v->1	
ak: g	e->1	
ak?Ne	j->1	
aka -	 ->1	
aka E	u->1	
aka a	l->1	v->1	
aka b	e->2	i->1	
aka d	e->6	
aka e	n->2	t->1	
aka f	r->2	ö->1	
aka g	e->2	i->1	
aka i	 ->3	n->1	
aka j	ä->1	
aka k	l->1	
aka m	e->2	o->2	ä->1	
aka o	c->7	n->1	
aka p	r->1	u->1	
aka r	i->1	ä->1	
aka t	i->9	r->1	
aka v	e->1	
aka ö	v->1	
aka.D	e->1	
aka.I	 ->2	
aka.L	å->1	
aka.M	e->1	
aka?I	 ->1	
akade	 ->2	.->1	m->1	
akadr	a->3	
akagå	n->4	
akamm	a->1	
akar 	F->1	f->1	m->1	r->1	v->3	ö->1	
akare	,->1	
akas 	a->2	e->1	f->1	
akass	e->1	
akat 	9->1	f->1	k->1	s->1	u->1	
akat.	D->1	H->1	
akats	 ->2	
akavi	s->4	
akdör	r->1	
ake, 	s->1	
akel 	-->1	o->1	s->1	
aken 	b->1	m->1	t->4	u->1	
aken,	 ->2	
aken.	J->1	
aken:	 ->1	
aken?	J->1	
akens	 ->3	
aker 	f->1	h->2	i->2	j->2	m->1	n->1	o->5	s->10	t->1	
aker,	 ->3	
aker.	-->1	D->3	M->1	
aker:	 ->1	
akern	a->11	
aket 	f->1	g->1	i->1	k->1	m->1	o->1	
aket.	J->1	
akete	t->3	
akför	h->1	
akgru	n->31	
akien	 ->1	
akis 	f->1	i->1	p->1	
akis!	 ->1	
akisb	e->1	
akisk	a->1	
akist	a->5	
akkun	n->1	s->1	
aklas	s->1	
aklig	a->1	e->9	t->1	
akluk	t->1	
akna,	 ->1	
aknad	e->5	
aknar	 ->11	
aknas	 ->15	,->3	.->2	
aknat	 ->1	s->1	
aknin	g->14	
akolo	g->1	
akom 	-->1	d->10	e->1	f->1	l->1	m->2	o->2	p->1	r->2	
akom,	 ->1	
akoml	i->1	
akomr	å->2	
akonv	e->1	
akopo	u->5	
akpro	b->1	
akrer	a->1	
akroe	k->5	
akrof	i->1	
akry.	D->1	
akryg	g->1	
aks b	e->1	
aks d	e->1	
aks p	e->1	
aks s	a->1	
aksam	 ->3	h->2	m->4	
aksod	l->1	
aksta	n->1	
akt -	 ->1	
akt a	t->3	
akt b	l->1	
akt d	e->4	
akt e	f->1	
akt f	r->1	ö->6	
akt h	u->2	
akt i	 ->2	n->1	
akt l	ä->1	
akt m	e->8	o->1	
akt o	c->8	m->2	
akt p	å->5	
akt s	o->1	
akt u	t->2	
akt v	a->2	i->1	
akt ä	n->1	
akt, 	a->1	b->1	o->1	
akt.B	o->1	å->1	
akt.D	e->1	ä->1	
akt.J	a->2	
akt.M	a->2	
akt.V	a->1	
akt: 	d->1	
akta 	a->1	b->2	d->4	h->1	i->1	m->1	o->4	p->1	r->2	s->9	t->1	u->2	v->1	
akta.	F->1	
aktad	e->1	
aktai	n->2	
aktan	 ->4	d->5	s->1	
aktar	 ->12	.->1	e->6	n->5	
aktas	 ->15	.->1	
aktat	 ->4	s->4	
aktba	l->2	
aktbe	f->2	
aktde	l->1	
aktdi	k->1	
akten	 ->8	,->1	.->1	s->2	
akter	 ->11	.->2	i->3	n->4	
aktet	 ->1	
aktfa	r->1	
aktfö	r->1	
aktha	v->1	
akthe	t->1	
akthå	l->1	
aktie	b->1	ä->2	
aktig	 ->7	.->3	a->3	h->8	t->13	
aktik	 ->1	,->1	e->10	
aktio	n->17	
aktis	k->74	
aktiv	 ->5	.->1	a->4	e->1	i->9	t->17	
aktko	n->1	
aktli	g->14	
aktlö	s->3	
aktme	d->2	
aktmi	s->1	
aktor	 ->6	,->1	.->2	e->14	h->1	
aktta	 ->3	g->1	r->1	s->3	
aktua	l->1	
aktue	l->31	
aktum	 ->64	,->1	.->2	e->1	
aktär	 ->4	,->1	.->1	e->3	
aktör	 ->1	e->12	
akulä	r->1	
akuta	 ->1	
akuum	 ->1	t->1	
akämn	e->1	
akåt 	i->2	
akåts	t->1	
al - 	d->1	n->1	
al Co	u->1	
al De	n->1	
al In	t->2	
al Ka	n->1	
al Ul	s->1	
al ar	t->1	
al at	t->1	
al av	 ->25	
al be	r->1	s->1	t->2	v->1	
al bi	d->2	l->3	
al br	i->1	
al co	r->1	
al de	m->1	n->2	s->1	
al du	m->2	
al ef	f->2	
al el	l->1	
al en	d->1	
al fo	r->1	
al fr	a->1	å->8	
al få	r->1	
al fö	l->1	r->8	
al gö	r->1	
al ha	r->2	
al hä	r->1	
al i 	E->1	d->2	f->1	n->1	s->1	t->1	v->1	
al in	b->1	d->2	g->1	o->4	t->3	v->1	
al ka	n->2	
al ko	d->1	l->1	
al kv	i->2	
al lä	n->2	t->1	
al ma	r->1	
al me	d->9	l->7	
al mi	n->1	
al mo	t->1	
al mä	n->1	
al må	n->2	s->1	
al mö	j->1	
al ni	v->3	
al no	g->1	
al ny	a->1	
al oc	h->22	
al om	 ->10	v->1	
al or	d->1	
al pe	r->1	
al pl	a->3	
al po	l->1	s->1	
al pr	a->1	e->1	i->2	o->1	
al på	 ->2	
al ra	m->1	
al re	d->1	g->2	
al ri	k->1	
al ro	l->3	
al rä	t->2	
al sa	k->1	m->8	
al se	r->1	
al si	t->3	
al sj	ä->1	
al sk	a->2	u->1	
al so	c->1	l->1	m->24	
al st	a->4	ä->1	
al sv	a->1	å->1	
al sy	n->1	
al sä	k->2	
al ti	l->7	
al tr	y->3	
al ty	c->1	
al un	d->1	
al up	p->1	
al ut	a->2	s->7	v->2	
al va	r->2	
al ve	r->2	
al än	 ->1	
al är	 ->6	
al åk	l->1	
al ås	i->1	
al åt	 ->1	
al öv	e->3	
al!Hä	r->1	
al" m	e->1	
al" o	c->1	
al, T	y->1	
al, a	t->1	v->1	
al, d	e->1	i->1	
al, e	f->1	
al, g	r->1	
al, h	a->2	
al, l	a->1	
al, m	e->1	
al, n	å->1	
al, o	c->6	
al, r	e->1	
al, s	o->2	
al, t	i->1	
al, v	i->2	
al- o	c->7	
al-Fi	n->3	
al-Sh	a->1	
al-so	c->2	
al. J	a->1	
al.De	s->1	t->4	
al.En	l->1	
al.Fr	u->1	
al.Fö	r->4	
al.He	r->2	
al.Hu	r->1	
al.I 	u->1	
al.In	g->1	
al.Ja	 ->1	g->1	
al.Ka	n->1	
al.Ko	m->1	
al.Me	n->1	
al.Pe	r->1	
al.Sa	m->1	
al.Sj	ä->1	
al.St	r->1	
al.Så	 ->1	
al.Vi	 ->3	
al: O	s->1	
al: p	r->1	
al; a	t->1	
alFin	a->1	
ala E	u->1	
ala K	o->1	
ala a	k->2	l->2	s->2	v->2	
ala b	a->1	e->6	i->1	u->1	
ala d	e->4	i->5	ö->1	
ala e	k->5	l->3	n->5	r->1	t->2	u->1	x->1	
ala f	a->1	o->2	r->4	u->1	ö->5	
ala g	i->2	r->5	
ala h	a->1	i->1	o->1	
ala i	 ->1	d->3	n->6	
ala j	ä->1	
ala k	a->1	l->2	o->6	
ala l	e->3	i->2	ö->1	
ala m	a->3	e->4	i->9	o->2	y->15	ä->1	ö->2	
ala n	o->1	
ala o	b->3	c->29	j->1	l->1	m->44	p->2	r->3	s->1	
ala p	a->9	e->1	o->2	r->10	
ala r	e->2	u->1	ä->2	ö->2	
ala s	a->12	e->1	i->16	j->1	k->12	t->5	u->1	y->1	å->1	
ala t	i->2	j->1	r->1	
ala u	n->1	p->2	r->1	t->15	
ala v	e->1	i->2	ä->3	å->1	
ala ä	n->1	r->1	
ala å	 ->1	t->2	
ala ö	v->1	
ala";	 ->1	
ala, 	d->1	l->1	n->1	o->1	ä->1	
ala.D	e->4	
ala.I	 ->1	
ala.J	a->1	
ala.K	o->1	
ala.S	m->1	
ala?D	e->3	
alaci	o->15	
alad 	i->1	
alade	 ->33	s->1	
alafr	a->1	
alag 	n->1	o->1	s->1	
alag,	 ->1	
alage	n->1	
alai 	L->7	
alam,	 ->1	
alan 	f->1	v->1	
alan.	 ->1	J->1	
aland	e->52	
alang	e->1	
alank	l->1	
alans	 ->14	,->2	e->16	l->1	v->1	ö->1	
alar 	2->1	a->2	e->1	f->8	g->1	i->2	j->2	m->7	n->2	o->28	p->1	r->1	s->8	t->1	v->3	ä->1	
alar,	 ->2	
alar.	D->1	E->1	F->1	J->1	
alar?	K->1	
alare	 ->18	,->4	.->1	n->7	
alarn	a->13	
alars	t->1	
alart	i->2	
alas 	d->1	e->1	o->4	p->1	s->1	t->1	u->1	
alas,	 ->1	
alasi	a->2	e->4	
alat 	a->1	e->1	f->2	g->1	i->1	m->1	n->1	o->9	s->1	u->1	ö->1	
alat,	 ->3	
alat.	I->1	V->1	
alate	r->1	
alatl	a->1	
alats	 ->5	.->1	
alaya	b->1	
alban	 ->1	e->5	k->8	s->4	
albar	h->1	
albel	o->1	
albes	t->2	
alblo	c->1	
ald f	r->4	
ald i	 ->1	n->1	
ald k	o->1	
ald p	o->1	u->1	
ald r	e->1	
ald ä	r->1	
ald, 	d->1	k->1	m->2	o->2	
ald.J	a->1	
alda 	f->3	i->2	o->1	p->3	r->3	s->1	
alda,	 ->1	
alda?	F->1	
aldag	e->1	
alde 	e->2	
aldel	t->3	
aldem	o->16	
alden	 ->4	.->1	
aldes	 ->3	
aldez	,->1	-->2	
aldig	a->1	t->1	
aldir	e->17	
aldis	t->1	
aldju	r->1	
aldom	s->1	
aldri	g->31	
aleid	o->2	
alejd	o->1	
aleko	n->4	
alem 	h->1	o->1	
alen 	B->1	b->1	f->2	h->1	i->7	m->3	o->2	s->2	t->2	
alen,	 ->3	
alen.	M->2	V->1	
alen?	Ä->1	
alens	k->1	
alent	i->1	
aleot	e->1	
aler 	b->1	m->2	o->3	p->1	s->3	t->1	
aler,	 ->1	
aler.	D->1	J->1	M->1	
alerm	o->1	
alern	a->5	
ales 	e->2	f->1	h->1	p->1	s->2	u->1	
ales.	H->1	V->1	
ales;	 ->1	
alesa	r->1	
alese	 ->1	
alesm	a->1	ä->1	
alest	i->22	
alesä	t->2	
alet 	E->1	T->1	a->4	b->1	d->1	e->4	f->5	g->1	h->2	i->2	k->1	l->2	m->7	n->1	o->5	p->1	r->2	s->5	t->2	u->1	v->2	ä->1	å->1	
alet,	 ->11	
alet.	D->3	H->1	I->1	
alets	 ->3	
aleur	o->1	
alfab	e->1	
alfon	d->15	
alfor	d->3	
alfra	m->3	
alfri	h->2	
alfrå	g->5	
alfån	g->4	
alför	b->1	s->9	v->1	
alibe	r->1	
alibi	 ->1	
alici	e->2	
alien	 ->12	,->5	.->1	s->18	
alier	 ->4	
alies	t->1	
alifi	c->14	k->1	
alig 	e->1	o->1	
aliga	,->2	
aligt	 ->1	
alina	r->1	
alini	s->2	
alinr	i->1	
alise	r->64	
alisk	 ->1	a->4	
alism	 ->6	.->1	?->1	e->3	
alist	e->24	g->3	i->33	k->1	p->5	
alita	r->2	t->6	
alite	t->50	
aliti	o->14	
alj o	m->1	
alj ö	v->1	
alj, 	o->1	ä->1	
alj.V	i->1	
aljan	a->1	
aljer	 ->3	,->2	.->1	a->16	n->4	
aljfl	ö->1	
aljko	n->2	
alkan	 ->3	.->4	
alkem	i->1	
alkoh	o->1	
alkor	,->1	
alkre	t->4	
all 7	5->1	
all E	G->1	u->1	
all K	o->1	
all a	c->1	g->1	l->3	n->16	r->4	t->1	v->11	
all b	a->5	e->40	i->4	l->22	o->1	r->1	ä->3	ö->2	
all c	e->1	i->2	
all d	e->21	i->5	r->1	ä->4	å->3	
all e	f->1	k->1	n->3	r->2	t->1	x->1	
all f	a->5	e->1	i->4	o->4	r->8	u->8	y->2	å->9	ö->26	
all g	a->3	e->12	o->3	r->2	ä->7	å->7	ö->18	
all h	a->34	e->1	i->3	j->3	o->1	å->2	ö->2	
all i	 ->1	n->49	
all j	a->11	u->3	
all k	a->3	l->1	o->20	r->3	u->55	
all l	e->2	i->5	y->6	ä->8	å->1	ö->1	
all m	a->7	e->3	i->1	o->1	u->1	y->1	å->2	ö->2	
all n	a->2	i->1	u->2	ä->1	å->1	
all o	c->6	f->1	m->11	r->1	ä->2	
all p	a->2	e->3	o->1	r->4	u->1	å->1	
all r	a->1	e->3	i->1	y->1	ä->5	ö->1	
all s	a->4	e->10	i->2	k->15	l->2	o->11	p->2	t->14	ä->5	ö->1	
all t	a->19	i->8	o->1	r->6	v->1	y->1	ä->2	
all u	n->8	p->10	t->14	
all v	a->31	e->5	i->26	ä->1	å->1	
all ä	g->1	n->3	r->4	v->3	
all å	s->2	t->8	
all ö	k->3	v->8	
all",	 ->1	
all, 	d->1	h->1	i->1	j->1	m->2	o->1	s->2	v->2	å->1	
all. 	D->1	o->1	
all.B	i->1	
all.D	e->4	
all.E	n->1	
all.H	e->1	
all.J	a->3	
all.M	e->1	
all.S	a->1	
all.V	i->2	
alla 	-->1	E->3	H->1	a->29	b->10	d->60	e->16	f->30	g->5	h->12	i->10	j->1	k->18	l->10	m->29	n->8	o->15	p->16	r->12	s->34	t->10	u->2	v->17	ä->3	å->1	ö->4	
alla!	H->1	
alla,	 ->5	
alla.	D->3	J->1	
allad	 ->5	e->5	
allan	d->6	
allar	 ->7	
allas	 ->6	
allat	 ->5	
allde	l->23	
alleg	o->1	
alleh	a->3	
allel	e->3	l->5	s->2	
allen	 ->6	,->1	.->1	a->1	
aller	 ->41	,->1	.->2	a->1	
alles	a->5	
allet	 ->36	!->1	,->9	.->10	
alleu	r->2	
allfä	r->1	
allia	n->7	
allib	e->1	
allie	r->1	
allih	o->1	
allin	d->1	
allit	 ->4	
allkl	a->2	
allmo	s->1	
allmä	n->121	
allmö	s->1	
allok	e->1	
allpo	l->1	
allra	 ->9	
allri	n->1	
alls 	a->1	b->1	d->1	h->1	i->2	n->1	p->1	s->4	ä->1	ö->1	
alls,	 ->1	
alls.	F->1	T->1	
allsf	ö->1	
allsh	a->1	
allsi	d->1	
allsm	ä->1	
allss	t->3	
allst	r->4	u->1	
allsä	m->1	
allt 	-->1	a->10	b->5	d->25	e->3	f->19	g->4	h->1	i->17	k->14	m->7	n->5	o->5	p->8	r->2	s->21	t->2	u->6	v->11	ä->6	ö->1	
allt,	 ->7	
allt.	D->3	M->2	V->1	
allt:	 ->1	
alltf	l->1	ö->38	
allti	d->77	h->1	n->5	
alltj	ä->3	
alltm	e->1	
allts	a->1	e->1	å->61	
allva	r->74	
ally 	f->1	
ally!	 ->1	
ally.	A->1	
allyb	e->1	
allys	 ->1	
alman	 ->7	!->242	,->157	:->1	n->11	s->9	
almed	e->1	
alna 	k->1	
alnin	g->15	
alog 	a->1	m->9	o->1	s->5	ä->1	
alog,	 ->1	
alog.	D->1	F->2	H->1	J->2	N->1	
aloge	n->8	
alpar	l->1	
alpat	r->1	
alpol	i->44	
alpro	d->1	g->1	
alres	u->4	
alrik	a->4	
alräk	e->1	
als a	r->2	
als b	a->1	
als f	a->2	i->1	r->1	
als g	a->1	
als h	e->1	
als i	l->1	n->1	
als k	v->1	
als m	i->3	ä->2	
als o	c->2	r->2	
als p	r->2	
als s	e->1	o->1	
als å	r->2	
als.D	e->1	
alsek	r->2	
alsfa	s->1	
alska	 ->1	.->1	t->3	
alskn	i->1	
alsko	m->1	
alskt	 ->1	
alsku	l->1	
alslö	s->1	
alsoc	i->1	
alspa	r->1	
alspu	n->6	
alsru	n->1	
alsst	i->1	
alsta	t->3	
alstö	d->2	
alsum	m->1	
alsys	t->1	
alt 2	7->1	
alt 7	0->1	
alt 9	5->1	
alt E	U->1	
alt a	n->3	t->4	v->1	
alt b	e->1	
alt d	e->1	
alt f	i->1	ö->1	
alt h	a->5	
alt i	 ->7	n->2	
alt m	i->1	
alt n	o->1	
alt o	c->3	m->1	
alt p	l->3	r->1	
alt r	i->1	ä->2	
alt s	a->1	e->3	t->3	ä->2	
alt t	i->2	
alt u	p->2	t->1	
alt v	i->2	
alt ä	n->1	v->1	
alt, 	f->1	m->2	o->1	å->1	
alt.D	e->2	
alt.J	a->1	
alt.O	m->1	
alt.V	a->1	i->1	
alta 	i->1	o->2	s->1	u->1	ä->1	
alta,	 ->1	
altak	t->1	
altar	 ->1	e->1	
altas	 ->1	
alter	 ->1	n->12	
altes	i->3	
altid	e->1	
altni	n->47	
alts 	o->1	p->1	s->1	u->1	
alts.	K->1	
alufö	r->1	
alund	a->3	
aluta	 ->1	,->1	f->10	n->5	p->1	s->2	u->3	
alutb	i->2	
alv d	a->1	
alv m	e->1	
alv t	i->2	
alva 	t->2	v->2	
alver	s->1	
alvhj	ä->1	
alvin	i->1	
alvmi	l->1	
alvof	f->1	
alvol	y->1	
alvt 	å->2	
alvti	d->1	m->2	
alvvä	g->2	
alvår	 ->1	e->2	s->2	
alvö,	 ->1	
alvö.	D->1	
alvön	 ->1	
alyda	n->1	
alyde	l->2	
alys 	-->1	a->16	f->2	g->1	i->1	j->1	o->2	s->1	v->1	
alys,	 ->4	
alys.	D->2	F->1	G->1	H->1	
alys?	D->1	I->1	
alysa	t->2	
alyse	n->5	r->16	
alösa	 ->1	
am "K	u->1	
am - 	K->1	e->1	i->1	o->1	s->1	
am 19	9->1	
am 80	 ->1	
am De	t->1	
am ac	c->1	
am al	t->1	
am ar	m->1	
am as	y->2	
am av	 ->4	,->1	
am be	h->1	l->1	s->1	t->2	
am bl	i->1	
am bu	d->1	
am co	r->1	
am da	g->1	
am de	 ->5	b->1	f->1	n->3	t->11	
am di	p->1	s->1	
am ef	t->1	
am em	o->17	
am en	 ->13	b->1	o->1	
am er	f->1	
am et	t->23	
am eu	r->2	
am fl	e->1	
am fo	r->1	
am fr	a->1	
am fö	l->1	r->44	
am ge	r->1	
am gr	u->1	
am gö	r->2	
am ha	r->4	
am he	t->1	
am hä	n->1	r->3	
am hå	l->1	
am i 	C->1	T->1	d->2	e->1	f->1	k->1	p->1	r->1	s->1	t->2	ö->1	
am in	f->2	i->1	r->2	
am ka	n->1	
am ko	n->2	
am kv	a->1	
am la	g->2	
am li	k->1	
am lä	g->1	
am lö	s->2	
am ma	r->2	
am me	d->5	l->1	n->2	r->2	
am mi	l->1	
am mo	t->1	
am my	c->1	
am må	s->4	
am ni	 ->1	
am no	r->1	
am nu	 ->1	
am nä	r->2	
am nå	g->2	
am oc	h->8	k->1	
am om	 ->5	f->1	
am po	l->1	
am pr	o->1	
am på	 ->10	
am ra	m->1	
am re	d->1	g->2	k->1	s->4	
am ri	k->1	
am rä	t->1	
am sa	d->1	k->2	m->1	
am si	t->3	
am sk	a->3	u->1	
am sl	u->1	
am so	m->12	
am sp	e->1	
am st	a->1	r->1	å->5	
am sy	f->1	s->1	
am sä	k->3	
am så	 ->2	
am ta	n->1	
am ti	d->1	l->46	
am tr	a->1	e->2	
am un	d->1	
am ut	i->1	r->1	t->1	
am va	l->1	r->3	
am ve	r->2	
am vi	 ->1	d->2	
am vå	r->2	
am än	d->2	
am är	 ->2	
am äv	e->1	
am åk	l->1	
am ås	i->1	
am åt	g->1	
am ök	n->1	
am öv	e->3	
am!De	n->1	
am, K	u->1	
am, a	l->1	t->1	
am, b	l->1	ö->1	
am, d	e->3	
am, e	t->1	
am, f	i->1	r->1	
am, i	 ->1	
am, j	u->1	
am, m	e->2	
am, n	ä->1	
am, o	c->7	
am, p	r->1	
am, r	e->1	
am, s	o->2	ä->1	å->4	
am, u	t->2	
am, v	e->1	i->1	
am..(	F->1	
am.De	n->2	t->3	
am.Fr	u->3	
am.Fö	r->1	
am.Ge	n->1	
am.Gö	r->1	
am.He	r->1	
am.Hu	r->1	
am.I 	d->1	
am.Ja	g->2	
am.Ko	s->1	
am.Ku	l->1	
am.Me	n->2	
am.Na	t->1	
am.Nä	r->1	
am.Om	 ->1	
am.Re	f->1	
am.Sl	u->1	
am.St	a->1	
am.Sy	f->1	
am.Ti	l->1	
am.Vi	 ->2	
am?Ja	g->1	
am?Vi	l->1	
ama -	 ->1	
ama h	a->1	
ama o	c->1	
ama p	å->1	
ama s	ä->1	
ama u	p->1	
ama.J	a->1	
ama.V	i->1	
amaff	ä->1	
amans	v->1	
amar 	f->1	s->1	
amar,	 ->3	
amar.	J->1	
amarb	e->83	
amarn	a->2	
amas 	f->1	s->1	
amask	u->1	
amati	s->6	
amavt	a->3	
ambal	a->1	
amban	d->47	
ambas	s->1	
ambit	i->26	
ambul	a->1	
ambur	g->2	
ame-f	a->1	
amels	 ->1	
amen 	f->54	k->1	o->4	v->1	
amen,	 ->4	
amens	b->2	
ament	 ->58	,->10	.->9	a->24	e->473	s->35	
amer 	o->41	
amera	 ->1	n->1	
ameri	k->15	
amete	r->1	
ametr	a->1	
amexi	s->2	
amfar	t->1	
amfin	a->1	
amfun	d->5	
amför	 ->97	a->23	d->36	h->1	k->1	s->9	t->12	
amgic	k->1	
amgå 	i->1	
amgån	g->38	
amgår	 ->12	
amgåt	t->1	
amhet	 ->56	,->5	.->7	?->1	e->21	s->7	
amhäl	l->49	
amhär	d->1	
amhäv	a->3	e->1	
amhål	l->17	
amhöl	l->2	
amidi	s->1	
amik 	e->1	
amilj	 ->1	e->14	
amina	t->2	
amine	r->10	
aming	 ->4	"->1	)->3	
amini	s->1	
amisk	 ->2	a->2	
amkar	 ->1	
amkas	t->1	
amkat	 ->1	,->1	
amkom	m->10	
amla 	U->1	b->7	d->1	f->6	h->1	i->5	k->5	l->1	m->2	o->1	r->1	s->5	t->1	u->1	
amlad	e->2	
amlag	d->3	t->9	
amlar	 ->2	f->1	
amlas	 ->1	
amlat	 ->3	s->2	
amlev	n->1	
amlig	.->1	a->1	
amlin	g->25	
amläg	g->8	
amm a	v->1	
amma 	1->1	E->1	a->7	b->7	d->8	e->4	f->10	g->3	h->4	i->12	j->5	k->13	l->4	m->12	n->6	o->7	p->12	r->14	s->96	t->2	u->13	v->9	å->3	ö->2	
amma,	 ->4	
amma.	H->1	J->1	
ammad	e->1	
ammal	 ->4	
amman	 ->18	,->1	.->1	b->6	d->1	f->15	h->101	j->1	k->12	l->2	s->57	t->35	
ammar	 ->2	,->1	e->63	n->2	
ammas	 ->2	
ammat	 ->3	s->1	
amme 	k->1	s->1	
ammen	 ->24	,->4	.->8	
ammer	f->22	
ammet	 ->53	)->2	,->6	.->9	:->1	s->2	
amn K	o->1	
amn b	y->1	
amn i	 ->1	
amn k	a->1	
amn m	e->1	å->2	
amn o	c->1	
amn p	å->1	
amn s	o->1	v->1	
amn, 	m->1	u->1	
amn.D	e->1	
amn.M	e->1	
amn.V	i->1	
amna 	h->1	i->1	p->1	
amnad	e->1	
amnar	 ->14	.->2	n->6	
amnav	g->2	
amnbe	s->1	
amnen	 ->1	.->1	
amnet	 ->2	
amnin	g->2	s->1	
amnko	n->2	
amnup	p->4	
amo, 	d->1	
amod 	m->1	ä->1	
amord	n->38	
amot 	J->2	L->1	R->2	W->1	a->8	f->3	h->2	i->3	k->1	s->2	
amot!	 ->7	
amot,	 ->16	
amote	n->26	
amp J	ö->1	
amp f	ö->2	
amp i	 ->3	
amp m	e->1	o->4	
ampag	n->1	
ampan	j->6	
ampen	 ->14	,->1	.->1	
amper	i->3	
ampla	n->8	
ampor	,->1	
ampro	g->12	
ampål	e->1	
amrat	 ->1	
amre 	h->1	
amres	t->1	
amrun	d->1	
amrät	t->1	
amråd	 ->3	,->1	.->1	a->2	e->1	s->1	
ams B	l->1	
amskj	u->1	
amskr	i->1	
amsky	d->4	
amste	g->32	
amstä	l->10	m->4	
amstå	 ->1	e->3	r->1	
amstö	t->1	
amsyn	 ->2	,->1	
amt G	a->1	
amt H	e->1	
amt a	n->1	s->1	t->7	v->3	
amt b	e->3	ö->1	
amt d	e->2	
amt e	k->2	n->1	t->2	u->2	
amt f	o->1	r->2	ö->9	
amt h	a->1	
amt i	 ->2	n->1	
amt j	ä->1	
amt k	o->3	u->1	v->1	
amt l	u->1	ä->2	
amt m	e->1	i->1	o->1	å->2	
amt n	e->1	
amt o	c->4	m->5	
amt p	a->1	å->1	
amt r	e->3	y->1	ä->2	
amt s	i->1	k->1	t->4	y->1	
amt t	a->1	i->3	
amt u	n->1	p->2	t->5	
amt v	a->1	
amt y	t->1	
amt ä	n->1	v->2	
amt å	t->1	
amt ö	v->1	
amt, 	ä->2	
amt.P	å->1	
amt.U	n->1	
amt.Å	r->1	
amtag	a->3	i->1	n->1	
amtal	 ->4	a->1	e->9	s->2	
amtid	 ->7	,->3	.->6	:->1	a->22	e->64	i->67	s->4	
amtli	g->25	
amträ	d->2	
amtvi	n->2	
amtyc	k->6	
amus 	e->1	
amutf	o->1	
amver	k->4	
amvet	e->1	s->1	
amvil	l->3	
amål 	f->1	
amål,	 ->2	
amål.	I->1	M->1	
amåle	t->6	
amåls	e->2	
amåt 	i->5	m->3	o->2	p->1	v->1	
amåt,	 ->3	
amåt.	D->3	F->1	H->1	J->1	V->1	
amöte	r->84	
amöve	r->2	
an "e	n->1	
an - 	'->1	m->1	n->1	ä->2	ö->1	
an 10	0->2	
an 15	0->1	
an 17	 ->1	
an 19	6->3	7->1	8->3	9->15	
an 4 	e->1	
an 8 	o->2	
an Al	t->1	
an Am	o->1	
an Br	o->2	
an CE	N->1	
an Ce	n->1	
an Da	m->2	n->1	
an De	 ->1	
an EG	-->1	
an EK	S->1	
an EM	U->1	
an EU	,->1	
an Er	i->1	
an Eu	r->13	
an Fl	o->1	
an Fo	n->1	
an Ga	z->1	
an Go	r->1	
an Ha	i->1	r->1	
an Hu	l->23	
an Im	b->2	
an Is	a->1	r->10	
an Ju	n->1	
an Ko	c->2	
an La	n->1	
an Ni	e->1	
an Pa	l->1	
an Pl	a->1	
an Po	r->2	
an Pr	o->1	
an Ro	v->1	
an SP	Ö->1	
an Sc	h->1	
an Se	b->1	
an Sh	a->1	
an Sy	r->2	
an Ve	l->1	
an Wi	e->3	
an a 	p->1	
an ab	s->1	
an ac	c->10	
an ag	e->2	
an ak	t->1	
an al	d->2	l->10	
an am	b->1	
an an	a->2	d->6	g->2	l->1	n->1	s->12	t->5	v->12	
an ap	p->1	
an ar	b->7	k->1	
an at	t->102	
an av	 ->24	d->1	g->2	s->5	v->1	
an ba	d->1	n->1	r->11	
an be	a->5	d->2	f->4	g->3	h->5	k->4	n->1	r->4	s->8	t->10	v->4	
an bi	d->8	l->2	
an bl	a->2	e->3	i->7	
an bo	r->4	s->1	t->1	
an br	o->2	
an by	g->1	t->1	
an bä	r->1	t->1	
an bö	r->20	
an ce	n->2	
an ch	a->1	
an da	g->3	
an de	 ->32	b->6	c->3	f->1	l->4	m->2	n->27	r->8	s->17	t->40	
an di	r->2	s->4	
an do	c->2	m->1	
an dr	a->5	i->1	u->1	ö->2	
an dy	k->1	
an dä	r->13	
an då	 ->9	
an dö	l->1	p->2	
an ef	f->2	t->5	
an ek	o->3	
an el	e->1	l->3	
an em	e->6	i->1	
an en	 ->31	a->2	b->2	d->3	g->1	h->1	l->2	v->1	
an er	 ->1	b->1	h->1	k->3	s->3	t->1	
an et	t->10	
an ex	 ->1	e->1	i->2	
an fa	k->1	l->1	n->1	s->5	t->5	
an fe	m->1	
an fi	c->1	n->14	
an fl	e->4	o->1	
an fo	r->12	
an fr	a->7	e->1	o->1	ä->2	å->20	
an fu	l->2	n->2	
an fy	l->1	r->2	
an fä	s->2	
an få	 ->15	,->1	r->3	s->1	
an fö	d->1	l->1	r->100	
an ga	m->1	n->1	r->8	
an ge	 ->14	m->1	n->10	r->1	t->2	
an gi	v->1	
an gj	o->3	
an gl	ä->1	
an go	d->10	
an gr	a->2	i->1	u->1	
an gä	l->5	
an gå	 ->7	r->4	t->1	
an gö	r->36	
an ha	 ->5	d->7	f->2	n->3	r->98	
an he	j->1	l->6	
an hi	n->2	t->5	
an hj	ä->5	
an ho	p->3	s->1	
an hu	r->4	v->1	
an hä	l->1	n->9	r->9	v->2	
an hå	l->1	
an hö	g->2	r->1	
an i 	B->2	E->4	I->1	K->1	L->1	P->1	V->1	a->3	b->4	d->18	e->1	f->8	g->2	j->2	k->1	l->3	m->7	p->4	r->1	s->10	u->2	v->4	ä->1	å->1	
an ib	l->1	
an id	e->3	
an if	r->2	
an ig	n->1	
an in	b->2	d->1	f->10	g->1	h->1	k->2	l->4	n->5	o->5	r->1	s->6	t->114	v->1	
an is	r->1	t->1	
an it	a->1	
an ja	g->41	n->1	
an ju	 ->3	l->1	r->1	s->2	
an jä	m->2	
an ka	b->1	l->3	n->38	p->1	t->2	
an kl	a->2	i->1	
an kn	a->1	
an ko	m->56	n->10	r->1	s->3	
an kr	i->1	ä->6	ö->1	
an ku	l->1	n->5	
an kv	a->1	i->4	o->2	
an ky	l->1	
an kä	n->1	
an kö	n->3	r->1	
an la	d->1	g->5	
an le	d->10	v->2	
an li	d->1	g->1	k->2	t->1	
an lo	k->3	v->1	
an ly	c->5	s->2	
an lä	g->9	m->2	n->3	r->1	s->5	t->2	
an lå	n->1	t->1	
an lö	s->5	
an ma	j->1	k->1	n->32	
an me	d->42	l->5	r->1	
an mi	n->3	s->1	
an mo	t->6	
an my	c->3	n->4	
an mä	n->1	t->1	
an må	s->42	
an mö	j->2	t->1	
an na	t->10	
an ni	 ->8	v->1	
an no	m->1	t->2	
an nu	 ->14	
an ny	 ->1	s->2	
an nä	m->8	r->2	s->1	
an nå	 ->3	g->11	
an nö	d->1	
an oc	h->54	k->53	
an of	f->1	t->1	
an ol	i->3	
an om	 ->114	"->1	,->1	e->1	p->2	r->1	s->2	ö->3	
an op	e->1	p->1	
an or	d->2	o->2	s->3	
an os	s->1	
an ov	i->2	
an pa	r->6	
an pe	l->2	
an pl	a->2	ö->1	
an po	l->3	o->1	ä->2	
an pr	a->1	e->5	i->1	o->1	
an pu	n->1	
an på	 ->42	b->1	m->1	p->3	s->3	t->1	v->2	
an ra	d->1	m->1	p->1	
an re	d->8	f->1	g->15	k->2	p->1	s->8	v->1	
an ri	g->1	k->5	s->3	
an ro	s->1	
an ru	s->1	
an rä	d->1	k->2	t->2	
an rå	d->5	
an rö	r->3	s->4	
an sa	d->10	g->9	k->4	m->6	n->1	t->2	
an se	 ->7	d->4	r->6	
an si	g->6	t->7	
an sj	ä->1	
an sk	a->54	e->2	j->1	r->1	u->17	ä->1	ö->1	
an sl	u->5	å->1	
an sn	a->9	
an so	m->20	
an sp	a->1	e->4	l->1	
an st	a->4	i->1	o->2	r->5	y->1	ä->9	å->4	ö->7	
an sv	a->2	å->1	
an sy	n->1	r->2	
an sä	g->16	k->1	r->5	t->1	
an så	 ->5	l->1	
an ta	 ->12	c->2	g->6	l->19	p->1	r->3	s->5	
an te	c->1	k->1	n->1	
an ti	b->1	d->4	l->42	t->3	
an tj	ä->2	
an to	g->1	
an tr	a->1	e->1	o->1	ä->2	
an tv	e->13	i->17	ä->3	å->2	
an ty	c->2	d->1	n->1	v->1	
an tä	n->5	
an un	d->17	i->4	
an up	p->31	
an ur	 ->1	m->1	s->1	
an ut	,->1	a->2	b->2	e->1	f->6	g->2	l->1	n->4	r->2	s->2	t->6	v->6	ö->3	
an va	d->1	l->1	n->2	r->38	
an ve	k->1	r->11	t->7	
an vi	 ->55	d->20	k->5	l->13	n->1	s->8	
an vo	r->1	
an vr	i->1	
an vä	c->1	g->4	l->1	n->5	
an vå	r->1	
an yt	t->2	
an Ös	t->1	
an äg	a->2	e->1	n->3	t->1	
an än	 ->3	d->3	n->1	
an är	 ->71	,->1	:->2	
an äv	e->15	
an å 	e->2	
an år	 ->2	l->1	
an ås	i->1	t->4	
an åt	e->8	f->1	g->1	m->3	
an ök	a->1	
an ön	s->1	
an öp	p->2	
an öv	e->19	
an! A	l->2	t->1	v->2	
an! B	e->2	
an! D	a->1	e->30	ä->1	í->1	
an! E	U->1	n->1	u->3	
an! F	r->3	å->1	ö->8	
an! G	r->2	
an! H	e->1	
an! I	 ->9	n->1	
an! J	a->74	
an! K	o->5	
an! L	i->1	å->5	
an! M	a->1	i->4	
an! N	u->1	ä->4	
an! O	l->1	m->1	
an! P	a->1	r->1	å->2	
an! R	e->1	o->1	å->2	
an! S	c->1	e->3	k->1	o->3	t->1	
an! T	a->1	h->1	i->4	o->1	r->1	
an! U	n->2	t->2	
an! V	a->3	i->12	å->2	
an! Ä	n->1	v->6	
an! Å	 ->3	
an! Ö	s->1	
an!Am	s->1	
an!De	t->2	
an!Ef	t->1	
an!En	 ->1	
an!Ja	g->6	
an!Mi	n->1	
an!Sa	n->1	
an!Ta	c->1	
an!Ti	l->1	
an!Un	d->1	
an!Vi	 ->2	
an" a	t->1	
an" g	e->1	
an", 	s->1	
an".R	å->1	
an, K	a->1	o->1	
an, U	z->1	
an, a	n->5	t->7	
an, b	ä->2	
an, d	e->9	ö->1	
an, e	f->4	l->1	n->3	t->1	
an, f	a->1	r->16	å->1	ö->8	
an, g	a->1	e->1	j->1	
an, h	e->42	
an, i	 ->4	n->2	
an, j	a->4	
an, k	a->1	o->9	r->2	ä->22	
an, m	e->5	i->15	
an, n	ä->7	
an, o	c->10	m->2	
an, p	a->1	r->1	å->3	
an, r	å->1	
an, s	a->3	k->3	o->9	å->2	
an, t	a->1	i->2	r->1	
an, u	n->1	p->1	t->5	
an, v	a->2	e->1	i->5	ä->1	
an, ä	n->1	r->12	v->1	
an- o	c->1	
an-Cl	a->1	
an-Ke	e->1	
an. D	e->1	
an.(L	i->1	
an.(P	a->2	
an.) 	T->1	
an.Al	l->1	
an.Av	s->1	
an.De	 ->2	n->1	t->13	
an.Dä	r->2	
an.Då	 ->1	
an.Ef	t->1	
an.En	l->1	
an.Fr	u->1	
an.Fö	r->4	
an.He	r->3	
an.Hu	r->2	
an.I 	a->1	d->1	
an.Il	l->1	
an.In	t->1	
an.Ja	g->14	
an.Ko	m->3	
an.Lå	t->1	
an.Me	n->3	
an.Ni	 ->1	
an.Nä	r->1	
an.Oc	h->1	
an.Se	d->1	
an.Sk	u->1	
an.Sl	u->2	
an.So	m->1	
an.Så	 ->2	l->1	
an.Ta	c->1	
an.Ty	 ->1	
an.Un	d->2	
an.Ut	s->1	
an.Va	d->2	n->1	
an.Vi	 ->1	d->1	l->2	
an.Vå	r->2	
an: A	t->1	
an: K	o->1	
an: V	a->1	i->1	
an: n	ä->2	
an: v	i->1	
an; J	a->1	
an; d	e->1	
an; s	k->1	
an? 2	1->1	
an?Fr	u->1	
an?He	r->1	
an?Hu	r->1	
an?Ja	g->1	
an?Om	 ->1	
an?Se	d->1	
an?Ve	t->1	
an?Är	 ->1	
anNäs	t->1	
ana -	 ->2	
ana E	l->1	
ana M	o->1	
ana T	e->1	
ana a	t->2	v->2	
ana b	e->3	u->1	
ana d	e->6	r->2	y->1	ä->1	
ana e	f->1	n->1	r->1	
ana f	a->4	o->2	r->2	ö->2	
ana g	a->1	r->1	
ana h	a->2	ä->3	
ana i	 ->2	
ana k	o->1	
ana l	ä->1	
ana m	i->1	å->1	
ana o	c->1	m->2	
ana p	a->2	r->3	
ana r	e->4	ä->1	
ana s	i->1	k->2	o->4	t->1	å->1	
ana t	r->1	
ana v	i->1	ä->1	
ana å	s->1	t->1	
ana, 	d->2	
anada	,->2	
anade	 ->2	n->2	
anal,	 ->1	
anal.	 ->1	F->1	
anale	r->4	
analf	a->1	
anali	s->3	
analy	s->58	
anamm	a->4	
anand	e->1	
anane	r->1	
anar 	d->7	e->3	h->1	i->1	j->3	k->9	m->2	o->1	t->1	v->2	Ö->1	
anar,	 ->1	
anas 	a->1	d->1	k->1	n->1	
anat 	d->1	t->2	v->1	
anati	o->1	
anber	 ->2	
anbil	a->8	
anbin	d->1	
anbla	n->2	
anbli	c->1	
anboe	n->1	
anbro	t->1	
anbry	t->1	
anbud	s->4	
anbul	 ->1	
anbun	d->1	
anc, 	d->1	
anca,	 ->1	
ancas	 ->1	
ance,	 ->1	
ance.	.->1	
ancer	!->1	a->1	b->1	
ancis	 ->1	
and -	 ->4	
and 8	0->1	
and E	U->1	
and S	v->1	
and T	i->1	
and a	c->1	l->4	n->21	t->4	v->1	
and b	e->4	i->1	y->1	å->1	
and d	e->15	ä->5	
and e	l->2	n->3	r->1	
and f	o->1	y->1	ö->3	
and g	e->2	o->1	r->1	
and h	a->11	
and i	 ->12	n->4	v->1	
and k	o->2	v->3	ä->1	
and l	a->1	ä->2	
and m	e->51	y->1	å->3	
and n	y->1	ä->4	ö->1	
and o	c->16	m->14	s->6	
and p	a->1	å->4	
and r	e->2	
and s	i->1	j->1	k->3	m->1	o->19	t->4	y->1	ä->4	å->2	
and t	.->1	a->1	i->6	v->1	
and u	n->3	t->3	
and v	a->4	e->1	i->2	ä->1	å->1	
and ä	n->1	r->13	
and ö	v->1	
and),	 ->1	
and, 	5->1	D->1	F->1	I->2	N->1	S->2	d->3	f->2	h->2	k->1	l->1	m->3	o->4	p->1	r->1	s->5	u->2	v->2	
and.A	n->1	
and.D	e->4	i->2	
and.E	m->1	
and.G	e->1	
and.I	 ->2	n->3	r->1	
and.J	a->6	
and.K	o->1	
and.L	å->1	
and.M	e->1	i->1	
and.N	u->1	ä->1	
and.O	m->2	
and.S	o->1	
and.U	p->1	
and.V	i->1	
and.Å	 ->1	
and?F	ö->1	
anda 	a->5	e->1	f->2	l->1	o->1	r->1	s->5	
anda,	 ->5	
anda.	D->1	F->1	H->1	M->1	N->1	
andad	 ->1	e->8	
andah	å->43	
andal	!->1	,->1	a->1	e->5	ö->1	
andam	a->1	
andan	 ->4	
andar	 ->3	d->24	
andas	 ->1	
andat	 ->7	,->3	e->5	p->9	
ande 	"->2	(->30	-->11	1->1	A->2	D->1	E->2	G->5	I->1	J->1	K->3	L->2	M->3	N->1	O->1	P->14	R->3	S->4	a->180	b->55	d->53	e->30	f->147	g->17	h->32	i->97	j->1	k->44	l->20	m->67	n->8	o->132	p->77	r->81	s->116	t->51	u->36	v->29	ä->30	å->36	ö->8	
ande!	 ->6	A->1	J->1	N->1	
ande(	A->1	
ande,	 ->101	
ande.	 ->3	-->1	.->1	A->2	D->21	E->6	F->3	G->1	H->8	I->4	J->23	K->3	L->3	M->8	N->3	O->3	P->2	S->4	T->5	U->1	V->9	Å->1	
ande:	 ->15	
ande;	 ->3	
ande?	F->1	H->2	V->1	
andeb	e->1	ä->1	
andef	r->1	ö->10	
andeh	ö->1	
andek	o->9	
andel	 ->12	,->4	.->3	a->6	e->1	n->2	s->17	
andem	e->5	
anden	 ->146	"->1	,->29	.->23	:->3	;->1	a->37	b->2	s->9	
ander	 ->2	a->5	e->3	l->2	ä->3	
andes	k->114	t->1	
andet	 ->323	)->1	,->17	.->30	;->1	?->1	a->1	s->12	
andev	i->2	
andfu	l->1	
andic	a->1	
andid	a->14	
andie	,->1	
andig	t->2	
andik	a->4	
andin	a->1	
andis	 ->1	
andla	 ->21	.->2	d->10	r->118	s->14	t->7	
andli	g->1	n->186	
andlä	g->1	
andmä	n->1	
andni	n->10	
andom	r->14	
andra	 ->283	,->21	.->7	:->4	;->2	b->2	d->2	g->1	h->1	k->1	r->10	s->2	
andre	 ->1	
andri	n->7	
ands 	b->1	d->1	e->1	g->1	i->2	l->1	n->1	p->1	r->1	å->1	
ands,	 ->1	
andsa	n->1	v->3	
andsb	e->1	y->43	
andsk	a->9	o->5	
andsm	e->6	ä->3	
andsp	l->3	
andsv	ä->1	
andsä	n->1	
andup	p->2	
andut	y->1	
andvi	n->2	
andzi	o->4	
ane o	c->2	
ane, 	R->1	
anele	r->1	
anen 	"->1	f->5	g->1	k->2	m->1	o->4	s->2	
anen,	 ->2	
anen.	 ->1	D->1	E->1	F->1	P->2	V->1	
anens	 ->2	
anent	 ->6	a->2	
aner 	b->1	d->1	f->8	h->1	i->2	o->6	s->2	v->1	
aner"	)->1	
aner,	 ->2	
aner.	-->1	J->1	R->1	V->1	
anera	 ->4	d->14	n->1	r->7	s->6	t->5	
aneri	n->20	
anern	a->22	
anesi	s->1	
anet 	f->1	o->1	t->1	
anet,	 ->2	
anet.	J->1	V->1	
anfal	l->2	
anfat	t->12	
anfly	k->1	
anför	 ->33	a->13	s->1	t->3	
ang a	v->1	
ang b	e->1	
ang e	n->1	
ang f	i->1	r->1	ö->2	
ang g	e->1	l->1	
ang h	a->3	
ang i	n->1	
ang j	a->1	
ang k	a->1	
ang m	e->1	å->1	
ang n	i->1	
ang o	c->4	
ang s	i->1	k->2	t->1	ä->1	
ang u	t->1	
ang ä	r->4	
ang, 	b->1	e->1	i->1	m->2	n->1	o->1	s->1	
ang..	 ->1	
ang.D	e->3	ä->1	
ang.E	n->1	
ang.H	u->1	
ang.J	a->2	
ang.O	c->1	m->1	
ang.Ä	r->1	
angav	 ->1	
ange 	a->2	e->1	h->2	n->1	o->5	p->1	s->2	v->1	
ange,	 ->1	
angel	ä->22	
angem	a->4	
angen	 ->10	,->4	.->1	I->1	b->1	s->3	ä->1	
anger	 ->6	a->2	
anges	 ->6	,->2	.->1	
anget	 ->12	
angiv	a->3	e->1	n->1	
angre	p->6	
angri	p->7	
angrä	n->1	
angåe	n->26	
angår	 ->2	
anhan	g->47	
anhed	r->2	
anhän	g->5	
anhål	l->54	
anhöj	d->4	
ani s	a->1	
ani, 	f->1	i->1	o->1	t->1	
anien	 ->4	,->2	.->1	?->1	s->1	
anife	s->1	
anifr	å->1	
anik 	s->1	
anine	r->1	
aning	 ->17	,->1	.->1	a->6	e->6	s->2	
aninv	å->1	
anio;	 ->1	
anisa	t->43	
anise	r->18	
anism	 ->1	.->1	e->9	
anist	i->2	
anite	t->1	
anitä	r->1	
anium	 ->1	.->1	
anivå	,->1	
anj f	ö->2	
anj m	o->1	
anj.D	e->1	
anjen	 ->1	
anjer	,->1	
anjor	 ->1	
anjäm	k->1	
ank e	n->1	
ank v	ä->1	
ank" 	f->1	
ank- 	e->1	
anka 	o->1	v->1	
anka.	E->1	
ankal	l->9	
ankar	 ->10	,->1	.->4	n->2	
anke 	a->1	l->1	o->1	p->40	r->1	t->2	ä->2	
anke,	 ->2	
ankeb	a->1	
ankef	r->1	
ankeg	å->1	
anken	 ->19	,->2	.->1	:->1	s->1	
ankep	o->1	
anker	 ->3	,->1	n->3	ä->1	
ankes	i->1	
ankfa	r->7	
ankfo	r->1	
ankfö	r->1	
ankir	e->1	
ankla	g->4	
ankny	t->1	
anko.	T->1	
ankom	m->1	s->2	
ankop	p->1	
ankra	 ->1	d->3	r->5	
ankre	n->2	
ankri	k->39	
anksc	h->1	
ankse	k->1	
ankt 	v->1	
ankti	o->8	
anlag	t->1	
anled	e->2	n->48	
anlig	 ->3	a->8	g->1	t->3	
anlit	a->1	
anläg	g->13	
anlän	k->1	t->1	
anlöp	a->1	e->3	
anman	ö->1	
anmar	k->26	
anmäl	a->3	d->1	e->1	n->11	s->2	t->1	
anmär	k->10	
ann d	e->1	
ann e	u->1	
ann o	c->1	
ann t	i->1	
ann ä	r->1	
ann, 	e->1	
ann-g	r->1	
anna 	k->3	m->1	p->1	s->1	v->2	
annab	i->1	
annak	i->2	
annal	a->1	
annan	 ->37	,->4	.->1	s->2	
annar	 ->4	e->1	s->15	
annat	 ->67	,->1	.->4	
annen	 ->15	,->1	.->2	s->7	
anner	l->4	
annes	m->1	
annhe	t->1	
annie	n->14	
annin	g->10	
anniv	å->1	
annla	n->1	
annly	s->1	
annlä	n->1	
annol	i->9	
annor	l->2	s->2	
anns 	a->2	d->1	e->2	f->1	m->3	n->1	o->2	t->1	v->1	
annsa	k->1	
annsk	a->1	
annäm	n->2	
ano P	r->2	
ano o	c->1	
ano u	n->1	
anois	e->1	
anon 	e->1	o->1	
anon,	 ->1	
anon.	E->1	
anon?	K->1	
anone	r->1	
anony	m->4	
anor.	D->1	F->1	J->1	V->1	
anord	n->9	
anos 	t->1	
anos!	 ->1	
anpas	s->14	
anpå 	d->1	
anröj	a->5	t->1	
ans -	 ->1	
ans H	e->1	
ans a	g->1	m->1	n->2	r->5	t->6	v->3	
ans b	a->1	e->15	
ans d	a->2	e->1	
ans e	f->1	g->2	n->1	u->1	
ans f	a->1	i->1	l->1	r->4	u->1	ö->13	
ans g	e->1	r->1	ä->1	
ans h	ä->1	å->1	
ans i	 ->4	n->4	
ans k	o->6	u->1	
ans l	a->2	ä->2	
ans m	a->2	e->28	y->1	
ans n	a->1	
ans o	b->1	c->7	m->1	
ans p	a->3	o->1	å->2	
ans r	e->1	
ans s	k->3	l->3	n->1	o->5	t->2	v->1	
ans t	i->1	
ans u	p->1	t->8	
ans v	a->2	e->1	i->1	o->1	
ans ä	r->1	
ans å	s->1	
ans, 	d->2	e->1	f->1	j->1	m->1	n->2	o->4	s->2	t->1	v->1	ä->2	
ans.D	e->1	ä->1	
ans.E	u->1	
ans.L	å->1	
ans.M	e->1	
ans; 	v->1	
ans?.	H->1	
ansat	 ->2	s->5	t->3	
ansch	 ->2	.->1	e->4	
ansde	p->1	
anse 	a->1	
anse.	E->1	
ansee	n->2	
ansen	 ->19	.->2	l->1	s->1	
anser	 ->197	,->3	.->1	a->8	i->1	n->5	
anses	 ->5	
anset	t->2	
anseu	r->1	
ansie	l->28	r->50	
ansik	t->1	
ansin	n->1	
ansio	n->1	
ansit	i->2	l->3	r->1	t->1	
ansiä	r->1	
ansjo	v->17	
ansk 	d->1	l->2	n->1	p->2	r->1	
anska	 ->117	,->2	.->2	d->3	f->1	r->5	s->5	t->4	
anske	 ->64	,->1	
anskl	i->1	
anskn	i->23	
ansko	n->9	
anskr	ä->1	
anskt	 ->4	.->1	a->1	
ansku	l->1	
ansla	g->23	
ansle	r->1	
ansli	e->1	
anslo	g->1	
anslu	t->29	
anslå	 ->1	d->1	r->1	s->2	
ansmi	n->1	
ansmä	l->1	n->5	
anspe	l->1	
anspo	r->108	
anspr	å->7	
ansrä	t->22	
ansta	l->1	n->2	t->5	
ansto	r->2	
anstr	ä->46	
anstä	l->33	n->5	
anstå	e->1	
ansva	r->306	
ansvä	r->11	
ansät	t->5	
ansåg	 ->12	
ansåt	g->1	
ansök	a->8	n->1	t->1	
ansöv	n->1	
ant -	 ->3	
ant E	u->2	
ant a	n->1	r->1	t->9	v->1	
ant b	e->2	i->1	
ant c	e->1	
ant d	e->3	i->1	
ant f	a->4	i->1	r->2	u->1	ö->9	
ant g	a->1	
ant h	a->2	
ant i	 ->2	f->1	n->2	
ant k	o->3	r->1	
ant m	ö->1	
ant n	u->1	y->1	ä->1	
ant o	c->2	m->3	
ant p	r->3	å->1	
ant s	a->1	e->1	k->1	l->1	o->7	t->3	y->2	ä->7	å->1	
ant t	e->1	i->2	
ant u	n->1	t->1	
ant ä	m->1	r->1	
ant ö	v->1	
ant!"	J->1	
ant, 	d->2	f->1	h->2	i->1	o->1	
ant.D	e->2	
ant.H	e->1	
ant.S	a->1	
ant.V	i->1	
ant: 	v->1	
anta 	-->1	1->1	M->1	S->1	a->1	b->1	d->4	e->7	f->2	k->4	l->1	m->3	n->1	o->1	s->2	t->1	u->1	ä->2	å->1	
antab	r->3	
antag	 ->12	,->4	.->2	?->1	a->13	e->6	i->18	l->1	n->4	s->10	
antal	 ->40	,->1	e->17	
antar	 ->9	
antas	 ->10	,->2	.->1	i->2	t->9	
antat	i->1	
ante 	e->1	f->2	
ante,	 ->2	
anten	 ->6	)->1	.->1	?->1	
anter	 ->8	,->1	-->1	.->3	a->80	i->20	n->1	
anti 	f->5	i->1	o->2	s->1	
anti,	 ->1	
anti-	g->1	i->1	r->1	
anti.	H->1	
antib	e->1	
antid	e->1	
antie	l->2	r->15	u->1	
antif	a->3	i->4	o->3	
antik	a->1	o->1	r->2	
antim	ö->1	
antin	 ->3	g->11	
antiq	u->1	
antis	e->5	k->6	y->1	
antit	a->4	r->1	
antku	s->1	
antli	g->3	
antni	n->1	
antog	 ->13	s->10	
antor	,->1	
antra	 ->2	t->1	
anträ	d->34	t->1	
antve	r->2	
antyd	d->2	
antör	e->2	s->1	
anuar	i->16	
anuts	-->1	
anvap	e->4	
anvis	a->1	
använ	d->174	t->10	
anyon	 ->2	,->1	
anz F	i->3	
anzes	-->1	
ançoi	s->1	
anöst	e->19	
anövr	a->1	
ao ti	l->1	
aordi	n->1	
aos n	ä->1	
aos o	c->1	
ap - 	o->1	
ap at	t->2	
ap av	 ->20	
ap bö	r->2	
ap de	n->1	
ap dä	r->2	
ap el	l->1	
ap fr	å->1	
ap fö	r->2	
ap gr	u->1	
ap ha	r->1	
ap i 	f->1	r->2	u->1	v->1	
ap in	l->1	t->1	
ap ko	m->1	
ap me	l->1	
ap må	s->1	
ap nä	r->1	
ap oc	h->12	
ap om	 ->3	
ap sk	a->1	u->1	
ap so	m->9	
ap ti	l->1	
ap un	d->1	
ap up	p->1	
ap va	d->1	
ap är	 ->1	
ap" f	r->1	
ap"!I	 ->1	
ap", 	v->1	
ap, d	e->1	ä->1	
ap, e	n->3	
ap, f	o->1	ö->1	
ap, h	a->1	
ap, i	n->1	
ap, o	c->2	m->1	
ap, u	t->1	
ap, v	a->1	i->1	
ap, ä	v->1	
ap. S	k->1	
ap.Da	g->1	
ap.De	t->6	
ap.Eu	r->1	
ap.I 	d->1	o->1	
ap.Ja	g->2	
ap.Sl	u->1	
ap.Ti	l->1	
ap.Vi	 ->2	
ap: K	o->1	
apa O	L->1	
apa a	r->2	
apa b	e->2	ä->1	
apa d	e->3	r->1	
apa e	f->1	n->22	r->1	t->14	u->1	
apa f	l->2	r->1	ö->5	
apa g	e->1	
apa h	å->1	ö->2	
apa i	m->1	n->2	
apa j	ä->1	
apa k	l->1	o->2	u->1	v->1	
apa l	u->1	
apa n	y->5	å->3	
apa o	c->1	m->1	
apa r	ä->1	
apa s	n->1	p->1	t->1	y->5	å->1	
apa t	i->1	r->3	v->2	
apa v	ä->1	
apa y	t->1	
apa ä	n->1	
apaci	t->5	
apade	 ->2	s->3	
apan 	e->1	o->1	
apan,	 ->1	
apand	e->24	
apans	k->1	
apar 	a->1	b->1	d->1	e->6	f->1	i->2	k->1	m->1	n->1	o->1	s->3	v->5	ö->1	
apar.	D->1	I->1	
apare	 ->2	
aparl	a->166	
apas 	a->2	e->2	f->3	i->4	l->1	m->1	
apat 	d->1	e->3	n->2	s->1	
apat.	F->1	
apats	 ->2	
apaya	n->2	
apeau	"->1	
apen 	(->2	-->1	a->2	b->1	e->4	f->2	g->2	h->3	i->2	k->2	m->3	n->2	o->10	p->1	s->6	u->3	v->2	ä->4	å->2	
apen,	 ->10	
apen.	 ->1	D->1	H->1	J->1	K->1	M->2	N->2	S->1	T->1	
apen?	.->1	
apenh	a->1	
apeni	n->1	
apens	 ->71	p->1	
apent	e->1	
apenu	t->1	
aper 	h->1	o->2	v->1	
aper,	 ->1	
aper.	E->1	
aperi	f->1	
apern	a->16	
apest	 ->1	
apet 	(->1	-->1	a->1	b->2	d->2	f->6	g->1	h->3	i->2	k->11	l->1	m->5	n->2	o->8	p->2	r->1	s->6	t->3	v->3	
apet)	 ->1	
apet,	 ->13	
apet.	H->1	J->1	M->2	N->1	P->1	
apet?	R->1	
apets	 ->15	
apita	 ->6	,->1	.->3	l->17	
apite	l->6	
apitu	l->2	
apkay	 ->3	,->3	.->1	D->1	b->1	s->2	
aplan	,->1	
aplig	 ->10	a->25	h->1	t->1	
apnen	 ->2	
apoli	t->2	
app d	ä->1	
app h	ö->1	
app u	t->1	
app, 	i->1	
app.V	i->1	
appa 	e->1	i->1	m->1	r->1	
appad	e->3	
appar	 ->2	a->1	
appas	t->9	
appel	l->1	
appen	 ->1	
apper	 ->4	.->1	:->1	e->1	s->1	
apphe	t->3	
appja	k->1	
appla	n->2	
applå	d->6	
appni	n->1	
appor	t->112	
appss	t->1	
appt 	e->2	i->1	s->1	t->1	
appve	r->2	
appy 	e->1	
april	 ->2	.->1	
aprob	l->1	
aproc	e->2	
aprod	u->1	
aproj	e->1	
aprop	å->1	
aps f	a->1	
aps- 	o->1	
apsav	t->2	
apsbe	f->1	g->1	s->1	
apsdi	r->1	
apsfr	å->1	
apsin	i->7	s->6	t->1	
apsko	n->3	
apsla	g->3	
apsma	s->2	
apsme	d->1	
apsmä	n->16	
apsmå	l->1	
apsni	v->11	
apsor	g->1	
apspe	l->2	
apspo	l->2	
apspr	o->3	
apsra	m->1	
apsre	g->9	
apsrä	t->8	
apsst	r->1	ö->2	
apssy	s->1	
apsåt	g->2	
apten	 ->2	
ar "ö	v->1	
ar (C	5->2	
ar (F	I->1	
ar - 	a->1	d->1	e->2	f->1	h->1	k->1	m->1	s->2	u->1	v->1	ä->1	
ar 1,	4->1	
ar 10	 ->1	
ar 13	0->1	
ar 15	 ->2	
ar 17	4->1	
ar 19	2->1	9->2	
ar 26	2->1	
ar 3-	4->1	
ar 40	 ->1	
ar 97	.->1	
ar Al	b->1	t->1	
ar BN	P->1	
ar Br	o->2	
ar Ce	n->1	
ar Eu	r->14	
ar Ev	a->1	
ar Fl	o->1	
ar Fö	r->1	
ar Go	l->1	
ar In	t->1	
ar Ku	m->1	
ar La	n->1	
ar Lo	t->2	
ar Ly	n->1	
ar Pa	l->1	
ar Po	n->1	
ar Pr	o->1	
ar RE	P->1	
ar Rh	ô->1	
ar Ro	t->1	
ar Rå	d->1	
ar Se	g->1	
ar So	l->1	
ar Sw	o->1	
ar Th	e->1	
ar Wa	l->1	
ar ab	s->1	
ar ac	c->2	
ar ag	e->1	
ar ak	t->3	
ar al	d->5	l->39	
ar an	a->5	d->1	k->1	l->1	m->1	o->1	s->22	t->11	v->6	
ar ar	b->6	t->1	
ar as	"->1	
ar at	t->128	
ar av	 ->55	g->4	i->2	l->1	s->5	v->2	
ar ba	n->2	r->9	
ar be	a->2	d->1	f->7	g->8	h->7	k->1	l->2	r->4	s->16	t->12	v->3	
ar bi	d->5	f->1	l->4	s->1	
ar bl	a->3	i->18	
ar bo	m->1	
ar br	a->1	i->3	o->1	u->1	å->2	ö->1	
ar bu	d->1	
ar by	g->3	r->1	
ar bä	t->4	
ar bå	d->2	
ar bö	r->7	
ar ci	r->1	
ar co	p->1	
ar da	g->1	
ar de	 ->61	,->1	b->17	f->1	l->11	m->9	n->63	r->1	s->29	t->109	
ar di	r->1	s->10	
ar do	c->5	m->2	
ar dr	a->8	i->1	
ar dä	r->33	
ar då	 ->5	
ar dö	r->1	t->1	
ar ef	f->2	t->13	
ar eg	e->1	
ar ek	o->2	
ar el	l->10	
ar em	e->4	o->5	
ar en	 ->94	a->2	d->4	e->5	g->1	h->2	i->1	l->6	o->1	s->3	
ar er	 ->7	,->3	.->1	a->1	f->1	h->2	k->1	s->2	t->1	
ar et	a->1	t->56	
ar eu	r->2	
ar ex	a->1	e->2	i->1	p->1	t->5	
ar fa	k->3	l->2	r->4	s->3	t->4	
ar fe	l->2	
ar fi	n->4	s->2	
ar fl	a->1	e->5	y->4	
ar fo	r->6	
ar fr	a->29	i->4	ä->2	å->19	
ar fu	l->1	n->7	
ar fä	s->1	
ar få	t->28	
ar fö	l->5	r->207	
ar ga	g->2	r->1	
ar ge	m->2	n->15	t->11	
ar gi	l->1	v->5	
ar gj	o->46	
ar gl	ö->2	
ar go	d->8	
ar gr	a->2	i->1	u->1	
ar gä	l->1	r->2	
ar gå	n->1	r->2	t->11	
ar gö	m->1	r->1	
ar ha	 ->4	f->16	k->1	l->1	m->1	n->6	r->8	v->1	
ar he	l->20	n->3	t->1	
ar hi	t->10	
ar hj	ä->1	
ar ho	n->4	s->3	t->1	
ar hu	r->4	
ar hä	n->7	r->10	v->3	
ar hå	l->6	
ar hö	g->1	r->13	
ar i 	E->15	I->1	K->2	L->1	T->1	W->1	a->7	b->3	d->34	e->10	f->12	g->1	h->1	i->1	k->2	m->6	n->2	o->4	p->4	r->1	s->17	t->3	u->5	v->5	Ö->1	ä->1	ö->2	
ar i.	A->1	
ar ia	n->1	
ar id	e->4	
ar if	r->1	
ar ig	e->4	
ar ih	o->1	
ar in	 ->3	b->1	d->1	f->9	g->18	i->2	k->1	l->5	n->4	o->7	r->1	s->2	t->99	v->2	
ar is	c->1	
ar it	u->6	
ar iv	ä->1	
ar ja	g->78	
ar ju	 ->13	r->1	s->10	
ar ka	l->3	m->1	n->9	
ar kl	a->3	i->1	o->1	y->1	
ar ko	m->66	n->14	r->3	s->1	
ar kr	a->2	e->1	i->3	ä->1	
ar ku	l->3	n->12	
ar kv	a->2	i->1	
ar kä	m->1	
ar kö	r->2	
ar la	g->36	n->1	
ar le	 ->1	g->2	t->7	
ar li	d->3	g->1	k->2	s->1	t->1	v->2	
ar lo	v->4	
ar lu	r->1	
ar ly	c->13	f->1	s->4	
ar lä	c->1	g->1	m->8	n->5	r->1	s->1	t->1	
ar lå	n->1	s->1	t->1	
ar lö	n->2	p->3	s->1	
ar ma	n->41	r->3	
ar me	d->90	l->4	n->2	r->4	t->1	
ar mi	g->23	l->8	n->16	s->3	t->1	
ar mo	d->3	n->1	t->11	
ar my	c->12	n->2	
ar mä	n->4	
ar må	n->5	r->1	s->3	
ar mö	j->8	
ar na	k->1	t->7	
ar ne	d->2	k->1	
ar ni	 ->11	v->1	
ar no	r->1	t->4	
ar nu	 ->16	,->1	.->1	
ar ny	a->4	l->2	t->3	
ar nä	m->10	r->13	s->1	
ar nå	g->30	t->4	
ar nö	d->3	j->2	
ar oa	c->1	v->1	
ar ob	s->1	
ar oc	h->110	k->44	
ar oe	n->1	
ar of	f->2	t->4	
ar ok	u->1	
ar ol	i->4	ö->1	
ar om	 ->125	,->5	.->6	b->1	v->1	
ar or	d->9	s->2	ä->1	
ar os	s->24	
ar pa	p->1	r->13	
ar pe	k->3	n->3	r->2	
ar pl	a->1	
ar po	l->4	
ar pr	a->1	e->4	i->1	o->9	
ar pu	n->4	
ar på	 ->90	b->2	f->1	p->7	s->1	t->3	v->5	
ar ra	p->1	t->3	
ar re	a->1	d->24	f->2	g->6	j->1	k->1	n->2	s->2	
ar ri	k->1	s->2	
ar ry	c->1	
ar rä	d->1	k->3	t->18	
ar rå	d->14	
ar rö	r->4	s->6	
ar sa	g->18	k->2	m->17	n->1	t->4	
ar se	 ->2	d->7	g->1	n->1	t->8	x->1	
ar si	g->45	n->15	t->3	
ar sj	ä->5	
ar sk	a->17	e->5	i->5	j->4	o->1	r->5	u->6	y->2	ö->1	
ar sl	a->1	u->6	
ar sm	u->1	
ar sn	e->1	
ar so	m->101	
ar sp	e->7	r->1	å->1	
ar st	a->4	i->1	o->10	r->3	y->2	ä->7	å->6	ö->9	
ar su	b->3	
ar sv	a->3	å->1	
ar sy	s->4	
ar sä	g->2	k->7	r->5	t->1	
ar så	 ->13	,->1	d->2	l->5	
ar ta	 ->1	g->23	l->7	s->1	
ar te	k->1	m->1	n->1	
ar ti	d->7	l->113	o->2	
ar tj	ä->2	
ar to	l->1	
ar tr	a->2	e->2	o->3	ä->1	å->1	
ar tu	s->1	
ar tv	u->4	ä->1	å->4	
ar ty	d->4	v->4	
ar tä	n->1	r->1	
ar un	d->20	g->1	i->3	
ar up	p->43	
ar ur	 ->1	
ar ut	 ->2	,->1	.->1	a->9	f->6	g->3	i->2	l->2	n->2	r->1	s->2	t->3	v->17	ö->1	
ar va	d->4	l->5	n->2	r->39	
ar ve	l->1	r->18	t->4	
ar vi	 ->123	,->3	d->10	g->1	k->1	l->2	s->17	t->1	
ar vu	n->1	
ar vä	c->4	l->8	n->3	s->2	x->1	
ar vå	r->14	
ar yt	t->2	
ar ÖV	P->1	
ar äg	n->2	t->3	
ar äl	d->1	
ar äm	n->1	
ar än	 ->6	d->11	n->5	
ar är	 ->26	a->2	
ar äv	e->10	
ar å 	a->1	
ar ål	a->1	
ar år	 ->3	
ar ås	a->1	t->1	
ar åt	 ->1	e->3	g->1	s->1	t->1	
ar ök	a->6	
ar ön	s->2	
ar öp	p->1	
ar ös	t->2	
ar öv	a->1	e->28	
ar! A	v->1	
ar! B	l->1	
ar! D	e->2	
ar! E	r->1	
ar! F	ö->3	
ar! H	i->1	
ar! J	a->4	
ar! N	å->1	
ar! P	P->1	
ar! S	o->2	
ar! T	i->1	
ar! V	i->1	
ar!De	t->1	
ar!Ja	g->1	
ar!Me	d->1	
ar!Mi	n->1	
ar!Ti	l->1	
ar" m	å->1	
ar" o	c->1	
ar).)	B->1	
ar, P	a->1	
ar, T	y->1	
ar, W	a->1	
ar, a	l->3	n->2	r->1	t->5	v->1	
ar, b	i->1	l->1	å->1	
ar, d	e->5	v->4	ä->2	å->2	
ar, e	f->4	l->1	n->2	r->1	t->1	
ar, f	o->1	r->3	ö->9	
ar, g	e->1	y->1	
ar, h	a->1	e->1	
ar, i	 ->4	c->1	n->5	
ar, j	a->3	ä->2	
ar, k	a->1	o->7	r->2	ä->4	
ar, l	i->5	ä->1	å->2	
ar, m	a->2	e->14	y->1	å->1	
ar, n	e->1	i->1	ä->2	å->1	
ar, o	c->32	l->1	m->5	
ar, p	r->1	å->3	
ar, r	ä->1	
ar, s	a->2	n->1	o->13	å->4	
ar, t	i->3	
ar, u	n->3	t->7	
ar, v	a->2	i->8	
ar, ä	n->1	r->6	v->2	
ar, å	t->3	
ar- s	o->1	
ar. A	l->1	
ar. E	f->1	
ar. M	e->1	
ar. V	å->1	
ar.)S	ä->1	
ar.- 	(->1	
ar.. 	(->2	
ar...	H->1	
ar.Am	e->1	
ar.At	t->1	
ar.Ba	r->1	
ar.Be	f->1	
ar.Bl	a->1	
ar.Bo	s->1	
ar.De	 ->10	n->10	s->2	t->37	
ar.Dä	r->4	
ar.Då	 ->1	
ar.Ef	t->2	
ar.En	 ->1	l->1	
ar.Er	f->1	
ar.Eu	r->2	
ar.FP	Ö->1	
ar.Fr	e->1	
ar.Fö	r->14	
ar.Ge	m->1	n->1	
ar.Gö	r->1	
ar.He	r->7	
ar.Hu	r->1	
ar.Hä	r->1	
ar.I 	I->2	R->1	a->2	d->1	r->1	s->2	v->1	
ar.In	d->1	g->1	r->1	t->1	
ar.Ja	g->32	
ar.Ko	m->2	n->1	
ar.Kr	a->1	
ar.Li	k->1	
ar.Lå	t->2	
ar.Ma	n->2	
ar.Me	d->1	l->1	n->6	
ar.Mi	n->1	
ar.Na	t->1	
ar.Ni	v->1	
ar.Nå	g->1	
ar.Ob	e->1	
ar.Oc	h->2	
ar.Om	 ->6	
ar.På	 ->2	
ar.Re	n->1	
ar.Ri	s->1	
ar.Rä	k->1	
ar.Rå	d->1	
ar.Se	d->2	
ar.Sk	u->1	
ar.So	m->1	
ar.St	ö->1	
ar.Så	 ->2	
ar.Ta	c->2	
ar.Ti	l->3	
ar.Un	d->1	
ar.Ut	e->1	
ar.Va	r->1	
ar.Vi	 ->27	d->1	
ar.Vå	r->1	
ar.Än	d->2	
ar: D	e->1	
ar: F	r->1	
ar: P	å->1	
ar: a	n->2	
ar: d	e->3	
ar: f	ö->1	
ar: o	p->1	
ar: u	t->1	
ar: v	i->2	
ar; i	 ->1	n->1	
ar; m	e->1	
ar; o	c->1	
ar?I 	e->1	
ar?Ja	g->1	
ar?Ka	n->1	
ar?Ko	m->1	
ar?Na	t->1	
ar?Ni	 ->1	
ara "	b->1	u->1	
ara 1	 ->1	0->1	5->1	
ara 2	 ->1	
ara 5	5->1	
ara 7	0->1	
ara B	a->1	
ara D	a->1	
ara E	u->2	
ara I	s->1	
ara a	d->1	k->1	l->2	m->1	n->4	r->1	t->16	u->1	v->15	
ara b	a->1	e->15	i->1	l->2	r->4	ä->2	
ara c	e->2	
ara d	a->1	e->24	i->1	j->2	o->1	r->1	u->1	ö->1	
ara e	f->3	l->1	m->1	n->75	r->1	t->28	u->4	x->2	
ara f	a->7	e->3	l->1	o->1	r->4	u->2	ä->1	å->1	ö->43	
ara g	e->5	i->1	l->2	o->2	r->1	ä->3	å->1	ö->2	
ara h	a->5	e->6	i->1	o->1	u->4	ä->3	
ara i	 ->13	a->1	c->1	h->1	l->2	n->4	
ara j	a->1	u->2	ä->1	
ara k	a->4	l->1	n->1	o->16	r->2	v->1	ä->1	
ara l	a->4	e->1	i->6	ä->6	ö->1	
ara m	e->23	i->5	o->4	y->17	ä->1	å->5	ö->4	
ara n	a->3	y->2	ä->9	å->11	ö->8	
ara o	b->4	c->8	f->2	m->10	n->1	r->3	s->1	t->1	
ara p	a->2	e->1	o->1	r->3	å->12	
ara r	e->5	i->4	o->1	ä->3	
ara s	a->7	i->3	j->1	k->11	m->1	n->1	t->6	u->1	v->1	y->2	ä->8	å->14	
ara t	a->4	e->1	i->19	j->1	o->1	r->3	v->1	y->2	
ara u	n->6	p->5	r->1	t->7	
ara v	a->8	i->14	o->1	ä->7	å->1	
ara y	t->3	
ara Ö	s->1	
ara ä	g->1	n->1	r->16	
ara å	 ->1	t->2	
ara ö	n->1	v->6	
ara".	D->1	
ara, 	a->1	b->1	f->2	m->1	o->1	u->1	
ara.A	l->1	v->1	
ara.D	e->2	
ara.F	ö->1	
ara.J	a->2	
ara.M	å->1	
ara.P	å->1	
ara.V	i->1	
ara: 	V->1	s->1	
ara?D	e->1	
arabi	s->6	
arabl	a->1	
arabs	t->2	
arad 	e->1	ä->1	
arade	 ->10	.->1	r->1	s->3	
arado	x->6	
aragr	a->3	
arak 	h->2	i->1	l->1	v->1	
arak.	T->1	
araks	 ->3	
arakt	e->2	i->4	ä->9	
arall	e->5	
arame	t->2	
aran 	f->2	v->1	
aran.	D->1	
arand	a->2	e->275	r->10	
arann	a->1	
arans	v->6	
arant	 ->2	e->57	i->34	
arar 	E->2	R->1	S->1	a->8	b->1	d->26	f->8	h->2	i->2	j->2	k->1	m->4	n->1	p->2	s->1	u->1	v->3	ä->1	
arar,	 ->1	
arare	 ->26	
aras 	a->3	b->1	f->1	i->1	m->1	o->1	r->1	s->2	
arast	 ->12	.->1	
arat 	a->1	d->1	e->1	f->1	k->2	s->1	t->1	
arate	n->1	
arati	o->1	
arats	 ->4	
arav 	4->1	8->1	d->1	e->1	
arbar	i->2	
arbas	t->1	
arbet	a->133	e->214	s->217	
arcel	o->2	
arcou	r->1	
ard C	o->1	
ard K	o->1	
ard e	u->1	
ard f	ö->1	
ard o	c->1	
ard p	å->1	
ard s	j->1	k->1	
ard v	a->1	
ard, 	d->1	o->2	
ard-a	f->1	
ard.D	e->1	
ard; 	i->1	
ardag	,->1	e->1	l->2	
arde-	l->1	
ardem	o->1	
arden	 ->3	
arder	 ->16	.->1	a->2	
ardis	e->9	
are -	 ->3	
are 1	1->1	5->1	
are 2	1->1	
are 3	5->1	
are 4	,->1	
are D	e->1	i->1	
are E	u->2	
are a	d->1	l->1	n->4	t->23	v->10	
are b	a->1	e->20	i->2	l->4	y->2	ö->1	
are d	a->2	e->6	i->2	o->1	y->1	ä->1	å->1	
are e	f->1	k->2	l->6	m->1	n->8	t->4	
are f	a->2	e->1	i->2	l->1	o->1	r->26	y->2	å->3	ö->53	
are g	e->4	j->1	o->1	r->1	å->1	ö->1	
are h	a->18	e->1	i->2	u->2	å->1	ö->2	
are i	 ->33	n->14	
are j	o->1	
are k	a->12	o->17	r->2	u->2	ä->1	
are l	i->1	ä->1	ö->1	
are m	a->1	e->11	i->1	o->3	å->5	
are n	i->1	u->1	ä->7	å->2	
are o	c->35	m->7	r->1	
are p	a->1	e->2	l->1	o->2	r->5	å->12	
are r	e->7	i->1	o->1	ä->1	
are s	a->5	e->2	i->13	k->13	o->34	t->4	y->2	ä->1	å->1	
are t	a->6	i->21	r->1	v->3	
are u	n->2	p->3	t->7	
are v	a->3	e->1	i->5	ä->1	
are ä	n->23	r->8	
are å	r->3	t->2	
are ö	k->2	
are!S	k->1	
are" 	s->2	
are",	 ->1	
are, 	F->1	H->1	a->3	b->5	d->2	e->1	f->3	h->4	i->3	j->1	k->2	m->10	n->3	o->10	p->5	s->10	u->2	v->6	ä->3	å->2	
are. 	D->1	O->1	Ä->1	
are.A	l->1	t->1	
are.B	å->1	
are.D	e->15	ä->2	å->2	
are.E	f->2	u->2	
are.F	ö->2	
are.H	e->1	
are.I	 ->2	m->1	
are.J	a->6	
are.K	o->2	
are.M	a->2	e->2	i->2	
are.N	u->1	
are.P	å->1	
are.R	o->1	
are.S	o->2	
are.T	i->1	r->1	
are.U	r->1	
are.V	a->1	i->4	å->1	
are.Ä	n->2	r->1	v->1	
are: 	d->1	
are?D	e->1	
are?K	a->1	
are?O	c->1	
arebe	f->2	h->1	
areft	e->1	
arela	 ->1	
arelä	g->2	
arems	a->2	
aren 	H->1	K->1	V->1	a->9	b->2	e->5	f->7	g->1	h->3	i->6	k->1	l->1	m->2	o->10	p->3	r->2	s->10	t->1	v->2	ä->7	å->1	ö->1	
aren)	.->1	J->1	
aren,	 ->17	
aren.	)->5	.->1	A->1	D->4	F->1	H->2	I->2	J->2	M->1	O->2	T->1	V->1	
aren;	 ->1	
aren?	Ä->1	
arend	a->2	
arenh	e->24	
arens	 ->4	/->1	
arent	s->1	
arepr	e->1	
arer 	a->1	e->1	h->1	i->3	m->1	o->5	s->2	v->1	
arer,	 ->3	
arer.	T->1	V->1	
arera	 ->4	
arern	a->1	
ares 	a->2	d->1	f->1	i->2	l->2	n->1	o->2	p->1	r->3	å->1	ö->1	
ares,	 ->3	
aret 	a->3	f->24	h->1	i->3	l->2	o->9	p->1	r->1	s->1	t->1	v->1	ä->6	å->1	
aret,	 ->2	
aret.	D->4	E->1	F->1	I->1	J->3	L->1	M->1	T->2	V->2	
areur	o->1	
areut	b->1	v->3	
arfor	d->1	
arfär	g->1	
arför	 ->46	,->1	:->1	?->3	m->1	
arga 	f->1	
argan	i->5	
argar	i->1	n->1	
argin	a->6	
argo 	s->1	
argot	 ->1	
argum	e->17	
argör	 ->2	a->13	s->2	
arhet	 ->11	.->3	e->7	
arhus	,->1	
arhän	g->1	
arhåg	o->2	
arhål	l->2	
ari 1	9->4	
ari 2	0->5	
ari e	n->1	t->1	
ari f	ö->1	
ari i	 ->1	n->2	
ari m	å->1	
ari n	ä->1	
ari o	c->2	m->1	
ari!H	e->1	
ari, 	m->2	o->4	s->3	v->1	
ari.H	u->1	
ari.V	i->1	
aria 	d->1	
ariat	 ->1	.->1	
arici	o->1	
arie 	C->1	
arien	.->1	
arier	,->1	a->2	
ariet	s->1	
arig 	a->1	b->1	f->14	k->1	m->1	
arig,	 ->3	
ariga	 ->25	,->2	.->2	
arige	 ->1	
arigh	e->5	
arigt	 ->5	,->1	
arike	r->9	t->15	
arin 	o->1	
aring	 ->13	,->1	.->3	a->4	e->6	
arinh	o->6	
arinn	a->1	
ario 	f->1	
arior	.->1	
ariot	 ->2	
aris 	s->1	
aris,	 ->1	
arise	r->3	
arisf	ö->1	
arisk	 ->7	a->9	t->2	
arism	 ->2	.->2	e->2	
arist	i->2	
arit 	a->2	b->2	d->1	e->13	f->7	g->1	h->3	i->5	k->4	l->2	m->8	n->2	o->2	p->4	r->2	s->9	t->3	u->1	v->2	
arite	t->53	
ariti	m->3	
arium	 ->2	
arje 	1->1	E->1	a->3	b->3	d->9	e->7	f->15	g->5	h->2	i->3	k->2	l->9	m->11	o->1	r->3	s->6	å->10	
ark -	 ->1	
ark b	e->1	
ark e	l->2	n->1	
ark f	ö->2	
ark h	a->1	
ark i	 ->1	n->2	
ark k	o->3	ä->1	
ark l	y->1	
ark m	å->1	
ark o	c->5	f->1	
ark p	o->2	å->2	
ark s	k->2	o->2	å->1	
ark t	i->2	r->1	
ark v	i->3	
ark, 	d->1	g->1	o->1	ä->1	
ark.D	e->1	å->1	
ark.F	r->1	
ark.J	a->1	
arka 	i->2	k->1	l->1	m->1	n->1	o->3	p->1	r->1	s->1	t->1	
arka,	 ->1	
arkan	t->3	
arkar	 ->1	e->6	
arkas	s->2	t->5	
arkbo	r->1	
arke 	m->1	
arken	 ->19	.->1	
arker	a->7	i->3	
arket	 ->1	
arki.	D->1	
arkin	 ->1	.->1	
arkis	k->1	
arkiv	 ->1	e->1	
arkla	s->1	
arkna	d->191	
arkol	l->1	
arkom	a->1	
arkon	f->1	t->2	
arkot	i->7	
arkov	 ->1	
arks 	o->1	t->1	
arkt 	E->1	b->3	d->1	f->2	m->5	p->1	s->4	v->1	ö->3	
arkt,	 ->1	
arkt.	D->1	
arl H	e->1	
arl v	o->3	
arl-H	e->1	
arlag	d->1	t->2	
arlam	e->600	
arlan	d->3	
arled	i->1	
arlig	 ->14	,->2	:->1	a->43	e->12	t->62	
arlik	a->1	
arlsr	u->2	
arläg	g->2	
arläk	t->1	
arlän	d->7	
arløn	,->2	
arm e	l->4	
arm-e	l->1	
arma 	f->1	k->1	å->1	
armac	e->1	
armad	e->4	
armak	o->1	
arman	d->1	
armat	 ->6	
armod	 ->1	
armon	i->18	
armra	p->2	
armsi	g->2	
armst	a->1	
armt 	a->1	d->1	e->1	o->3	t->5	v->1	
armyn	d->14	
armé 	o->1	
armén	 ->1	.->1	
arn -	 ->1	
arn i	n->1	
arn k	o->1	
arn o	c->2	
arn s	k->1	o->1	å->1	
arn, 	m->2	o->1	
arna 	-->4	1->1	6->1	8->8	a->30	b->6	d->9	e->10	f->43	g->7	h->15	i->61	k->12	l->2	m->13	n->5	o->47	p->9	r->1	s->33	t->10	u->5	v->6	ä->13	ö->3	
arna!	O->1	
arna"	.->1	i->1	
arna,	 ->43	
arna.	 ->1	(->1	A->1	D->19	E->2	F->8	H->2	I->3	J->5	K->2	L->1	M->4	O->1	S->2	T->1	U->3	V->6	Ä->1	
arna?	H->1	J->1	V->1	
arnad	e->1	
arnag	e->1	
arnar	 ->3	
arnas	 ->65	,->1	
arnba	r->1	
arnhi	l->1	
arnie	r->14	
arnin	g->7	
arnpo	r->2	
arns 	f->1	
aro -	 ->1	
aro i	 ->1	
aro n	å->1	
aro v	a->1	
aro, 	t->1	
aron 	a->2	
aron,	 ->1	
aror 	o->1	s->2	
aror,	 ->1	
aror.	N->1	V->1	
arouk	 ->1	
arpar	t->1	
arpeg	n->1	
arpol	-->1	
arpt 	d->1	f->1	
arr i	 ->1	
arran	g->6	
arres	t->2	
arris	 ->1	
arriä	r->4	
arrog	a->2	
ars 1	9->1	
ars 2	0->1	
ars E	U->1	
ars a	n->1	
ars b	e->3	
ars d	ö->1	
ars e	f->1	k->1	
ars f	l->4	ö->2	
ars g	i->1	r->1	
ars h	a->2	j->1	ä->1	
ars i	 ->3	n->1	
ars k	a->2	o->3	
ars l	ä->1	
ars m	å->3	
ars n	a->1	i->1	
ars o	a->1	c->1	f->1	r->1	
ars p	a->1	r->1	
ars r	e->1	o->1	
ars s	i->1	k->3	o->1	y->1	
ars t	a->1	r->1	
ars u	p->1	t->3	
ars v	ä->1	
ars ä	g->1	r->1	
ars å	t->1	
ars, 	e->1	k->1	o->2	
ars.D	e->1	
ars.N	u->1	
ars.V	i->1	
arsam	m->6	
arsav	g->1	
arsbe	f->2	
arsbu	d->1	
arsch	e->1	
arsei	l->1	
arsfr	i->43	å->4	
arsfu	l->4	
arsfö	r->4	
arska	p->9	
arsku	l->1	
arskä	n->3	
arsla	n->1	
arsma	k->1	
arsme	d->1	
arsmi	n->1	
arsom	r->6	
arsor	d->1	
arsot	 ->1	
arspo	l->4	s->1	
arsta	d->1	g->1	
arsti	d->1	
arsto	l->1	
arstå	r->6	t->1	
arsyd	d->1	
art -	 ->3	
art E	u->2	
art a	g->1	t->53	v->4	
art b	a->1	e->3	ä->1	
art d	e->2	
art e	m->1	n->3	
art f	a->4	i->1	r->1	å->2	ö->17	
art g	e->3	
art h	a->1	o->3	u->2	
art i	 ->6	n->6	
art k	o->5	
art l	y->1	ä->1	
art m	a->4	e->3	å->1	
art n	ä->1	å->1	
art o	c->12	m->3	
art p	a->1	o->1	r->1	å->1	
art r	e->1	
art s	k->3	l->1	o->15	p->1	t->2	y->1	ä->6	å->2	
art t	e->2	i->1	o->1	r->1	
art u	n->1	t->2	
art v	a->1	i->1	
art Ö	s->1	
art ä	r->4	
art!H	e->1	
art, 	h->1	l->1	m->2	o->2	s->1	v->1	
art. 	7->1	
art.A	r->1	
art.D	e->1	
art.F	r->1	ö->1	
art.H	ä->1	
art.I	 ->1	
art.J	a->1	
art.K	o->2	
art.M	e->1	
art.S	t->1	
art.V	a->1	i->2	
art.Ä	v->1	
art: 	e->1	
arta 	e->1	f->1	k->1	o->2	p->1	ä->1	
artad	 ->1	e->2	
artan	n->3	
artar	.->2	
artas	 ->2	
artat	s->2	
artec	k->4	
artel	l->15	
artem	e->9	
arten	 ->7	d->1	
arter	 ->10	,->2	.->3	n->10	
artex	t->3	
arthy	 ->1	
arti 	a->1	d->1	f->2	h->2	i->4	k->1	m->1	p->1	s->7	t->2	å->1	
arti,	 ->7	
arti.	.->1	D->1	H->1	K->1	
artid	 ->2	
artie	l->2	r->10	t->30	
artif	i->2	
artig	h->1	
artii	n->1	
artik	e->93	l->14	r->1	
artil	e->1	
artin	e->1	
artip	r->2	
artis	 ->1	k->3	p->1	
artlä	g->1	
artne	r->28	
arton	h->1	
artpl	a->1	
artra	n->1	r->1	
artsi	n->1	
artsm	e->1	y->1	
artso	r->2	
artss	e->3	
artyg	 ->28	)->1	,->3	.->4	;->1	e->20	s->12	
arv o	c->1	
arv, 	a->1	e->1	s->1	
arv."	D->1	
arv.B	a->1	
arv.E	n->1	
arvat	t->9	
arven	.->1	
arver	 ->1	
arvet	 ->3	,->1	
arvid	 ->3	
arvli	g->1	
arvsi	n->1	
arvss	t->2	
arvär	l->1	
ary o	c->1	
arzwa	l->1	
arämb	e->1	
aråda	n->1	
aråde	t->1	
arébe	t->1	
arón 	C->2	
as - 	o->2	
as 40	0->1	
as Eu	r->8	
as Sj	ö->2	
as ag	e->1	
as al	l->1	
as an	d->2	g->1	m->1	s->23	t->2	
as ar	b->6	
as at	t->72	
as au	t->1	
as av	 ->102	g->1	s->1	t->1	
as ax	l->1	
as be	f->1	h->1	r->1	s->3	t->5	
as bi	d->1	
as bl	a->3	i->2	
as bo	r->5	
as br	i->1	
as bä	r->1	s->1	t->1	
as bö	r->1	
as ce	n->5	
as da	 ->5	g->1	
as de	 ->4	l->4	m->3	n->5	r->1	t->6	
as di	p->1	r->2	s->1	
as dj	u->1	
as du	b->1	
as dä	r->7	
as dö	d->1	
as ef	f->1	t->8	
as eg	e->1	n->3	
as ek	o->6	
as el	l->9	
as en	 ->20	d->3	h->3	l->1	s->1	
as et	t->9	
as ev	e->1	
as ex	a->1	e->2	
as fa	b->1	k->1	r->1	v->1	
as fi	s->1	
as fl	a->1	e->1	
as fo	l->2	r->1	
as fr	a->7	i->2	å->14	
as fu	l->4	n->2	
as få	 ->3	
as fö	l->1	r->73	
as ga	n->1	r->1	
as ge	m->3	n->14	o->1	
as gr	u->1	
as gu	v->1	
as ha	n->1	r->2	v->3	
as hi	s->1	
as hj	ä->2	
as hu	v->2	
as hy	c->1	
as hä	l->1	n->1	r->3	
as hå	r->3	
as i 	B->1	E->4	K->1	M->2	S->2	U->1	b->3	d->21	e->5	f->12	g->1	h->4	k->4	l->1	m->1	n->1	o->1	p->7	r->6	s->8	t->3	v->2	Ö->1	ö->1	
as id	e->1	
as ig	e->1	
as in	 ->4	,->2	b->1	d->2	f->1	g->1	k->1	l->2	n->1	o->8	s->2	t->23	
as ir	r->1	
as ja	g->10	
as ju	r->3	s->1	
as jä	m->1	
as ka	b->1	l->2	p->2	t->1	
as kl	a->2	
as ko	m->13	n->8	p->1	r->3	
as kr	a->3	
as ku	l->1	m->1	s->1	
as kv	a->3	
as kä	n->1	
as kö	p->1	
as la	g->4	n->1	
as le	 ->1	d->1	g->4	v->3	
as li	k->3	t->1	v->2	
as lä	m->1	n->1	
as ma	k->1	n->1	s->1	
as me	d->58	l->2	r->3	
as mi	l->2	
as mo	t->4	
as my	c->5	
as mä	r->1	
as må	l->1	s->2	
as mö	j->4	t->1	
as na	c->1	m->2	t->9	
as ne	d->1	
as ni	 ->1	o->1	v->1	
as no	r->1	
as nu	 ->3	v->1	
as nä	r->9	
as nå	g->9	
as ob	l->1	
as oc	h->59	k->6	
as of	f->3	t->2	ö->2	
as oh	j->1	
as oi	n->2	
as ol	a->1	i->2	j->1	y->1	
as om	 ->17	.->1	
as or	d->3	g->1	o->2	
as ov	a->1	
as pa	r->3	
as pe	n->1	r->1	
as pl	a->2	
as po	l->5	t->1	
as pr	o->6	
as på	 ->58	,->1	
as ra	d->1	t->1	
as re	a->1	f->1	g->4	s->1	
as ri	g->1	
as ro	l->2	
as ru	n->3	
as rä	d->1	k->1	t->12	
as rö	s->1	t->1	
as sa	d->1	k->3	m->9	
as se	d->1	k->1	n->1	
as si	d->4	t->1	
as sj	ä->2	
as sk	a->7	e->1	i->1	o->1	r->1	u->2	y->1	
as sl	a->1	u->1	
as sn	a->3	
as so	c->4	m->23	
as sp	e->3	
as st	a->1	r->2	u->1	ä->2	å->2	ö->3	
as su	b->1	v->3	
as sv	a->1	å->2	
as sy	n->1	
as sä	k->4	l->1	r->1	t->1	
as så	 ->9	
as sö	n->2	
as ta	 ->1	l->1	n->1	
as ti	l->50	o->1	
as tj	ä->1	
as tr	a->1	o->3	
as tu	l->1	r->1	
as tv	ä->1	å->1	
as ty	d->2	v->1	
as un	d->19	
as up	p->22	
as ur	 ->1	
as ut	 ->4	,->1	.->1	a->5	f->1	g->1	t->2	v->2	
as va	c->1	l->1	r->10	t->1	
as ve	c->1	r->9	
as vi	 ->4	a->1	d->8	k->2	
as vä	g->4	l->1	r->3	s->1	
as vå	r->2	
as yr	k->1	
as yt	t->3	
as äg	a->2	
as än	 ->1	d->2	
as är	 ->6	
as äv	e->2	
as ål	d->2	
as år	l->2	
as ås	t->1	
as åt	 ->3	a->1	m->1	
as öd	e->1	
as ög	o->1	
as öm	s->1	
as ön	s->1	
as öp	p->1	
as ör	o->1	
as öv	e->8	
as!De	t->1	
as!Eu	r->1	
as!Ge	n->1	
as!He	r->1	
as".J	a->1	
as, M	i->1	
as, a	n->1	t->4	
as, b	e->1	ä->1	
as, d	å->1	
as, e	f->4	n->3	t->2	
as, f	r->2	ö->6	
as, g	e->1	
as, h	a->1	e->1	u->1	ä->1	
as, i	 ->4	n->2	
as, k	o->1	
as, l	e->1	
as, m	e->6	ä->1	
as, n	ä->1	
as, o	c->11	m->3	
as, p	å->2	
as, r	e->1	
as, s	a->1	k->1	o->2	p->2	ä->2	å->6	
as, u	r->1	t->6	
as, v	a->1	i->2	
as, ä	v->1	
as, å	t->1	
as. D	e->2	
as. M	e->1	
as. P	a->1	
as.- 	(->1	
as.Al	l->1	
as.At	t->1	
as.Be	t->1	v->1	
as.Bl	a->2	
as.Ce	n->1	
as.De	 ->2	n->5	t->18	
as.Dä	r->5	
as.Då	 ->1	
as.Ek	o->1	
as.En	l->1	
as.Et	t->3	
as.Fl	o->1	
as.Fr	u->2	å->1	
as.Fö	r->2	
as.Ge	n->2	
as.Gr	e->1	
as.He	l->1	r->5	
as.Hi	s->1	t->1	
as.I 	a->2	d->1	e->1	l->1	r->1	s->1	ö->1	
as.In	g->1	o->1	
as.Ja	g->8	
as.Jo	n->1	
as.Jä	m->1	
as.Ko	m->4	
as.Ma	n->1	
as.Me	d->3	n->4	
as.Mi	n->1	
as.Ni	 ->1	
as.Nä	r->2	
as.Om	 ->1	
as.Pa	r->3	
as.Pe	r->1	
as.Pr	e->1	o->1	
as.På	 ->1	
as.Re	s->1	
as.Sa	m->1	
as.Sl	u->1	
as.Sn	a->1	
as.Ta	l->1	
as.Ti	l->1	
as.Un	d->1	
as.Va	d->3	
as.Vi	 ->15	d->1	
as.Vå	r->1	
as.Yt	t->1	
as.Än	d->1	
as.Åt	a->1	g->1	
as: a	n->1	
as: e	n->1	
as; e	n->1	
as?Ha	r->1	
as?Sk	u->1	
asabl	a->1	
asaca	 ->1	
asade	 ->2	
asar!	D->1	
asar,	 ->1	
asas 	s->1	
asat 	o->1	
asatt	e->1	
asbou	r->5	
asche	n->2	r->1	
aschh	o->1	
ascis	m->3	t->9	
ase.O	m->1	
aseba	l->1	
asen 	"->1	i->5	k->1	
asen,	 ->1	
asen.	P->1	
aser 	f->1	o->1	
aser,	 ->1	
aser.	 ->1	
asera	d->4	r->2	s->2	
asern	a->2	
ashat	e->1	
ashin	g->3	
ashus	.->1	
asiat	i->2	
asien	 ->3	.->1	s->1	
asifu	l->1	
asili	e->1	
asin 	s->1	
asis 	a->2	o->1	
asis,	 ->1	
asism	 ->6	,->2	.->4	e->3	
asist	.->1	i->11	
ask f	o->1	
askad	 ->1	e->1	
askam	m->1	
askar	,->1	
asker	a->2	
askie	n->2	
askin	 ->3	e->3	
askis	k->4	
askra	r->1	
askus	 ->1	
asm f	ö->1	
asm p	å->1	
asm s	o->1	
asmat	t->1	
asmug	g->1	
asnin	g->3	
asoch	i->1	
asor,	 ->1	
aspek	t->34	u->2	
aspis	k->1	
ass e	l->1	
ass f	å->1	ö->1	
ass o	m->1	
ass t	j->1	
ass v	i->1	
assa 	d->1	h->1	o->1	p->2	r->1	v->1	
assad	 ->3	ö->1	
assag	e->1	
assak	r->1	
assan	d->2	
assar	 ->1	b->2	
assas	 ->6	
assav	g->1	
asse-	N->1	
assen	s->2	
asser	 ->1	a->3	i->1	n->1	
assif	i->9	
assig	t->1	
assio	n->2	
assis	k->5	t->2	
assiv	 ->1	.->1	a->1	t->1	
assla	t->1	
assme	d->3	
assni	n->4	
assoc	i->1	
asson	i->1	
assor	 ->1	,->1	
asspe	l->1	
asst 	m->1	
assus	e->1	
ast 1	 ->1	
ast 2	5->1	
ast 5	,->1	
ast 7	0->1	
ast 9	 ->1	
ast a	c->1	l->1	n->2	t->5	v->1	
ast b	e->2	
ast d	e->5	r->1	
ast e	n->6	r->1	t->5	
ast f	a->3	r->1	u->1	å->1	ö->5	
ast g	e->1	l->1	ä->1	å->1	ö->1	
ast h	a->2	
ast i	 ->10	n->3	
ast k	a->4	o->2	r->1	u->3	
ast l	ä->1	ö->1	
ast m	e->4	i->1	o->1	å->2	ö->3	
ast n	e->1	i->1	y->1	ä->2	å->1	
ast o	b->1	m->4	p->1	r->1	
ast p	e->1	r->1	å->3	
ast r	u->1	ä->1	ö->1	
ast s	a->1	o->2	y->1	å->2	
ast t	a->1	i->11	r->1	v->2	ä->1	
ast u	p->1	t->4	
ast v	a->1	i->11	ä->1	
ast ä	r->7	
ast å	r->1	t->3	
ast ö	v->2	
ast!D	ä->1	
ast, 	P->1	d->1	m->1	s->1	v->1	
ast- 	o->1	
ast.D	e->1	
ast.E	f->1	
ast.K	ä->1	
ast.N	u->1	
ast.V	i->1	
ast?V	i->1	
asta 	d->5	g->1	i->1	n->1	o->1	s->3	
astad	 ->1	.->2	e->1	
astan	d->2	
astar	 ->4	e->1	
astas	 ->1	,->1	t->1	
astat	 ->2	.->1	s->2	
aste 	-->1	E->2	a->5	b->3	c->1	d->10	e->6	f->12	g->2	h->2	i->3	j->1	k->6	l->1	m->16	n->1	o->3	p->4	r->10	s->13	t->15	u->5	v->6	ä->2	å->16	
aste,	 ->1	
aste.	D->1	F->1	V->1	
aste:	 ->1	
asten	 ->3	,->1	.->1	s->1	
aster	,->1	a->1	
astet	 ->1	.->3	
astia	n->1	
astig	a->1	h->1	
astin	d->1	
astio	n->1	
astis	k->12	
astku	b->1	
astla	g->1	n->2	
astlä	g->2	
astna	r->1	
astni	n->7	
astod	o->1	
astri	c->6	
astro	f->90	n->1	
astru	k->15	
astsl	a->2	o->2	å->17	
astst	ä->51	
astu 	m->1	
astän	 ->1	
aståe	n->2	
asune	r->1	
asus 	k->2	o->1	
asyl 	g->1	o->3	
asyl,	 ->2	
asyl-	 ->1	
asyl.	D->1	J->1	V->1	
asylb	e->1	
asylf	ö->2	
asylr	ä->2	
asyls	ö->6	
asäke	r->1	
asätt	a->13	e->3	s->3	
aså e	n->1	
aså h	a->1	
aså s	a->1	
aså v	i->1	
at "K	v->1	
at "e	k->1	
at - 	a->1	d->1	f->2	i->1	j->2	k->1	s->1	å->1	
at -,	 ->1	
at 39	 ->1	
at 90	 ->1	
at Ad	o->1	
at Br	o->1	
at Er	i->1	
at Eu	r->5	
at Fl	o->1	
at Fr	a->1	
at It	a->1	
at Ki	r->1	
at Sj	ö->1	
at ad	m->1	
at al	l->5	
at an	d->1	g->2	s->4	t->1	
at ar	b->1	t->1	
at at	t->41	
at av	 ->12	s->2	
at ba	k->1	
at be	g->2	h->2	k->1	r->1	s->1	t->6	
at bi	l->2	
at bl	i->1	
at bo	r->1	
at br	e->1	
at bö	r->1	
at de	 ->8	l->1	m->3	n->7	t->13	
at di	r->4	
at do	k->1	
at dr	a->2	
at dä	r->2	
at dö	d->1	
at ef	t->2	
at em	o->3	
at en	 ->21	a->1	o->1	
at er	 ->2	a->1	t->1	
at et	t->12	
at ex	t->1	
at fa	l->6	s->1	
at fi	n->1	s->2	
at fl	e->2	
at fo	l->1	r->1	
at fr	a->3	i->2	å->7	
at få	 ->1	.->1	g->2	r->2	
at fö	r->38	
at ge	n->5	
at gr	a->1	
at gå	 ->1	
at gö	r->5	
at ha	 ->2	d->1	n->2	r->6	
at he	m->1	
at hi	n->1	t->1	
at ho	n->1	s->1	t->1	
at hu	r->3	
at hä	r->2	
at hå	l->2	
at hö	g->2	r->1	
at i 	D->1	I->1	K->1	M->1	a->2	b->1	d->2	e->2	f->4	g->1	k->1	o->1	p->1	r->2	s->2	u->2	Ö->1	ä->1	
at ic	k->2	
at if	r->1	
at ig	e->2	
at in	 ->2	f->1	n->1	o->3	t->4	v->1	
at ja	g->1	
at ju	s->1	
at kl	a->1	
at ko	a->1	l->1	m->4	n->11	
at kr	a->1	
at kö	t->1	
at la	g->1	n->2	
at le	v->1	
at li	v->2	
at lä	g->2	m->1	n->1	
at lå	n->1	
at ma	n->1	r->1	
at me	d->11	n->1	
at mi	g->4	l->1	
at mo	d->1	t->6	
at my	c->4	
at mä	n->1	
at må	n->1	s->4	
at ne	d->1	
at nu	.->1	
at nä	r->2	
at nå	g->6	
at nö	j->1	
at oc	h->23	k->2	
at ol	y->1	
at om	 ->14	,->1	.->2	r->2	
at or	d->2	
at os	s->9	
at pa	r->1	
at pr	i->1	o->7	
at på	 ->18	,->1	b->1	p->1	
at re	s->2	
at rä	t->2	
at rå	d->2	
at rö	s->2	
at sa	m->2	
at se	n->1	
at si	g->26	n->4	t->4	
at sj	u->2	
at sk	a->2	o->1	r->1	
at so	m->21	
at st	ä->1	ö->8	
at sy	f->1	s->1	
at sä	k->2	n->1	t->8	
at så	 ->7	d->1	
at sö	k->1	
at ta	 ->2	g->1	l->1	r->1	
at ti	d->1	l->17	
at tr	a->1	u->1	
at tä	m->1	
at un	d->7	
at up	p->6	
at ur	a->6	
at ut	 ->2	,->1	b->2	f->1	p->1	s->1	t->1	
at va	d->2	l->1	r->2	t->1	
at vi	 ->1	a->2	k->1	l->2	s->4	
at vä	g->1	l->1	n->1	
at vå	r->3	
at yt	t->1	
at äm	n->1	
at än	 ->12	d->2	
at är	 ->1	
at år	,->1	.->2	
at åt	g->1	n->1	
at ök	a->1	
at öv	e->1	
at, a	t->2	
at, b	e->1	y->1	
at, d	ä->1	
at, e	f->3	l->1	n->2	
at, f	ö->1	
at, h	a->2	
at, i	 ->2	n->1	
at, k	o->2	r->1	
at, l	å->1	
at, m	e->4	
at, n	ä->2	
at, o	c->10	m->2	
at, p	r->1	å->1	
at, s	j->1	o->3	å->1	
at, u	t->3	
at, v	i->3	
at, ä	n->1	r->2	
at. F	r->1	
at. H	e->1	ä->1	
at. O	f->1	
at..H	e->1	
at.Be	r->1	
at.Bi	l->1	
at.De	 ->2	s->2	t->15	
at.Dä	r->3	
at.En	d->1	l->2	
at.FP	Ö->1	
at.Fö	r->2	
at.Ge	n->1	
at.Gr	u->1	
at.He	r->5	
at.Hu	r->2	
at.Hä	r->1	
at.I 	d->3	f->1	s->1	
at.Ja	g->10	
at.Ko	m->2	n->1	
at.Ku	l->1	
at.Lä	n->1	
at.Me	d->1	
at.Ni	 ->1	
at.Oc	h->1	
at.Om	 ->1	
at.Pr	o->1	
at.Ta	c->1	
at.Ti	l->1	
at.Tr	o->1	
at.Va	d->2	r->1	
at.Vi	 ->1	
at.Än	d->1	
at.Å 	a->1	
at.Öv	r->1	
at: "	a->1	
at: h	a->1	
at: j	a->1	
at; a	l->1	
at?.(	E->1	
at?Jo	 ->1	
ata a	k->1	
ata f	ö->6	
ata i	n->1	
ata k	ä->1	
ata m	e->1	o->1	
ata o	c->4	m->3	r->1	
ata s	e->4	
ata å	t->1	
ata, 	u->1	
ataba	s->1	
atal 	h->1	
atalo	g->2	
atals	 ->4	s->1	
ataly	s->2	
atane	n->3	
atar 	o->1	
atast	r->89	
atasä	k->1	
atcha	n->1	
atche	r->1	
ate c	o->2	
ategi	 ->17	,->3	.->3	e->14	n->8	p->1	s->17	
atego	r->8	
ateko	n->1	
atell	i->3	
atema	l->1	t->1	
aten 	-->1	B->1	a->7	b->1	e->1	f->4	g->1	h->1	k->1	m->3	o->2	s->2	t->1	u->1	
aten,	 ->7	
aten.	D->3	M->2	O->1	V->1	
atens	 ->5	
ater 	-->4	a->2	b->1	d->3	e->3	f->11	g->1	h->4	i->7	k->1	m->6	o->7	p->2	s->13	t->3	u->5	v->4	ö->1	
ater)	 ->2	
ater,	 ->10	
ater-	n->1	
ater.	B->1	D->3	J->3	K->1	L->1	M->2	O->1	S->2	U->1	V->2	Ä->1	
ater;	 ->1	
ater?	B->1	
atera	 ->28	,->1	.->1	d->6	l->8	n->2	r->5	s->1	t->3	
aterg	r->1	
ateri	a->23	e->4	n->1	
atern	a->219	
aters	 ->3	
ates-	 ->1	
atet 	a->17	b->1	f->12	i->1	k->2	m->2	o->4	s->2	ä->4	
atet,	 ->4	
atet.	.->1	D->1	H->1	J->1	V->1	
ateti	s->1	
atför	ä->4	
ath h	a->1	
ath n	ä->1	
ath o	c->1	
ath, 	o->1	
athie	s->2	
ati d	e->1	
ati f	ö->3	
ati i	n->1	
ati k	r->1	
ati m	e->1	
ati o	c->9	
ati s	o->1	
ati u	p->1	
ati" 	s->1	
ati, 	b->1	e->1	o->1	s->1	
ati.D	e->2	
ati.E	f->1	n->1	
ati.F	o->1	
ati.H	e->1	
ati.I	 ->1	
ati.K	u->1	
ati.M	i->1	
atien	t->4	
atier	 ->1	n->3	
atifi	c->13	
atifr	å->1	
atik,	 ->1	
atike	n->4	
atin 	a->1	b->1	h->1	i->1	o->3	s->3	v->1	
atin,	 ->1	
atin.	F->2	H->1	O->1	
atino	s->4	
atinr	i->1	
atins	 ->4	
ation	 ->139	,->14	.->30	:->3	?->3	a->41	e->454	s->38	
atire	f->1	
atis 	e->1	i->1	t->1	å->1	
atise	r->5	
atisk	 ->30	a->71	t->33	
atist	i->9	
ativ 	-->2	E->1	a->2	d->1	f->10	g->1	h->1	i->5	k->2	l->2	m->2	o->4	p->3	r->1	s->20	t->8	v->1	ä->2	
ativ,	 ->7	
ativ.	 ->1	.->1	B->1	D->1	E->1	M->1	R->1	S->1	Y->1	
ativ;	 ->1	
ativa	 ->46	,->2	.->1	n->1	
ativb	e->1	
ative	n->2	t->14	
ativf	ö->1	
ativi	s->1	t->1	
ativr	i->1	ä->4	
ativt	 ->22	,->2	.->2	
atjän	s->1	
atlan	d->1	t->2	
atlig	 ->8	a->67	h->2	t->23	
atlis	t->2	
atlän	d->10	
atnyt	t->1	
ato -	 ->1	
ato f	ö->2	
ato h	a->1	
ato i	 ->1	
ato o	m->1	
ato s	a->1	å->1	
ato t	i->1	
ato ö	p->1	
ato.J	a->1	
atoak	t->1	
atoba	s->1	
atobe	t->1	
atoge	n->2	
atoli	k->4	
atols	k->3	
atom 	o->3	
atom)	 ->1	
atome	n->3	
atomf	o->1	
aton-	H->1	
atons	 ->1	
ator 	f->1	
ator,	 ->1	
atorb	r->1	
atore	r->6	
atori	e->1	s->15	u->2	
atorl	ä->1	
atorn	 ->1	a->1	
ators	k->1	
atos 	b->9	e->1	f->1	o->1	v->1	
atpen	s->1	
atper	i->9	
atpro	t->1	
atrio	t->1	
ats -	 ->5	
ats E	u->1	
ats S	p->2	
ats a	v->32	
ats b	o->1	
ats d	e->2	ä->2	
ats e	l->1	n->2	r->1	x->1	
ats f	l->1	o->1	r->2	å->3	ö->15	
ats g	e->3	o->1	ö->2	
ats h	a->1	i->1	o->2	å->1	
ats i	 ->24	n->5	
ats k	o->1	
ats l	e->1	
ats m	e->7	i->1	o->2	å->1	
ats n	e->1	ä->1	
ats o	c->8	m->2	
ats p	r->1	å->9	
ats r	e->2	ä->1	
ats s	e->1	o->4	t->1	u->1	
ats t	i->24	
ats u	n->4	p->2	t->6	
ats v	a->2	i->4	
ats ä	n->1	r->1	
ats å	t->2	
ats, 	a->2	d->2	e->3	h->1	m->4	n->2	o->4	p->1	s->3	t->1	v->4	å->1	
ats- 	o->5	
ats.D	e->10	ä->1	å->1	
ats.E	n->2	r->1	
ats.F	a->1	
ats.H	e->1	o->1	
ats.J	a->2	
ats.K	o->2	
ats.M	e->1	
ats.R	e->1	
ats.S	å->1	
ats.V	i->1	
ats.Ä	n->1	
ats?F	r->1	
ats?K	o->1	
atsa 	a->1	m->1	p->4	s->1	
atsar	 ->3	
atsas	 ->2	
atsat	s->1	
atsba	n->2	
atsen	 ->19	!->1	,->1	.->3	;->1	
atser	 ->44	,->7	.->8	n->20	
atsfö	r->1	
atska	p->1	
atsma	k->2	
atsmi	n->2	
atsni	n->4	v->4	
atsos	 ->2	,->1	
atspr	i->1	
atsst	y->3	ö->19	
att "	P->1	
att -	 ->8	
att 1	9->3	
att 2	5->1	
att 4	0->1	
att 7	0->1	
att 8	0->1	
att A	l->1	m->2	
att B	a->3	o->1	r->1	
att C	E->1	
att D	a->3	
att E	G->9	I->1	K->1	L->1	U->12	r->1	u->64	v->1	
att F	E->1	N->1	P->1	l->1	ö->1	
att G	r->1	
att I	C->1	r->1	s->3	t->1	
att J	ö->3	
att K	o->2	
att M	a->2	
att N	a->1	
att O	L->3	
att P	a->1	o->2	
att R	I->1	a->1	o->1	
att S	a->1	o->1	t->1	
att T	h->2	o->1	u->13	
att V	ä->1	
att a	c->5	d->1	g->13	k->4	l->39	m->1	n->68	r->40	v->39	
att b	a->6	e->158	i->31	l->48	o->5	r->18	u->2	y->14	ä->1	å->4	ö->22	
att c	i->1	
att d	a->7	e->978	i->37	o->5	r->24	u->1	y->2	ä->8	ö->9	
att e	f->10	k->2	l->3	n->85	p->1	r->13	t->25	u->2	v->1	x->6	
att f	a->21	e->1	i->17	l->5	o->29	r->57	u->13	y->2	å->88	ö->241	
att g	a->18	e->106	i->1	l->2	o->11	r->20	y->4	ä->5	å->25	ö->106	
att h	a->96	e->6	i->7	j->14	o->8	u->2	y->1	ä->11	å->19	ö->9	
att i	 ->39	a->1	b->2	d->6	f->5	g->1	m->2	n->145	r->1	s->2	
att j	a->84	o->3	u->3	ä->1	
att k	a->5	l->11	n->4	o->207	r->24	u->57	v->5	ä->3	ö->2	
att l	a->15	e->20	i->14	o->2	u->3	y->13	ä->53	å->10	ö->18	
att m	a->220	e->38	i->37	o->14	u->1	y->16	ä->10	å->8	ö->8	
att n	a->2	e->1	i->45	o->6	u->2	y->3	ä->20	å->22	ö->1	
att o	c->18	f->6	k->2	l->4	m->43	n->1	p->1	r->13	s->2	
att p	a->34	e->13	l->6	o->6	r->37	u->1	å->47	
att r	a->6	e->61	i->11	o->2	u->1	ä->15	å->24	ö->32	
att s	a->35	e->57	i->7	j->6	k->125	l->12	m->1	n->6	o->13	p->13	t->104	u->2	v->6	y->6	ä->64	å->14	ö->3	
att t	.->1	a->102	e->1	h->1	i->96	j->3	o->6	r->7	u->3	v->8	y->4	ä->12	å->1	
att u	n->62	p->73	r->4	t->121	
att v	a->71	e->15	i->441	ä->26	å->20	
att y	t->6	
att z	o->1	
att ä	g->21	n->21	r->5	v->19	
att å	 ->3	k->1	r->3	s->6	t->41	
att ö	k->20	n->2	p->4	s->1	v->42	
att, 	E->1	d->1	e->3	f->2	g->1	i->2	l->1	o->3	s->3	t->1	u->1	v->1	ä->1	å->1	
att..	.->1	
att.D	e->6	ä->1	
att.F	ö->2	
att.H	e->2	
att.J	a->1	
att.K	o->1	
att.L	å->2	
att.M	e->3	
att.N	i->1	
att.P	P->1	a->1	
att.T	a->1	
att.U	t->1	
att.V	i->2	
att: 	"->1	o->1	
att?V	i->1	
attBe	t->1	
atta 	a->2	b->10	d->8	e->5	f->3	g->2	i->5	k->1	m->7	n->1	o->7	p->1	r->2	s->4	t->2	u->3	v->4	å->1	
atta.	J->1	P->1	S->1	V->1	
attac	k->2	
attad	 ->1	e->10	
attan	 ->1	d->40	t->1	
attar	 ->40	.->1	e->4	n->4	
attas	 ->29	.->1	
attat	 ->9	s->9	
attav	l->7	
atte 	i->2	j->1	
atte-	 ->1	
atteb	a->1	e->14	
attef	r->2	ö->1	
attei	n->2	
attel	ä->1	
atten	 ->68	!->2	,->16	.->17	;->1	?->1	F->1	d->2	f->2	p->1	r->2	s->3	t->5	v->8	
attep	o->1	
atter	 ->8	,->1	.->1	a->13	n->1	
attes	 ->4	.->2	a->1	y->1	
attig	a->18	d->12	
attin	n->1	
attit	y->5	
attkv	ä->1	
attle	 ->3	.->1	
attna	 ->1	r->2	s->3	
attne	n->2	t->6	
attni	n->68	
attra	k->1	
attre	t->1	
atts 	a->1	f->1	
atts.	N->1	
atuer	a->2	
atula	t->6	
atule	r->31	
atum 	d->1	f->2	o->1	s->4	å->1	
atum,	 ->2	
atum.	I->1	
atume	t->2	
atur 	-->1	e->1	o->3	
atur,	 ->3	
atur-	 ->1	
atur.	D->2	V->1	
atura	.->1	
ature	n->14	r->4	
aturf	ö->2	
aturk	-->1	a->13	
aturl	i->102	
aturn	ö->1	
aturo	m->1	
aturv	e->1	
atus 	a->1	e->1	q->2	
atus.	D->1	
atus?	O->1	
atuse	n->4	
atusf	ö->1	
atzid	a->2	
atäck	n->1	
atöre	n->1	r->3	
atöve	r->6	
atürk	d->1	
au du	 ->1	
au fö	r->4	
au oc	h->1	
au sa	 ->1	d->2	
au", 	d->1	
au, L	a->1	
au, a	n->1	
au, e	f->1	
au, h	a->1	
au, o	c->1	
au, s	o->2	
au.Et	t->1	
auMed	 ->1	
aubet	ä->1	
aucto	r->1	
aude 	M->1	
audro	n->1	
auen,	 ->1	
auer 	s->1	
auern	t->1	
aufma	n->1	
aukas	u->3	
aukto	r->6	
aumat	i->1	
auna 	ä->1	
aunio	n->3	
aurer	i->1	
auro,	 ->1	
aus b	e->3	
ausse	n->1	
ausul	 ->2	.->1	e->3	
autom	a->8	
autop	i->1	
autre	 ->1	s->1	
aux, 	n->1	
av "p	a->1	
av "r	e->1	i->1	
av - 	d->1	i->1	o->2	s->1	u->1	
av 14	 ->1	
av 19	 ->1	9->2	
av 20	0->1	
av 40	 ->1	
av 5 	0->1	
av 54	0->1	
av 8 	4->1	
av Ah	e->2	
av Am	e->1	s->1	
av Ar	a->1	
av BN	I->1	P->5	
av BS	E->1	
av Ba	r->2	
av Be	r->8	
av Bo	u->1	
av Br	o->2	
av Ca	n->1	
av Da	 ->1	v->1	
av De	m->1	
av Di	m->2	
av Du	b->1	
av Dü	h->1	
av EG	-->1	
av EU	 ->3	,->1	-->4	.->2	:->7	
av Er	i->1	
av Eu	r->70	
av Ex	x->2	
av FN	:->1	
av FP	Ö->2	
av Fl	o->1	
av Fö	r->8	
av Ga	z->1	
av Ge	n->2	
av Gr	a->2	o->1	
av Ha	i->1	
av He	n->1	
av Hi	t->1	
av Is	r->2	
av Ja	c->1	
av Je	r->1	
av Jo	n->2	
av Ki	n->3	
av Ko	c->3	s->7	
av Ku	l->1	
av La	n->3	
av Li	b->1	
av Lö	ö->1	
av Ma	r->2	
av Mc	N->1	
av Mo	r->1	
av OL	A->3	
av Os	m->1	
av Oz	 ->1	
av Pa	l->1	t->1	
av Po	r->1	
av Pé	t->1	
av Ra	p->1	
av Ri	i->1	
av Sa	m->1	
av Sc	h->6	
av Ta	c->1	
av Te	r->1	
av Th	e->3	y->1	
av Ti	b->1	
av To	t->1	
av UN	M->1	
av Va	n->1	r->1	
av Vä	s->1	
av Wa	l->1	
av Wi	e->1	
av Wy	e->1	
av ac	c->1	
av ad	m->1	v->1	
av ag	e->1	
av al	b->1	d->1	k->1	l->29	
av an	b->1	d->3	l->2	m->1	o->1	s->14	t->3	v->1	
av ap	r->2	
av ar	b->19	t->20	
av as	y->1	
av at	t->64	
av av	 ->1	f->1	g->3	p->1	t->2	v->1	
av ba	r->2	
av be	d->1	f->6	g->1	h->5	k->1	s->14	t->8	v->2	
av bi	d->2	l->11	o->1	
av bl	a->1	y->1	å->1	
av bo	l->1	m->2	
av br	e->1	i->4	o->4	u->1	
av bu	d->8	
av by	g->2	
av bå	d->2	
av bö	c->1	r->2	
av ce	n->2	
av ci	r->2	v->4	
av co	m->1	
av da	g->4	t->1	
av de	 ->164	b->3	f->1	l->3	m->26	n->172	r->6	s->45	t->124	
av di	p->1	r->20	s->4	v->1	
av dj	u->1	
av do	k->1	m->11	
av dr	i->1	
av ef	f->2	t->2	
av eg	e->2	
av ek	o->10	
av en	 ->98	b->1	e->5	h->1	i->1	o->1	t->2	
av er	 ->9	,->2	:->1	a->3	f->1	t->2	
av et	n->1	t->51	
av eu	r->7	
av ev	e->1	
av ex	a->6	p->1	t->1	
av fa	k->3	l->2	r->39	t->3	
av fi	n->3	s->3	
av fj	o->2	
av fl	e->9	o->1	y->6	
av fo	l->1	n->1	r->6	
av fr	a->1	e->1	i->11	ä->5	å->10	
av fu	l->2	n->1	s->2	
av fy	s->1	
av fä	d->1	
av få	 ->1	n->1	
av fö	l->2	r->105	
av ga	m->3	
av ge	m->28	n->2	o->1	
av gi	f->1	g->1	v->1	
av gl	o->1	
av go	d->1	
av gr	a->2	o->1	u->3	ä->4	ö->1	
av gö	r->1	
av ha	n->4	r->1	t->2	v->4	
av he	l->6	m->1	
av hi	e->1	g->1	s->3	
av ho	n->1	
av hu	n->1	r->7	
av hä	n->1	r->1	
av hö	g->2	
av i 	d->4	s->1	
av ib	e->1	
av ic	k->3	
av id	e->1	é->1	
av im	p->4	
av in	d->1	e->1	f->4	i->2	n->3	o->1	s->5	t->8	v->1	
av jo	r->5	
av ju	r->1	s->3	
av jä	m->2	
av ka	m->2	n->3	p->1	r->2	t->2	
av kl	a->4	
av kn	u->1	
av ko	a->2	l->4	m->57	n->38	r->2	s->6	
av kr	i->4	ä->1	
av ku	l->4	s->1	
av kv	i->4	o->1	
av kä	r->8	
av la	g->10	n->8	s->1	
av le	d->9	g->1	j->1	
av li	b->2	c->1	k->2	v->8	
av lo	j->2	k->3	
av lä	g->1	n->2	t->1	
av lå	n->1	
av lö	v->1	
av ma	k->2	n->2	r->10	t->4	
av me	d->23	r->3	
av mi	g->2	l->13	n->17	s->3	t->3	
av mo	d->2	n->1	t->2	
av my	c->3	
av mä	n->7	
av må	l->3	n->4	
av mö	j->1	
av na	t->13	z->1	
av ni	 ->1	
av no	r->1	
av ny	 ->2	a->6	b->1	h->1	n->1	
av nä	r->1	s->1	
av nå	g->6	
av nö	d->2	
av oa	c->1	n->1	
av ob	e->2	
av oc	h->7	
av of	f->4	r->1	
av ok	l->1	
av ol	i->8	j->3	y->3	
av om	 ->4	b->1	k->1	r->2	s->2	
av on	d->1	
av or	d->7	i->1	k->1	s->2	
av os	s->12	
av ot	r->1	v->1	
av ou	n->1	
av ov	a->1	
av pa	k->1	l->1	r->20	
av pe	n->7	r->5	
av pi	o->1	
av po	l->8	
av pr	e->1	i->8	o->28	
av på	 ->17	
av ra	m->2	p->3	s->1	
av re	f->2	g->17	k->1	n->1	p->1	s->8	t->1	v->1	
av ri	k->4	s->3	
av ry	s->1	
av rä	d->1	k->5	t->6	
av rå	d->12	
av rö	s->1	
av sa	m->12	
av sc	e->1	
av se	k->2	n->1	r->1	s->2	x->1	
av si	g->3	n->13	s->1	t->7	
av sj	u->1	ä->1	ö->1	
av sk	a->8	e->1	o->4	r->3	ä->3	ö->1	
av sl	u->2	
av sm	å->2	
av so	c->7	m->8	
av sp	e->1	l->1	
av st	a->19	i->1	o->14	r->14	y->1	ä->1	å->2	ö->20	
av su	b->3	c->1	
av sv	a->1	ä->1	
av sy	n->1	s->19	
av sä	k->9	r->5	
av så	 ->3	d->7	
av ta	l->2	
av te	k->4	l->1	r->3	
av ti	d->2	l->11	
av tj	ä->28	
av to	t->2	
av tr	a->7	e->2	y->1	ä->1	
av tu	n->5	r->1	
av tv	å->1	
av ty	d->1	p->1	
av tä	n->1	
av un	d->6	g->2	i->19	
av up	p->6	
av ut	a->5	b->2	f->1	g->3	n->1	r->2	s->7	t->3	v->9	
av va	d->12	n->3	p->1	r->5	t->1	
av ve	d->1	r->2	t->5	
av vi	c->4	k->3	l->4	s->8	t->1	
av vo	n->4	
av vä	g->1	l->3	n->1	r->8	x->6	
av vå	r->24	
av yt	t->5	
av Ös	t->2	
av äl	d->1	
av äm	n->1	
av än	d->4	n->1	
av är	 ->1	
av ål	d->1	
av år	 ->5	e->1	h->1	
av ås	i->1	
av åt	e->4	g->10	
av öb	o->1	
av öd	e->1	
av ök	a->4	
av öp	p->4	
av ös	t->2	
av öv	e->3	
av, d	e->1	ä->1	
av, e	f->1	
av, f	r->1	
av, m	e->1	
av, o	c->3	
av, s	o->1	
av, t	r->1	
av, ä	r->1	
av.(S	a->1	
av.. 	(->1	
av.De	 ->1	t->3	
av.Dä	r->1	
av.Ef	f->1	
av.Er	i->1	
av.Ja	g->1	
av.Me	n->1	
av.OL	A->1	
av.Rå	d->1	
av?Vi	l->1	
ava g	a->1	
avale	n->2	s->1	t->1	
avall	p->1	
avanc	e->1	
avand	e->1	
avano	s->2	
avant	 ->1	
avar 	p->1	
avar.	R->1	
avara	n->1	
avare	 ->1	
avarn	a->2	
avars	l->1	
avbro	t->3	
avbru	t->2	
avbry	t->3	
avbrö	t->6	
avdel	n->8	
ave (	C->2	
ave m	å->1	
ave ä	r->1	
ave, 	a->1	
ave- 	p->1	
ave-p	r->2	
aveNä	s->1	
avec 	l->1	
aven 	e->1	f->8	i->1	m->4	o->3	p->7	s->1	
aven,	 ->2	
aven.	D->1	N->1	S->1	V->1	
aven:	 ->1	
avera	n->4	
avere	r->1	t->1	
averi	 ->4	,->1	e->1	
avery	,->1	
avet 	a->3	b->1	f->1	h->2	o->3	p->9	s->1	u->3	
avet,	 ->1	
avet.	E->1	F->1	J->2	N->1	T->1	
avets	 ->2	
avett	e->1	
aveur	o->1	
avfal	l->22	
avfol	k->1	
avför	d->1	s->1	t->1	
avgas	e->1	
avgav	 ->1	
avge 	e->3	
avger	 ->5	
avges	 ->1	
avget	t->1	
avgic	k->4	
avgif	t->4	
avgiv	i->1	
avgjo	r->4	
avgrä	n->4	
avgå.	S->1	
avgåe	n->1	
avgån	g->2	
avgår	 ->1	
avgåt	t->1	
avgör	 ->1	a->57	s->3	
avhjä	l->2	
avhän	d->1	g->1	
avhål	l->1	
avi I	n->1	
avid 	B->2	L->1	
avien	s->1	
avisa	 ->1	n->1	r->2	
avise	r->4	
avisk	 ->1	
avkla	r->1	
avkrä	v->1	
avkun	n->1	
avla 	f->1	s->1	v->1	ä->1	
avla"	 ->2	
avlad	e->1	
avlag	t->1	
avlan	"->1	
avled	d->2	
avlig	e->1	
avliv	a->1	
avlop	p->1	
avläg	g->1	s->9	
avmat	t->1	
avori	t->1	
avpri	c->1	
avrap	p->1	
avreg	l->2	
avrun	d->1	
avrät	t->1	
avs a	v->1	
avs h	a->2	
avs i	 ->2	
avs m	e->1	
avs o	m->1	
avs u	t->1	
avs v	e->1	
avs, 	f->1	m->2	o->1	
avs.A	l->1	
avs.D	e->1	
avs.R	e->1	
avs.V	i->1	
avs?T	i->1	
avsak	n->4	
avsat	t->3	
avse 	f->1	
avsed	d->3	
avsee	n->47	
avser	 ->14	
avses	 ->1	
avset	t->14	
avsev	ä->13	
avsfo	r->1	
avsfö	r->1	
avsid	e->1	
avsik	t->38	
avska	f->19	
avske	d->5	
avski	l->1	
avskr	ä->2	
avsky	 ->1	v->1	
avsla	g->2	
avslo	g->2	
avslu	t->60	
avslä	n->2	
avslå	 ->2	r->1	
avslö	j->6	
avsmi	l->2	
avsni	t->4	
avsom	r->1	
avspe	g->5	
avsta	m->1	
avsto	d->2	
avstä	n->3	
avstå	 ->7	e->1	n->11	r->5	t->2	
avsva	t->1	
avsäg	a->1	
avsät	t->4	
avt s	k->1	
avtal	 ->51	"->1	,->2	.->5	:->1	e->28	s->1	
avtar	.->1	
avtvi	n->1	
avund	s->1	
avvak	t->6	
avvec	k->8	
avver	k->2	
avvik	a->4	e->4	
avvis	a->13	n->2	
avväg	d->2	n->1	
aw, s	o->1	
aw.Me	d->1	
ax av	s->1	
ax ef	t->1	
ax in	n->1	
ax-fr	e->3	
axa e	t->1	
axa u	t->1	
axbel	o->1	
axelr	y->1	
axeri	n->1	
axima	l->6	
axime	r->2	
aximi	å->1	
axis 	a->1	i->1	s->2	ä->1	
axis.	D->1	F->1	
axise	n->1	
axlar	.->1	
ay fö	r->2	
ay ha	r->1	
ay, J	o->1	
ay, a	t->1	
ay, h	a->1	
ay, s	o->1	
ay.Vi	 ->1	
ayDe 	f->1	
ayabe	r->1	
ayabu	k->2	
ayago	l->4	
ayann	a->2	
aybet	ä->1	
ayed 	i->2	
ayern	,->1	
ays b	e->2	
ays d	e->1	
ays-d	e->1	
aza o	c->1	
aza, 	d->1	
aza.D	e->1	
aza.S	i->1	
azaks	t->1	
azare	m->2	
azism	 ->2	.->1	e->5	
azist	 ->1	!->1	e->2	f->1	i->3	
aça M	o->5	
b Söd	e->2	
b eft	e->1	
b had	e->1	
b hjä	l->1	
b kan	 ->1	
b och	 ->3	
b ska	l->1	
b var	n->1	
b) in	f->1	
b) mi	n->1	
b, en	 ->1	
b, so	m->1	
b, sä	r->1	
b, vi	 ->1	
b-omr	å->1	
b.Ans	v->1	
b.Det	 ->1	
ba an	s->1	
ba be	h->1	
ba bi	l->1	
ba fr	a->1	
ba oc	h->1	
ba os	s->1	
ba på	 ->1	
ba re	a->1	
ba ti	l->1	
ba up	p->1	
ba va	r->1	
ba åt	g->1	
ba-, 	S->1	
bacil	l->1	
back-	p->1	
backn	i->1	
bacèt	e->1	
bad F	P->1	
bad e	r->1	
bad k	o->1	
bad o	m->1	
bada 	r->1	
bade 	F->1	T->1	a->1	b->2	d->1	f->1	h->1	i->1	k->1	m->3	o->4	r->3	s->1	
bade.	A->1	T->1	
bades	 ->4	
bads 	b->1	
bagat	e->2	
bain"	,->1	
bak i	 ->1	
bak, 	b->1	
baka 	a->2	b->1	d->5	e->1	f->2	g->2	i->3	j->1	k->1	m->3	o->5	t->9	
baka.	D->1	I->2	M->1	
baka?	I->1	
bakad	r->3	
bakag	å->4	
bakav	i->4	
bakdö	r->1	
bakgr	u->31	
bakom	 ->19	,->1	l->1	
baks 	d->1	
bakso	d->1	
bakte	r->1	
bakåt	 ->2	s->1	
bal n	i->1	
bala 	j->1	k->1	u->1	v->1	ö->1	
balam	,->1	
balan	s->33	
balis	e->5	
ballm	ö->1	
balt 	o->1	
balt,	 ->1	
ban s	o->1	
ban" 	a->1	
bana 	i->1	
banal	i->3	
banan	e->1	
banat	 ->1	
banbr	y->1	
band 	h->1	i->1	m->45	o->1	s->1	
bande	n->1	t->3	
baner	 ->2	,->1	.->1	n->1	
banes	i->1	
banie	n->1	
banis	e->1	
bank 	v->1	
bank"	 ->1	
banke	n->10	r->4	
bankf	ö->1	
banki	r->1	
banks	c->1	e->1	
bannl	y->1	
banon	 ->2	,->1	.->1	?->1	
banor	.->3	
bansk	 ->1	a->3	
banta	s->1	
bantn	i->1	
bar d	e->2	
bar e	n->5	r->1	
bar f	ö->1	
bar g	ä->1	
bar h	e->1	
bar k	o->3	
bar m	e->2	i->1	
bar n	i->1	
bar o	c->1	
bar p	o->2	
bar r	å->1	
bar s	e->1	k->1	t->1	y->2	
bar t	i->1	
bar u	t->12	
bar v	e->2	
bar, 	i->1	
bar.D	e->2	
bar.F	ö->1	
bar.H	e->1	
bara 	"->1	1->2	2->1	5->1	7->1	D->1	I->1	a->16	b->11	d->4	e->53	f->21	g->9	h->8	i->10	j->2	k->9	l->5	m->13	n->14	o->9	p->10	r->2	s->21	t->9	u->10	v->16	y->1	Ö->1	ä->15	å->3	ö->1	
bara,	 ->2	
bara.	A->1	F->1	P->1	
bara:	 ->1	
barba	r->2	
barde	r->1	
bare 	b->1	f->1	o->3	r->1	t->1	ä->1	
bare.	 ->2	E->1	
bargo	 ->1	
barhe	t->9	
barie	t->1	
baris	k->1	
barkb	o->1	
barli	g->12	
barma	n->1	
barn 	i->1	k->1	o->2	s->2	
barn,	 ->3	
barnb	a->1	
barnp	o->2	
barns	 ->1	
barri	ä->2	
bart 	-->1	E->2	a->21	b->2	e->3	f->13	g->3	h->3	i->4	k->2	l->1	m->6	n->1	o->3	p->2	s->11	t->3	u->1	Ö->1	ä->1	
bart!	H->1	
bart,	 ->4	
bart.	A->1	F->2	H->1	I->1	K->2	S->1	V->1	
baréb	e->1	
bas a	v->5	
bas f	ö->1	
bas h	å->1	
bas i	 ->1	
bas o	h->1	
bas p	å->1	
bas, 	h->1	
bas.D	e->1	
basar	!->1	,->1	
baseb	a->1	
basen	 ->5	
baser	a->8	
basis	 ->3	,->1	
baski	s->4	
baskr	a->1	
bassa	d->1	
bast 	t->1	v->1	
baste	 ->1	
basti	a->1	o->1	
bastu	 ->1	
basun	e->1	
bat F	r->1	
bat e	n->1	
bat f	å->1	
bats 	a->5	e->1	h->1	
bats.	J->1	V->1	
batt 	-->1	b->2	d->1	e->1	f->3	g->2	i->7	m->3	o->11	p->2	r->1	s->9	t->1	u->1	v->4	ä->4	
batt,	 ->9	
batt.	D->5	F->2	H->2	J->1	K->1	L->2	M->3	P->1	T->1	U->1	V->2	
batt:	 ->1	
batt?	V->1	
battB	e->1	
batta	n->1	
batte	n->65	r->18	
batti	n->1	
battk	v->1	
baxa 	u->1	
bayer	n->1	
bb ef	t->1	
bb hj	ä->1	
bb oc	h->3	
bb va	r->1	
bb, s	ä->1	
bb, v	i->1	
bba a	n->1	
bba b	e->1	i->1	
bba f	r->1	
bba o	c->1	s->1	
bba p	å->1	
bba r	e->1	
bba t	i->1	
bba u	p->1	
bba v	a->1	
bba å	t->1	
bbade	 ->21	.->2	s->4	
bbar 	d->2	k->1	r->1	
bbare	 ->8	.->3	
bbas 	a->5	h->1	o->1	p->1	
bbast	 ->2	e->1	
bbat 	F->1	e->1	f->1	
bbats	 ->7	.->2	
bbel 	e->1	
bbels	 ->1	k->2	
bbelt	 ->2	
bbelv	ä->1	
bbiga	 ->1	
bbla 	d->1	f->7	k->1	s->1	
bblas	 ->1	
bbpla	t->1	
bbt f	r->4	ö->1	
bbt g	e->2	
bbt h	å->1	
bbt k	a->2	o->1	
bbt l	ä->1	
bbt m	å->2	
bbt o	c->1	
bbt p	å->1	
bbt s	k->2	o->9	v->1	ä->2	
bbt t	a->1	
bbt u	t->1	
bbt v	i->1	ä->1	
bbt, 	a->1	h->1	k->1	
bbt.J	a->1	
bbt.M	e->1	
bbt.O	m->2	
bbt.T	y->1	
bbt.V	i->1	
bbvar	n->1	
bby, 	d->1	
bbyar	b->1	
bbybi	l->1	
bbygr	u->2	
bbyis	t->2	
bbyma	s->1	
bbyn 	h->1	l->1	å->1	
bbyve	r->1	
be Pr	o->1	
be er	 ->5	
be fr	u->1	
be he	r->1	
be ho	n->1	
be ko	m->6	
be om	 ->2	
be pa	r->1	
be st	a->1	
beakt	a->30	
bearb	e->2	
beboe	l->1	
bebyg	g->1	
bebåd	a->1	
bedd 	u->1	
bedre	v->1	
bedri	v->15	
bedrä	g->35	
beds 	a->1	
bedöm	a->15	b->1	d->1	e->4	n->26	s->3	t->1	
befar	a->5	
befat	t->6	
befin	n->31	t->10	
beflä	c->1	
befog	a->5	e->27	
befol	k->43	
befor	d->7	
befra	k->10	
befri	a->3	e->6	
befrä	m->1	
befäl	h->1	
befän	g->1	
befäs	t->10	
begag	n->4	
begra	v->1	
begre	p->13	
begri	p->21	
begru	n->2	
begrä	n->68	
begär	 ->11	.->1	a->34	d->3	s->1	t->10	
begå 	e->1	s->1	
begår	 ->3	
begås	 ->3	
begåt	t->3	
behag	l->2	
behan	d->85	
behov	 ->23	,->2	.->3	e->39	
behäf	t->1	
behål	l->29	
behöl	l->1	
behör	i->18	
behöv	a->16	d->2	e->99	s->27	t->3	
beivr	a->1	
bekan	t->3	
bekis	t->2	
bekla	g->42	
bekom	 ->1	
bekos	t->1	
bekrä	f->30	
bekvä	m->15	
bekym	m->6	r->10	
bekäm	p->41	
bekän	n->1	
bel H	i->1	
bel P	e->1	
bel e	n->1	
bel i	 ->1	
bel l	ö->1	
bel n	i->1	
bel o	c->1	
bel r	e->1	
bel u	t->1	
bel!M	e->1	
bel, 	e->1	o->1	s->2	
bel.D	e->1	
bel.V	i->3	
bel.Ä	r->1	
belag	d->4	
belas	t->10	
belgi	s->8	
bell 	f->3	s->1	
bell.	J->1	M->1	
belop	p->16	
bels 	v->1	
belsk	r->2	
belt 	-->1	E->1	a->3	f->2	m->1	o->3	s->6	t->1	v->1	
belt.	D->1	H->2	I->1	J->1	U->1	V->2	
belt;	 ->1	
belt?	J->1	
belvä	g->1	
belys	a->1	e->1	n->1	t->1	
beläg	g->3	n->4	
belön	a->2	
beman	n->2	
bemyn	d->1	
bemär	k->5	
bemöd	a->3	
bemöt	a->4	e->1	s->2	
ben i	 ->1	
benef	i->5	
benen	 ->1	
benga	 ->1	
benhå	r->1	
beni 	f->1	s->1	
beni.	A->1	
bensi	n->1	
benäg	n->1	
benåd	a->1	
beord	r->1	
ber 1	9->20	
ber V	i->1	
ber a	n->1	t->3	
ber d	e->3	
ber e	n->1	r->6	x->1	
ber f	ö->4	
ber h	a->1	
ber i	 ->2	n->1	
ber j	a->9	
ber k	o->4	
ber l	i->1	o->1	ä->1	
ber m	i->1	å->3	
ber n	ä->1	
ber o	c->4	m->6	s->2	
ber r	i->1	å->1	
ber s	a->1	
ber v	i->1	
ber, 	a->4	d->2	e->1	k->1	l->1	m->1	p->1	r->1	å->1	
ber. 	J->1	
ber.D	e->1	
ber.E	n->1	
ber.J	a->1	
ber.N	u->1	
ber.S	t->1	
berad	 ->1	
beral	 ->2	a->19	d->1	e->3	i->5	t->1	
berba	y->1	
bered	a->10	d->35	e->12	s->2	
beret	t->6	
berg 	f->1	k->1	o->1	
berge	n->1	
berik	a->8	
beris	k->1	
berna	 ->2	
berod	d->5	
beroe	n->68	
berop	a->1	
beror	 ->18	,->1	
berot	t->1	
bert 	C->1	G->1	
berve	c->1	
beryk	t->1	
beräk	n->4	
berät	t->31	
beröm	t->1	v->1	
berör	 ->9	d->21	s->8	t->4	
beröv	a->1	
bes a	t->1	
bes ä	r->1	
beseg	r->2	
besik	t->2	
besit	t->2	
beska	t->4	
beske	d->3	
beskr	e->2	i->21	
besky	d->3	l->2	
beslu	t->220	
beslä	k->1	
beslö	t->1	
bespa	r->5	
besto	d->1	
bestr	a->2	i->2	å->1	
besty	r->1	
bestä	l->4	m->159	n->2	
bestå	 ->4	e->4	n->27	r->18	
bestö	r->1	
besva	r->17	
besvi	k->8	
besvä	r->7	
besyn	n->1	
besät	t->3	
besök	 ->6	a->1	e->1	t->1	
besör	j->2	
bet F	ö->1	
bet d	e->1	
bet h	a->1	
bet m	e->1	
bet o	c->3	
bet s	k->1	o->1	
bet t	i->1	
bet u	t->2	
bet" 	ä->1	
bet",	 ->1	
bet, 	p->1	s->1	u->1	
bet-f	r->1	
bet.E	u->1	
bet.V	i->1	
bet?J	a->1	
beta 	b->1	d->1	e->9	f->13	i->7	k->2	m->16	n->1	o->2	p->6	s->2	t->3	ö->1	
beta,	 ->1	
beta.	 ->1	D->1	T->1	
beta?	V->1	
betad	e->2	
betal	a->73	n->15	t->2	
betan	d->11	e->5	s->5	
betar	 ->21	.->1	e->8	k->1	n->4	
betas	 ->1	.->1	
betat	 ->12	s->2	
bete 	(->2	-->3	a->2	b->3	d->2	f->9	h->6	i->9	k->6	l->3	m->22	o->14	p->6	r->1	s->22	t->1	u->1	v->2	ä->1	å->1	
bete,	 ->11	
bete.	 ->1	.->1	A->1	D->5	F->1	H->1	I->1	J->3	K->1	L->3	M->2	N->1	P->1	R->2	S->1	U->1	V->2	Å->1	
bete?	H->1	I->1	S->1	
betec	k->4	
betee	n->3	
beten	 ->6	a->3	
beter	 ->1	.->1	
betet	 ->39	"->1	,->3	.->7	s->1	
beth 	S->1	
betjä	n->1	
beton	a->45	i->1	
betra	k->23	
betry	g->1	
beträ	f->72	
bets-	 ->2	
betsa	n->4	v->1	
betsb	e->1	ö->5	
betsd	o->4	
betsf	o->1	ö->1	
betsg	i->8	r->5	
betsi	n->2	
betsk	l->1	o->1	r->4	
betsl	i->2	ä->1	ö->43	
betsm	a->13	e->2	ä->2	
betsn	o->3	
betso	r->11	
betsp	e->1	l->9	o->1	r->3	
betsr	a->1	u->2	ä->2	
betst	a->40	i->43	
betsv	i->5	
bett 	o->2	t->1	
betts	 ->2	
betun	g->1	
betvi	v->3	
betyd	a->17	d->1	e->91	l->13	
betän	k->268	
beund	r->3	
bevak	a->3	n->3	
bevar	a->22	
bevek	a->1	
bevil	j->48	
bevis	 ->22	,->1	.->2	a->6	b->7	e->4	n->1	
bevit	t->1	
bexpl	o->1	
bi de	n->1	
bi nä	r->1	
bibeh	å->11	
bibli	o->2	
bidra	 ->35	,->1	g->52	r->20	
bidro	g->3	
bieff	e->2	
bifal	l->3	
bifar	t->2	
biga 	o->1	
bigot	t->1	
bigå 	d->1	
bigåe	n->4	
bigås	 ->1	
bihan	;->1	
bikme	t->2	
bil e	l->1	
bil f	ö->1	
bil g	r->2	
bil i	 ->1	
bil k	o->1	
bil o	c->1	
bil s	o->4	
bil v	e->1	
bil, 	s->1	t->1	
bil- 	o->1	
bil. 	E->1	
bil.D	e->1	
bil.T	r->1	
bila 	b->1	
bilag	a->4	o->2	
bilar	 ->42	,->14	.->13	?->1	b->1	e->1	n->10	
bilat	e->6	
bilbe	s->1	
bilbr	a->1	
bild 	a->2	b->1	m->1	
bild,	 ->1	
bild.	D->1	N->1	
bilda	 ->6	d->3	n->5	r->6	s->5	t->3	
bilde	l->3	n->2	r->2	
bildn	i->66	
bilen	 ->3	,->2	.->2	
bilin	d->29	
bilis	e->10	t->1	
bilit	e->27	
biljo	n->1	
bilko	n->1	
bilky	r->1	
bilkö	p->2	
billi	g->6	
bilmä	r->1	
bilpa	r->6	
bilpr	o->1	
bils 	l->2	
bilse	k->1	
bilsk	r->2	ö->1	
bilsp	r->1	
bilt 	g->1	j->1	
bilti	l->15	
bilvr	a->6	
biläg	a->1	
bilåt	e->1	
bin, 	r->1	
binat	i->1	
binda	 ->2	n->12	
binde	l->15	r->8	
binet	t->3	
bio s	a->1	
biogr	a->1	
biolo	g->4	
biopl	a->1	
biosf	ä->1	
biosä	k->2	
bisee	n->1	
bisen	.->1	
bisk 	b->1	m->1	
bisk-	i->1	
biska	 ->9	
bistå	 ->1	n->21	t->1	
bit p	å->1	
biter	 ->1	
bitio	n->14	
bitiö	s->12	
bitte	r->2	
bittr	a->1	
bjekt	"->1	i->1	
bjuda	 ->15	n->5	s->2	
bjude	n->1	r->11	t->4	
bjudi	t->1	
bjudn	a->2	i->1	
bjöd 	f->1	
bjöds	 ->1	
bl.a.	 ->27	
bla a	t->1	
bla d	e->1	i->1	
bla e	f->1	
bla f	a->7	i->1	ö->1	
bla i	 ->1	n->1	
bla k	ö->1	
bla o	c->1	
bla s	a->1	i->1	k->1	n->1	
bla t	r->1	
bla".	H->1	
bla, 	v->1	
bla.D	e->1	
bla.M	e->1	
bla.N	ä->1	
bla.Ö	v->1	
blad 	s->1	
blame	r->1	
blanc	a->1	
bland	 ->69	a->18	e->1	n->10	s->1	
blank	o->1	t->1	
blare	 ->1	.->1	
blas 	t->1	
bleka	s->1	
blem 	-->1	a->1	d->2	e->3	f->3	h->2	i->11	k->2	m->12	n->4	o->5	p->1	s->17	v->3	ä->4	ö->1	
blem,	 ->13	
blem.	 ->1	.->1	A->1	D->6	F->1	H->2	I->1	J->3	P->1	S->2	V->3	
blem:	 ->1	
blem;	 ->2	
blem?	M->1	
blema	t->5	
bleme	n->17	t->48	
blemo	m->3	
bler 	o->1	
blera	 ->5	d->4	t->2	
bleri	n->3	
bles 	G->1	
blev 	a->3	d->2	f->2	i->2	k->1	o->3	t->1	u->1	
bli -	 ->1	
bli 2	0->1	
bli a	k->1	l->2	n->2	t->4	v->2	
bli b	e->3	r->1	ä->1	
bli d	e->3	o->2	
bli e	f->2	n->18	t->11	
bli f	l->2	r->1	ä->1	ö->8	
bli g	a->1	
bli h	e->1	
bli j	u->1	
bli k	l->3	o->1	
bli l	e->1	i->2	ä->1	
bli m	e->11	i->2	y->5	ö->3	
bli n	ä->1	å->2	ö->2	
bli o	b->1	m->1	t->1	
bli p	l->1	r->2	
bli r	i->1	
bli s	l->1	t->3	u->1	v->1	y->1	ä->1	å->1	
bli t	v->3	
bli v	a->1	e->2	å->1	
bli ä	m->1	
bli ö	v->2	
bli, 	e->1	
bli.U	t->1	
blic 	-->1	
blice	r->4	
blici	t->1	
blick	 ->4	,->1	.->2	a->2	b->5	e->10	
bliga	t->14	
blik 	h->1	p->1	
blika	n->6	
blike	n->10	r->2	
blin 	b->1	o->2	s->1	
blin.	L->1	
blind	a->1	
blink	o->2	
blint	 ->1	
bliot	e->2	
blir 	E->2	a->10	b->3	d->14	e->10	f->6	g->1	h->3	i->5	j->2	k->1	l->5	m->11	n->5	o->4	r->3	s->13	t->5	u->2	v->4	ä->1	å->1	ö->1	
blir,	 ->2	
blir:	 ->1	
bliva	n->1	
blivi	t->26	
blixt	r->1	
block	a->2	b->1	e->3	
blomm	a->1	o->2	
bloms	t->3	
blonm	ä->1	
blott	 ->1	a->2	
blund	a->4	
bly å	t->1	
bly, 	k->2	
bly.V	i->1	
blygs	a->4	
blå b	a->1	
blåse	r->2	
bning	a->1	
bo i 	l->1	
bo kv	a->1	
bo vi	l->1	
board	,->1	
bock"	 ->1	
bocka	r->1	
boda 	h->1	o->1	
bodas	 ->1	
boeli	g->1	
boend	e->3	
bogse	r->1	
bojko	t->1	
bok a	v->1	
bok h	e->1	
bok m	e->1	
bok o	m->7	
bok s	k->1	o->2	
bok t	i->1	
bok ä	r->2	
bok, 	d->1	
bok.D	e->1	
bok.H	u->1	
bok.J	a->1	
bok.T	a->1	
bok.V	i->1	
boken	 ->29	,->1	.->4	:->1	s->1	
boksl	u->1	
bokst	a->1	
bol f	ö->2	
bolag	 ->3	,->1	e->8	
bolis	k->6	m->1	
bolls	b->1	
bomb 	h->1	
bomb.	A->1	
bomba	r->1	t->1	
bombe	n->1	r->2	x->1	
bombn	i->1	
bomul	l->1	
bon f	ö->1	
bon g	ö->1	
bon k	o->1	
bon m	.->1	
bon, 	D->1	
bon.V	a->1	
bondg	å->2	
bonmö	t->2	
bor d	ä->1	
bor i	 ->4	
bor p	å->1	
borat	o->3	
bord 	i->1	o->2	
bord.	B->1	
borda	d->1	n->1	r->1	
borde	 ->65	.->1	t->4	
bordl	a->1	
bords	u->1	
borg 	t->1	
borga	r->168	
borge	r->3	
borgm	ä->2	
borre	n->1	
bort 	-->1	a->4	f->5	i->2	k->2	n->2	o->1	p->1	s->2	
bort,	 ->5	
bort.	D->4	V->2	
borta	 ->1	
bortf	a->6	
borto	m->2	
bortp	r->1	
borts	e->6	
bosat	t->3	
bosni	e->2	
bosta	d->1	
bostä	d->4	
bosät	t->4	
bot p	å->2	
botar	 ->2	
botte	n->5	
bottn	a->3	e->1	
bourg	 ->2	.->3	
bovar	 ->1	
boven	 ->1	
boxni	n->1	
bplat	s->1	
bra a	r->2	t->8	v->1	
bra b	a->1	e->3	i->1	
bra d	a->1	e->1	i->2	ä->1	
bra e	l->1	x->1	
bra f	ö->3	
bra i	 ->2	d->1	
bra j	o->1	
bra m	e->1	i->4	
bra n	y->2	
bra o	c->6	m->3	
bra s	y->1	ä->8	
bra t	i->1	
bra u	r->1	t->3	
bra v	i->1	
bra ä	n->2	
bra å	t->1	
bra!M	ä->1	
bra, 	d->2	e->1	g->1	i->1	m->2	o->1	
bra.D	e->1	
bra.E	n->1	
bra.J	a->1	
bra.P	a->1	
bra.S	o->1	
bra.V	i->1	
brand	 ->1	e->1	m->1	
brans	c->7	
bred 	b->1	d->1	e->1	l->1	
breda	 ->1	,->1	r->3	s->1	
bredd	e->2	
brede	r->1	
bredn	i->4	
breis	k->1	
brepu	b->1	
breta	g->1	
brett	 ->6	
brev 	d->1	f->1	s->1	t->1	
brev.	F->1	
brevl	å->1	
brief	i->1	
brien	 ->2	.->1	
brigh	t->1	
brike	r->3	
bring	a->13	
brist	 ->19	a->12	e->23	f->8	
brita	n->14	
britt	e->2	i->15	
bro m	e->1	
bro o	c->1	
broar	 ->1	
brode	r->2	
broki	g->2	
brome	r->4	
broms	 ->1	a->4	v->1	
bron-	 ->1	
bror,	 ->1	
broth	e->1	
brott	 ->10	,->6	.->4	a->2	e->4	m->1	s->26	
brotu	l->1	
bruar	i->16	
bruk 	a->1	m->1	o->5	p->1	s->1	
bruk!	A->1	
bruk,	 ->9	
bruka	d->2	r->14	s->1	
bruke	n->1	t->19	
brukn	i->1	
bruks	e->1	f->2	l->1	o->2	p->9	r->2	s->6	
bruna	 ->1	
bruta	l->1	
brute	n->1	t->1	
bruti	t->2	
brutt	o->1	
brygg	a->3	
bryos	t->1	
bryr 	e->1	j->1	
bryta	 ->6	n->1	s->1	
bryte	l->2	r->6	
brytn	i->2	
bränd	a->2	e->1	
bränn	a->3	i->2	
bräns	l->7	
bräsc	h->2	
bråds	k->20	
bråke	t->1	
brås 	f->2	
bröd.	-->1	D->2	
bröst	t->1	
bröt 	h->1	t->4	
bröts	 ->2	
bserv	a->1	e->1	
bsida	r->1	
bsidi	a->21	ä->1	
bsolu	t->40	
bsorb	e->1	
bstan	s->2	t->2	
bstat	 ->1	e->1	
bstra	k->1	
bsurd	 ->1	
bsurt	 ->2	
bt fr	a->3	i->1	
bt fö	r->1	
bt ge	n->1	t->1	
bt hå	l->1	
bt ka	n->2	
bt ko	m->1	
bt lä	m->1	
bt må	s->2	
bt oc	h->1	
bt på	 ->1	
bt sk	a->1	u->1	
bt so	m->9	
bt sv	a->1	
bt sä	g->1	t->1	
bt ta	 ->1	
bt ut	t->1	
bt vi	l->1	
bt vä	x->1	
bt, a	t->1	
bt, h	o->1	
bt, k	r->1	
bt.Ja	g->1	
bt.Me	l->1	
bt.Om	 ->2	
bt.Ty	 ->1	
bt.Vi	 ->1	
bu in	l->1	
bud e	l->1	
bud f	a->1	ö->4	
bud m	e->2	o->7	
bud o	c->4	
bud r	e->1	
bud v	i->1	
bud ä	r->1	
bud, 	a->1	e->1	h->1	s->1	
bud.D	e->2	
bud.V	a->1	
buddh	i->1	
budet	 ->7	,->1	?->1	
budge	t->106	
budor	d->1	
budsf	ö->3	
budsi	n->3	
budsk	a->10	
budsm	a->10	
budsp	r->1	
bugge	n->1	
bukte	n->2	
bul f	ö->1	
bulan	s->1	
bular	y->1	
bulte	n->1	
bunde	n->4	t->9	
bundi	t->3	
bundn	a->4	
bunds	k->1	l->2	r->5	
buret	 ->1	
burg 	f->1	i->1	m->1	u->1	
burg,	 ->4	
burg.	D->1	
burga	r->1	
burgh	.->1	
burit	 ->1	
burna	.->1	
bus ä	r->1	
bussa	r->2	
butik	 ->1	
butio	n->1	
bvarn	i->1	
bvent	i->12	
bvärl	d->1	
by, d	e->1	
byarb	e->1	
bybil	a->1	
byens	 ->1	
bygd 	i->1	o->1	
bygd.	D->2	
bygde	n->31	
bygds	b->1	k->1	o->4	r->2	t->1	u->1	
bygga	 ->32	n->22	s->3	
byggd	 ->2	e->2	
bygge	 ->1	l->1	r->7	t->3	
byggn	a->19	
byggs	 ->2	t->1	
byggt	 ->4	s->1	
bygru	p->2	
byist	e->2	
bymas	k->1	
byn h	a->1	
byn l	y->1	
byn å	l->1	
byrå 	s->1	ä->1	
byråe	r->1	
byråk	r->30	
byrån	 ->2	
byta 	e->1	h->1	
byte 	a->3	f->2	k->1	m->3	s->1	
byte,	 ->1	
bytet	 ->6	
bytts	 ->1	
byver	k->1	
byxfi	c->1	
bälte	 ->2	,->2	n->2	t->4	
bänke	n->1	
bär a	l->1	n->5	t->45	
bär b	a->1	ö->1	
bär d	e->3	i->2	
bär e	n->11	t->4	
bär f	r->1	ö->4	
bär i	 ->4	n->5	
bär l	ä->1	
bär m	e->1	i->1	
bär n	å->1	
bär o	c->3	l->1	
bär p	å->4	
bär s	k->1	t->1	å->1	
bär u	p->1	
bär v	i->1	
bär ä	r->1	
bär ö	v->1	
bär, 	i->1	
bär.D	ä->1	
bär.F	ö->1	
bära 	a->10	e->3	f->1	h->3	i->1	k->2	m->1	p->1	s->3	
bäran	d->2	
bäras	 ->3	
bärli	g->4	
bärs 	f->1	s->1	
bäst 	a->1	g->1	k->1	r->1	t->1	
bästa	 ->34	.->3	
bättr	a->60	e->75	i->18	
bävni	n->10	
båda 	a->1	b->1	d->4	e->1	f->5	i->1	l->2	m->1	o->3	p->1	s->3	
båda,	 ->1	
bådad	e->1	
bådan	d->1	
både 	D->1	S->2	a->1	b->2	d->6	e->2	f->2	g->1	h->2	i->6	k->1	m->5	n->1	p->4	r->2	s->4	t->1	v->2	ö->1	
båtar	 ->5	,->2	n->1	
båten	s->1	
bé av	e->1	
bébé 	a->1	
böcke	r->3	
bödel	s->1	
böjel	s->1	
böjt 	s->1	
böld 	m->1	
bör "	i->1	
bör -	 ->1	
bör E	u->3	
bör a	b->2	l->3	n->1	r->2	v->2	
bör b	e->4	i->2	l->2	
bör d	e->12	i->1	o->2	ä->1	
bör e	m->1	r->4	
bör f	a->1	i->2	o->2	r->1	u->2	å->3	ö->7	
bör g	e->3	r->1	ö->8	
bör h	a->4	å->1	ö->1	
bör i	 ->2	n->12	
bör k	o->5	r->1	u->1	
bör l	i->2	ä->4	
bör m	a->23	i->1	
bör n	i->1	o->3	
bör o	c->5	m->1	
bör s	a->2	e->3	j->1	l->1	n->1	p->1	t->1	
bör t	.->1	a->3	v->1	y->1	
bör u	n->4	p->3	t->5	
bör v	a->14	e->3	i->10	ä->1	å->1	
bör ä	g->1	v->3	
bör å	t->4	
bör ö	v->2	
bör, 	o->1	
bör.F	ö->1	
böran	d->1	
börd.	D->1	
börda	 ->5	,->1	.->2	?->1	n->8	
börde	n->6	
bördo	r->2	
börja	 ->59	d->8	n->19	r->17	t->12	
börli	g->10	
börse	n->1	r->1	
böter	 ->1	
c - o	c->1	
c Bra	v->1	
c bli	r->1	
c bör	 ->1	
c då 	d->1	
c i E	K->1	
c i d	e->1	
c l'e	a->1	
c osv	.->1	
c ser	 ->1	
c", f	ö->1	
c) li	k->1	
c, dv	s->1	
c-dir	e->1	
c-sys	t->1	
c-tra	n->1	
c. oc	h->1	
c. Äm	n->1	
c. Äv	e->1	
c.Det	 ->1	
c.En 	v->1	
c?Att	 ->1	
cCart	h->1	
cNall	y->5	
ca 30	 ->1	
ca Co	l->1	
ca Mo	u->3	
ca sa	d->1	
ca, o	c->1	
ca. 1	2->1	
cal c	o->1	
calvi	n->1	
cance	r->2	
canna	b->1	
cante	 ->1	
cao t	i->1	
cap ä	r->1	
capit	a->10	
cas s	k->1	
case.	O->1	
cayab	u->2	
cayag	o->4	
ccept	a->44	e->45	
ccess	i->5	
ce bö	r->1	
ce de	l->2	n->2	
ce fö	r->1	
ce na	t->1	
ce oc	h->1	
ce or	d->11	
ce ta	l->2	
ce, D	a->1	
ce...	)->1	
ce.Al	l->1	
ce.De	n->1	
ce.Ja	g->2	
ce.Of	f->1	
ce.St	ä->1	
cedo 	a->1	
cedur	r->1	
cekor	t->1	
cekva	l->1	
celon	a->2	
cembe	r->19	
cemen	t->2	
cemis	-->1	
cen m	e->1	
cen, 	o->1	
cenar	i->5	
cenen	.->1	
cenni	e->6	u->1	
censa	t->1	
censi	n->1	
cent 	(->1	-->1	1->1	a->44	b->1	e->4	f->1	g->1	h->1	i->4	k->4	m->3	o->3	p->2	s->1	t->3	u->1	v->1	
cent,	 ->2	
cent.	D->4	F->1	H->1	M->2	S->1	V->1	
centa	n->8	
cente	n->6	r->8	
centi	m->1	
centr	a->84	e->16	u->9	
cents	 ->3	a->1	i->1	
cept 	i->1	k->1	
cept.	D->1	H->1	
cepta	b->37	n->7	
cepte	r->45	t->3	
cepti	o->6	
cer!D	e->1	
cer, 	h->1	
cera 	a->1	d->1	e->1	f->1	l->1	m->3	o->1	t->1	u->2	
cerad	 ->14	.->3	e->14	
ceran	d->3	
cerar	 ->5	.->2	
ceras	 ->5	
cerat	 ->11	,->2	.->2	s->2	
cerbö	l->1	
cerin	g->13	
cerne	r->2	
certi	f->6	
cess 	a->4	f->1	i->2	k->2	m->4	o->1	s->8	
cess"	.->1	
cess,	 ->2	
cess.	A->1	D->4	H->1	M->2	N->1	V->4	
cess?	J->1	
cesse	n->54	r->12	
cessi	v->5	
cessr	e->1	ä->2	
cessu	e->1	
ceuti	q->1	
ch "U	r->1	
ch "s	k->1	
ch "t	i->1	
ch (A	5->1	
ch - 	e->1	s->2	
ch -o	r->3	
ch 0 	p->1	
ch 1-	2->1	
ch 10	 ->1	0->1	
ch 13	8->1	
ch 14	 ->1	
ch 16	 ->1	
ch 17	 ->1	.->1	
ch 19	 ->1	4->1	9->11	
ch 2 	i->1	
ch 2,	 ->1	
ch 2.	D->1	
ch 20	 ->2	0->1	
ch 21	 ->3	
ch 22	.->1	
ch 25	.->1	
ch 27	 ->1	
ch 29	 ->1	
ch 3.	I->1	
ch 30	 ->1	0->1	
ch 33	 ->1	
ch 34	 ->1	
ch 35	.->1	
ch 3:	 ->1	
ch 4.	J->1	
ch 41	 ->2	
ch 45	 ->2	,->1	.->1	
ch 47	 ->1	
ch 48	 ->2	
ch 5 	v->1	
ch 5.	E->1	
ch 53	 ->1	
ch 60	-->1	
ch 68	 ->1	
ch 7 	-->1	f->1	i->1	o->1	
ch 7,	 ->2	
ch 8 	ä->1	
ch 8,	 ->1	
ch 82	 ->2	)->1	,->3	
ch 86	 ->2	
ch 89	 ->1	
ch 9 	i->1	m->1	
ch 92	/->1	
ch 94	 ->1	
ch Al	b->1	t->1	
ch Am	s->1	
ch An	k->1	
ch BP	,->1	
ch Ba	s->1	
ch Be	l->1	
ch Br	a->1	o->1	
ch Bu	l->1	
ch C.	 ->1	
ch CE	C->1	
ch Ca	u->1	
ch Cy	p->1	
ch Da	n->2	
ch De	 ->1	m->1	
ch EL	D->2	
ch EU	 ->2	-->1	G->1	
ch Ed	i->1	
ch El	m->2	
ch Em	i->1	
ch Er	k->1	
ch Et	i->1	
ch Eu	r->24	
ch FN	:->1	
ch FP	Ö->1	
ch Fi	n->2	
ch Fr	a->10	u->1	
ch Ga	l->1	z->1	
ch Ge	m->1	
ch Go	l->1	
ch Gr	a->1	e->1	u->1	
ch He	l->1	
ch Hi	t->1	
ch Hu	h->1	
ch II	 ->1	,->1	
ch In	d->2	t->2	
ch Ir	l->2	
ch Is	r->5	
ch It	a->1	
ch Ja	c->1	
ch Jö	r->1	
ch Ka	s->1	
ch Ki	n->5	r->1	
ch Ko	u->1	
ch Ku	l->1	
ch La	n->3	
ch Le	i->5	
ch MA	R->1	
ch Ma	d->3	
ch Me	d->1	
ch No	r->1	
ch Ny	a->1	
ch OL	A->1	
ch On	e->1	
ch PP	E->1	
ch PS	E->2	
ch Pa	c->1	k->3	l->4	r->1	
ch Po	r->2	
ch Pr	í->1	
ch Ra	f->2	p->1	
ch Sa	m->10	
ch Sc	h->1	
ch Si	m->1	
ch Sj	ö->1	
ch So	c->1	
ch Sp	a->1	
ch St	o->2	
ch Sw	o->1	
ch Sy	d->1	r->7	
ch Ta	d->1	i->1	m->2	
ch Ts	a->1	
ch Tu	r->1	
ch Ty	s->2	
ch Uz	b->1	
ch Vi	t->1	
ch Vä	s->1	
ch Wy	e->1	
ch X 	o->1	
ch ab	s->1	
ch ac	c->1	
ch ad	m->1	v->1	
ch ag	e->2	
ch ak	t->4	
ch al	d->2	l->16	
ch am	b->4	
ch an	a->3	d->27	g->3	n->3	p->2	s->12	t->5	v->3	
ch ap	r->1	
ch ar	b->14	t->1	
ch as	s->1	y->3	
ch at	t->150	
ch av	 ->14	d->1	g->3	l->1	r->2	s->6	t->3	v->2	
ch ba	d->1	g->1	l->3	n->1	r->7	
ch be	a->1	d->8	f->7	g->2	h->7	k->4	l->4	m->1	r->3	s->5	t->6	v->4	
ch bi	d->6	l->4	
ch bl	.->2	a->2	i->3	u->1	
ch bo	r->2	s->2	t->1	
ch br	a->1	i->2	o->2	u->2	ä->3	å->5	
ch bu	d->3	
ch by	r->2	
ch bä	s->2	t->2	
ch bå	t->1	
ch bö	r->6	
ch ca	l->1	n->1	
ch ce	n->6	
ch ch	e->1	o->1	
ch da	g->2	m->1	t->1	
ch de	 ->83	b->2	c->1	l->8	m->10	n->108	r->12	s->35	t->208	
ch di	a->1	o->1	r->3	s->4	t->2	
ch dj	u->3	ä->1	
ch do	m->9	
ch dr	a->2	i->2	
ch du	k->1	
ch dy	r->1	
ch dä	r->83	
ch då	 ->22	,->1	l->1	
ch dö	t->1	
ch ef	f->16	t->18	
ch eg	e->1	
ch ej	 ->1	
ch ek	o->22	
ch el	e->1	
ch en	 ->70	,->1	a->1	d->2	e->2	g->2	h->5	k->1	l->2	s->1	t->2	v->1	
ch er	 ->2	.->1	a->2	b->2	f->3	h->1	k->2	s->3	t->1	
ch et	i->1	t->32	
ch eu	r->9	
ch ex	a->2	p->1	t->1	
ch fa	k->2	l->2	r->3	s->1	t->5	u->1	
ch fe	d->1	l->1	m->1	
ch fi	e->1	n->8	r->1	s->2	
ch fl	e->8	o->1	y->1	
ch fo	d->1	l->2	r->4	
ch fr	a->25	e->2	i->6	o->2	u->4	ä->34	å->10	
ch fu	l->5	n->2	s->2	
ch fy	r->1	s->1	
ch fä	l->1	
ch få	 ->4	g->1	r->5	t->2	
ch fö	l->5	r->163	
ch ga	g->1	r->6	
ch ge	 ->10	m->6	n->20	o->1	r->3	s->3	
ch gi	v->4	
ch gj	o->1	
ch gl	a->1	o->1	ä->1	
ch go	d->1	t->1	
ch gr	a->2	u->5	ä->2	ö->1	
ch gä	l->1	
ch gå	 ->2	r->2	
ch gö	r->17	
ch ha	 ->2	m->1	n->27	r->14	
ch he	l->7	n->4	r->43	
ch hi	t->1	
ch hj	ä->4	
ch ho	b->1	n->1	p->5	t->4	
ch hu	m->1	n->1	r->11	s->1	v->1	
ch hy	g->1	l->1	
ch hä	l->1	r->8	
ch hå	l->16	
ch hö	g->4	j->2	
ch i 	G->1	M->1	N->1	S->1	T->2	a->1	b->1	d->13	e->3	f->5	g->4	h->1	i->1	j->1	k->1	l->1	m->1	n->1	o->1	p->2	r->1	s->16	u->2	v->8	ö->4	
ch ib	l->3	
ch ic	k->2	
ch id	e->2	r->3	
ch if	r->1	
ch ik	r->1	
ch il	l->1	
ch im	a->1	m->1	
ch in	d->6	f->11	g->7	h->1	i->2	k->1	l->1	n->3	o->7	p->1	r->12	s->12	t->72	v->6	
ch ir	l->1	
ch is	r->2	
ch ja	g->149	
ch jo	r->5	
ch ju	r->3	s->4	
ch jä	m->1	
ch ka	b->1	m->1	n->14	p->1	r->2	t->2	
ch ki	n->1	
ch kl	a->3	o->1	
ch kn	u->1	
ch ko	h->1	l->2	m->61	n->57	r->5	s->3	
ch kr	a->5	e->1	i->6	y->1	ä->4	å->1	
ch ku	l->3	n->4	
ch kv	a->2	i->8	
ch kä	l->1	m->1	r->4	
ch kö	r->1	
ch la	g->6	n->10	r->1	
ch le	d->13	g->1	m->1	v->1	
ch li	k->7	t->1	v->3	
ch lj	u->1	
ch lo	c->1	k->4	s->1	v->3	
ch lu	k->1	
ch ly	c->3	
ch lä	c->1	g->6	m->2	n->1	r->1	t->3	
ch lå	n->11	s->1	t->7	
ch lö	s->2	
ch ma	k->1	n->18	r->1	t->1	
ch me	d->121	k->1	l->3	n->2	r->15	t->1	
ch mi	g->1	l->18	n->17	s->3	
ch mo	d->4	n->6	r->3	t->11	
ch mu	s->1	
ch my	c->7	n->1	
ch mä	n->11	r->1	
ch må	h->1	l->6	n->10	s->5	
ch mö	j->8	r->1	
ch na	t->11	
ch ne	d->1	g->1	o->1	p->4	u->1	
ch ni	 ->8	v->1	
ch no	g->3	r->1	t->1	
ch nu	 ->11	
ch ny	a->5	e->1	l->3	n->2	t->2	
ch nä	r->14	t->2	
ch nå	g->5	
ch nö	d->6	
ch oa	c->4	
ch ob	e->2	
ch oc	h->1	k->8	
ch od	e->1	
ch oe	g->1	k->1	
ch of	f->3	t->2	ö->1	
ch oj	ä->1	
ch ok	l->3	r->1	
ch ol	i->5	j->1	y->2	
ch om	 ->22	b->2	e->3	f->5	g->3	r->2	s->4	
ch on	t->1	
ch op	e->1	p->1	
ch or	d->3	g->2	i->1	s->1	ä->1	
ch os	s->2	t->1	ä->2	
ch ot	v->1	
ch ou	m->1	n->1	t->1	
ch pa	p->1	r->23	s->1	
ch pe	k->2	r->7	
ch pl	a->1	i->2	
ch po	l->15	s->2	
ch pr	a->1	e->3	i->8	o->19	ä->1	
ch på	 ->22	m->1	p->1	s->2	t->1	v->2	
ch ra	p->1	s->4	t->2	
ch re	c->1	d->2	f->4	g->34	j->1	k->2	l->3	n->5	p->1	s->11	v->2	
ch ri	g->1	k->6	n->1	s->1	
ch ro	l->1	m->3	
ch ru	t->1	
ch rä	d->1	k->1	t->59	
ch rå	d->39	
ch rö	s->1	
ch sa	m->40	n->3	
ch se	 ->6	d->9	k->3	l->1	n->1	r->5	t->1	x->3	
ch si	f->1	n->3	s->3	t->3	
ch sj	u->1	ä->3	ö->2	
ch sk	a->14	i->1	o->1	r->1	u->3	y->4	ä->2	ö->4	
ch sl	a->1	u->20	ä->3	
ch sm	u->1	å->1	
ch sn	a->3	å->1	
ch so	c->40	l->2	m->92	
ch sp	a->1	e->4	r->4	
ch st	a->12	i->1	o->3	r->19	ä->7	å->5	ö->14	
ch su	c->1	v->4	
ch sv	a->4	å->8	
ch sy	f->2	n->1	r->1	s->12	
ch sä	g->7	k->12	n->1	r->11	t->2	
ch så	 ->21	d->4	l->2	s->1	
ch sö	d->1	r->1	
ch t.	o->1	
ch ta	 ->5	c->6	k->1	l->4	n->1	r->1	s->2	
ch te	k->2	l->4	
ch th	e->1	
ch ti	d->3	g->1	l->52	n->2	s->1	t->1	
ch tj	o->1	ä->3	
ch to	g->1	l->3	p->1	t->1	
ch tr	a->9	e->2	o->5	å->2	
ch tu	n->1	r->14	s->2	
ch tv	å->3	
ch ty	d->13	v->1	
ch tä	m->1	n->1	p->1	
ch un	d->17	g->6	i->2	
ch up	p->24	
ch ut	a->5	b->4	e->1	f->2	g->4	i->1	l->1	n->2	o->1	r->2	s->4	t->3	v->26	ö->1	
ch va	d->10	l->13	n->4	p->3	r->22	
ch ve	k->1	m->2	r->9	t->11	
ch vi	 ->86	a->1	d->6	k->3	l->13	n->1	s->13	
ch vä	d->1	g->2	l->12	n->2	p->1	r->4	x->4	
ch vå	l->1	r->11	
ch vö	r->1	
ch yn	g->1	
ch yr	k->1	
ch yt	l->1	t->4	
ch ÖV	P->1	
ch Ös	t->6	
ch äg	a->1	n->1	
ch än	 ->4	d->5	n->3	
ch är	 ->9	e->1	
ch äv	e->31	
ch å 	a->4	
ch åk	l->1	
ch ås	a->1	i->1	t->1	
ch åt	e->26	g->3	
ch ök	a->3	
ch öm	s->1	
ch ön	s->1	
ch öp	p->13	
ch ör	e->1	
ch ös	t->4	
ch öv	e->16	r->4	
ch! U	r->1	
ch)De	t->1	
ch, d	e->1	
ch, f	r->1	ö->2	
ch, h	e->1	
ch, i	 ->1	
ch, n	å->1	
ch, r	e->1	
ch, s	l->1	o->3	
ch, t	r->1	
ch, u	t->1	
ch.Ef	t->1	
ch.Ja	g->1	
ch/el	l->1	
ch: V	e->1	
ch?Fr	u->1	
chI o	k->1	
chII.	 ->1	
chabl	o->1	
chand	e->1	
chans	 ->6	e->6	
chape	a->1	
chara	d->1	
chard	 ->1	-->1	
chart	r->1	
che B	a->1	
check	 ->1	
chef 	h->1	
chefe	n->1	r->15	
chema	 ->1	
chen 	f->1	i->1	s->1	v->1	
chen.	F->1	
chen;	 ->1	
cheng	e->10	
cher 	i->1	o->1	v->1	
chera	r->1	
chern	a->2	
chez 	t->1	
chhof	e->1	
chiel	 ->1	
chist	i->1	
chler	 ->1	,->1	.->1	s->1	
chner	 ->3	,->3	s->6	
chock	 ->1	a->1	e->2	
chokl	a->1	
chrey	e->3	
chroe	d->14	
chröd	e->1	
chs i	 ->1	
cht m	e->1	
cht o	c->1	
cht.D	e->1	
chter	s->2	
chtfö	r->3	
chtid	 ->1	
chulz	 ->3	
chwar	z->1	
chwei	z->1	
chwit	z->1	
chyre	g->1	
chörl	i->1	
chüss	e->4	
cial 	d->2	o->4	r->2	s->11	t->3	u->8	
cial-	 ->1	
ciala	 ->78	
cialb	e->2	
ciald	e->15	o->1	
cialf	o->17	r->5	ö->6	
ciali	n->1	s->40	
cialp	o->4	r->1	
cialt	 ->16	,->1	.->1	
cialu	t->1	
ciden	t->1	
ciell	 ->4	a->21	t->24	
cien,	 ->2	
cient	e->1	i->1	
cieri	n->1	
ciety	 ->1	
cific	e->2	
cifik	 ->3	a->17	t->7	
cil -	,->1	
cill 	a->1	
cilov	o->1	
ciner	 ->1	
cio S	á->1	
cio V	a->3	
cio f	ö->1	
cio h	a->1	
cio s	k->1	å->1	
cio, 	a->1	s->1	t->1	
cio.J	a->1	
cio.N	ä->1	
cio: 	v->1	
cioek	o->3	
cios 	i->1	å->1	
cip a	l->1	t->2	
cip e	l->1	n->2	
cip f	ö->1	
cip i	 ->2	n->5	
cip o	c->2	m->2	
cip r	å->1	
cip s	o->4	å->1	
cip ä	r->3	v->1	
cip, 	g->1	m->1	o->1	
cip.J	a->1	
cip.S	j->1	
cip.V	i->2	
cipen	 ->72	,->11	.->16	:->2	N->1	
ciper	 ->28	,->4	.->5	:->1	n->10	
cipes	 ->1	
cipie	l->8	
cipli	n->14	
cipsk	ä->1	
cirka	 ->4	
cirke	l->1	
cirkl	a->2	
cirku	l->3	
cis W	u->1	
cis a	n->1	
cis d	e->4	
cis e	t->1	
cis f	u->1	ö->1	
cis h	a->1	
cis i	n->1	
cis l	i->5	
cis p	å->1	
cis s	a->1	k->1	o->19	
cis v	a->1	
cis-p	r->1	
cisa 	i->1	
ciser	a->7	i->4	
cism,	 ->1	
cisme	n->2	
cist 	b->1	n->1	s->1	
ciste	r->3	
cisti	s->5	
cit.F	ö->1	
citam	e->8	
citat	.->1	
citer	a->7	
citet	 ->4	,->1	.->1	e->1	
civil	 ->5	-->1	a->3	b->2	f->2	i->2	r->1	s->2	t->1	
ck - 	v->1	
ck Ki	r->1	
ck al	l->1	
ck an	v->1	
ck at	t->12	
ck av	 ->7	
ck ba	k->1	r->1	
ck be	s->1	
ck de	 ->1	n->1	t->4	
ck ef	t->3	
ck ej	 ->1	
ck em	e->1	
ck en	 ->3	
ck et	t->1	
ck fr	u->2	å->5	
ck få	 ->1	
ck fö	r->21	
ck ga	v->1	
ck gr	a->1	
ck gå	r->2	
ck ha	r->4	
ck hu	r->1	
ck hö	r->2	
ck i 	T->1	e->1	f->1	k->1	s->1	u->1	
ck in	 ->1	g->1	l->1	o->1	t->7	
ck ja	g->3	
ck ju	 ->2	
ck ka	n->3	
ck kl	a->1	
ck ko	m->3	
ck kä	n->1	
ck lä	g->1	n->1	
ck me	d->2	
ck mi	s->1	
ck mo	t->2	
ck my	c->2	n->1	
ck må	s->1	
ck mö	j->1	
ck ne	d->1	
ck nu	 ->1	
ck ny	a->1	
ck nå	g->3	
ck oc	h->8	k->2	
ck os	s->2	
ck pa	r->1	
ck på	 ->2	
ck se	 ->1	
ck sk	a->1	y->1	
ck sn	a->1	
ck so	m->3	
ck st	a->1	r->2	
ck sv	å->1	
ck sä	g->1	k->1	r->1	
ck så	 ->15	
ck ti	l->15	
ck tv	u->1	
ck tä	n->1	
ck up	p->1	
ck ut	t->1	
ck va	r->8	
ck vi	 ->1	d->2	k->1	l->4	
ck vä	r->1	
ck än	n->1	
ck är	 ->1	
ck åt	m->2	
ck" -	 ->1	
ck, 1	5->1	
ck, R	e->1	
ck, f	i->1	r->5	
ck, h	e->6	
ck, i	 ->1	n->2	
ck, k	o->3	ä->1	
ck, m	e->2	
ck, n	ä->1	
ck, s	o->2	å->1	
ck, t	r->1	
ck-po	s->1	
ck. M	e->1	
ck.Av	g->1	
ck.De	t->2	
ck.Fr	u->1	
ck.He	r->2	
ck.Ja	g->2	
ck.Ki	n->1	
ck.Ko	m->1	
ck.Äv	e->1	
cka A	h->1	
cka G	r->2	
cka K	a->1	o->1	
cka L	a->1	
cka P	a->1	o->1	
cka S	c->1	
cka a	l->6	t->1	v->1	
cka d	e->7	
cka e	n->2	r->5	
cka f	o->1	r->3	ö->20	
cka h	a->1	e->8	
cka i	 ->3	n->2	
cka k	o->11	
cka l	e->3	
cka m	e->3	i->12	
cka n	y->1	ä->2	
cka o	c->2	r->3	
cka p	a->2	r->1	å->2	
cka r	e->2	å->3	ö->1	
cka s	e->1	i->7	k->2	o->1	
cka t	a->1	i->4	j->1	r->1	
cka u	n->1	p->1	t->3	
cka v	a->7	i->1	o->1	å->5	
cka ä	g->1	v->1	
cka å	t->1	
cka",	 ->1	
cka, 	e->1	o->1	t->1	v->2	
cka.(	I->1	
cka.B	o->1	
cka?"	J->1	
ckad 	a->2	
ckad.	D->1	
ckade	 ->5	s->10	
ckadi	n->1	
ckan 	-->2	d->1	f->1	h->2	i->4	m->1	o->4	p->1	s->3	u->1	v->3	
ckan.	(->1	
ckand	e->21	
ckar 	L->1	a->1	b->1	d->1	e->2	f->6	i->1	k->7	r->2	t->1	u->1	
ckars	 ->1	
ckas 	b->1	e->1	f->1	i->1	k->1	m->10	n->1	o->1	r->1	s->1	u->1	ä->1	å->1	ö->1	
ckas!	H->1	
ckas,	 ->3	
ckas.	J->1	
ckat 	a->1	e->1	k->1	t->1	
ckats	 ->20	.->1	
ckbar	h->4	t->1	
ckbil	d->1	
ckbär	a->1	
ckdel	 ->5	,->1	.->1	e->1	
cke b	i->1	
cke e	n->2	
cke f	r->1	ö->2	
cke i	 ->1	n->1	
cke k	o->1	u->1	
cke l	a->1	i->1	
cke o	f->1	
cke s	e->1	o->1	p->1	
cke t	e->1	i->2	
cke u	t->1	
cke v	a->1	
cke ö	n->1	
cke-a	l->1	v->1	
cke-d	a->1	i->2	
cke-f	o->1	
cke-m	e->1	
cke-s	p->3	t->9	
cke.F	r->1	
cke.H	e->1	
cke.V	i->1	
ckelf	r->2	u->1	
ckeln	 ->3	
ckelp	r->1	
ckelr	o->1	
cken 	a->1	f->2	k->1	m->2	p->7	s->1	t->3	v->1	
cken.	F->1	H->1	
ckens	 ->1	
cker 	C->1	a->31	b->2	d->13	e->1	f->3	g->1	h->3	i->11	j->11	k->2	m->7	o->5	p->1	s->4	t->4	u->1	v->2	ä->2	
cker,	 ->2	
cker.	H->1	
cker:	 ->1	
ckera	n->1	r->2	
ckeri	n->1	
ckert	 ->2	
cket 	a->43	b->16	d->2	e->11	f->15	g->16	h->9	i->12	j->2	k->34	l->25	m->17	n->12	o->25	p->20	r->9	s->72	t->18	u->8	v->73	ä->3	å->2	ö->1	
cket!	(->1	
cket,	 ->22	
cket.	D->1	E->2	M->1	O->1	
cket;	 ->1	
cket?	O->1	
cketm	a->1	
ckfri	t->1	
ckför	e->7	
ckhee	r->14	
ckhet	e->1	
ckhol	m->3	
ckit 	a->1	
ckla 	a->2	d->1	e->9	f->1	h->1	i->1	k->1	l->1	n->3	o->2	r->1	s->4	t->1	u->1	v->1	ö->1	
ckla.	M->1	
cklad	 ->1	e->9	
cklan	d->5	
cklar	 ->3	
cklas	 ->18	.->3	:->1	
cklat	 ->2	,->1	s->3	
ckler	i->4	
cklig	 ->25	,->1	a->14	e->11	h->3	t->52	
cklin	g->175	
ckna 	d->1	s->1	v->1	
cknad	 ->1	e->5	
cknan	d->1	
cknar	 ->2	
cknas	 ->6	
cknat	 ->6	,->1	s->4	
cknes	 ->1	
cknin	g->47	
ckor 	d->2	e->1	f->1	i->5	m->2	n->1	o->3	s->5	t->3	v->1	ä->1	
ckor,	 ->2	
ckor.	B->1	J->1	
ckorn	a->9	
ckors	 ->1	
ckosa	m->1	
ckpro	v->3	
ckra 	f->1	o->2	s->1	v->1	
ckras	t->1	
cks a	n->1	v->3	
cks d	e->1	o->1	
cks e	f->1	
cks i	n->1	
cks m	i->2	
cks n	a->1	
cks o	c->1	
cks p	a->1	
cks r	e->1	
cks s	t->1	
cks t	y->1	
cks u	p->1	t->1	
cks v	a->1	e->1	
cks ö	v->1	
cks.P	å->1	
cks.U	t->1	
cks; 	d->1	
cksam	 ->5	.->1	m->3	
cksbå	d->1	
cksce	n->1	
cksdr	a->3	
cksfa	l->2	
cksil	v->3	
ckskö	r->1	
ckson	 ->2	
cksri	s->2	
cksva	t->1	
ckså 	"->1	-->2	1->1	E->3	F->1	M->1	a->73	b->28	d->25	e->32	f->43	g->18	h->26	i->37	j->1	k->33	l->2	m->38	n->13	o->11	p->18	r->6	s->48	t->31	u->18	v->35	z->1	ä->20	å->3	ö->3	
ckså,	 ->10	
ckså.	D->1	I->1	J->1	N->1	P->1	
cksöd	e->1	
ckt e	r->1	
ckt f	r->1	
ckt h	a->2	
ckt k	a->1	
ckt n	ä->2	
ckt s	i->1	ä->1	å->1	
ckt u	t->1	
ckt v	i->1	
ckt ä	n->1	
ckte 	J->1	a->5	d->2	e->1	i->1	j->1	m->2	o->1	s->1	u->1	v->1	
cktes	 ->5	
ckts 	o->1	u->2	
ckts!	F->1	
ckupa	n->1	t->1	
ckupe	r->3	
ckvid	d->3	
cköns	k->5	
cling	 ->1	
co, e	t->1	
co-af	f->1	
cob S	ö->2	
comba	t->1	
commo	n->1	
compa	s->1	
condi	t->1	
contr	o->2	
copyr	i->1	
coreb	o->1	
corpu	s->4	
corre	c->1	
cost-	b->5	
coup 	d->1	
cours	 ->1	
cover	i->1	
cques	 ->3	
cquis	i->1	
crick	e->1	
ct. D	e->1	
ctnes	s->1	
ctori	t->1	
ctort	a->1	
cu me	d->1	
cu, e	n->1	
cy, s	t->1	
cyavt	a->1	
cycli	n->1	
cydel	 ->1	
cyför	s->1	
cykel	 ->1	,->1	.->1	
cykla	r->4	
cète 	s->1	
d "al	l->1	
d "an	g->1	
d "en	 ->1	
d (ar	t->1	
d (at	t->1	
d (ef	t->1	
d (ko	m->1	
d (rå	d->1	
d - E	U->1	
d - a	t->1	
d - d	ä->1	
d - e	n->1	
d - m	a->1	e->1	
d - o	c->1	
d - u	n->1	
d - v	i->1	
d - Ö	s->1	
d - ä	r->1	
d 12 	m->1	s->1	
d 13 	n->1	s->1	
d 14,	 ->1	
d 164	 ->1	
d 199	5->1	
d 2 i	 ->1	
d 2 m	i->1	
d 2 p	r->1	
d 20 	0->1	
d 200	6->1	
d 24 	p->1	
d 27 	l->1	o->1	
d 28 	n->1	
d 30 	p->1	
d 367	 ->1	
d 5 0	0->1	
d 7 p	å->1	
d 700	 ->1	
d 80 	p->2	
d A. 	G->1	
d Ade	n->1	
d Amo	c->1	
d Ams	t->1	
d BNI	 ->1	
d BSE	 ->1	
d Bal	f->1	
d Bar	a->2	
d Byr	n->2	å->1	
d Cor	b->1	
d Dal	a->1	
d Dav	i->1	
d E-k	o->1	
d EDD	-->1	
d EG-	d->3	
d EU-	l->1	m->1	t->1	
d Eri	k->4	
d Eur	o->17	
d FPÖ	 ->1	
d Fra	n->4	
d GA-	s->1	
d Gen	e->1	
d Gui	g->1	
d Haa	r->1	
d Hai	d->4	
d Ing	l->2	
d Int	e->1	
d Isl	a->1	
d Isr	a->1	
d Jör	g->1	
d Kou	c->3	
d Kul	t->2	
d Kyo	t->1	
d LTC	M->1	
d Lan	d->1	g->3	
d Lea	d->1	
d Lib	a->1	
d Lit	a->1	
d Maa	s->1	
d Mad	r->1	
d Mal	t->1	
d Med	e->1	
d Mid	d->1	
d OLA	F->1	
d Osl	o->1	
d Pad	d->1	
d Pat	t->1	
d Rys	s->1	
d Sav	e->1	
d Sve	r->1	
d Syd	a->1	
d Syr	i->4	
d The	a->1	
d Tib	e->1	
d Tur	k->2	
d USA	 ->2	,->1	:->1	
d Van	d->1	
d Ver	h->1	
d Wid	e->1	
d a) 	a->1	
d acq	u->1	
d adm	i->2	
d all	 ->11	a->18	m->7	t->3	v->2	
d alt	e->1	
d ana	l->1	
d and	a->1	r->17	
d ang	e->1	
d ank	n->1	
d anl	e->5	ä->1	
d ann	a->19	
d ans	e->3	t->5	v->4	å->1	
d ant	a->5	i->1	o->1	
d anv	ä->6	
d arb	e->5	
d arg	u->2	
d art	i->8	
d att	 ->188	
d aut	o->2	
d av 	B->1	E->1	T->1	a->25	b->6	d->36	e->8	f->8	g->1	i->3	j->1	k->4	l->4	m->6	n->5	o->3	p->1	r->3	s->10	t->2	u->3	v->4	
d av.	D->1	
d avf	a->1	
d avs	e->13	i->3	k->1	l->3	
d avt	a->1	
d bak	o->2	
d bal	a->1	
d bar	a->2	
d bas	i->1	
d bed	r->2	ö->2	
d beg	a->1	
d beh	a->3	o->3	å->1	ö->4	
d bek	r->1	v->3	
d ber	i->1	o->1	
d bes	k->2	l->1	t->2	ö->1	
d bet	a->1	r->23	y->3	
d bev	i->4	
d bib	e->2	
d bid	r->3	
d bil	 ->1	,->1	d->2	
d bin	d->1	
d bla	n->1	
d bli	r->3	
d blo	c->1	
d bom	b->2	
d bra	 ->1	,->1	n->1	
d bri	s->3	
d bro	t->1	
d bry	t->1	
d brä	s->1	
d brå	k->1	
d bud	g->1	
d byg	g->2	
d bät	t->1	
d båd	a->1	e->1	
d bör	 ->6	j->1	
d ca.	 ->1	
d cir	k->1	
d dag	e->3	o->5	
d dat	u->1	
d de 	"->1	1->1	a->5	b->4	d->2	f->8	g->3	h->1	i->6	k->4	m->8	n->7	o->6	p->6	r->3	s->9	t->4	v->4	ä->1	å->1	ö->3	
d def	i->1	
d del	 ->2	s->1	t->2	
d dem	 ->8	.->4	o->4	
d den	 ->83	,->1	.->1	n->24	
d der	a->4	
d des	s->29	
d det	 ->52	,->1	t->37	
d dir	e->7	
d dis	k->1	
d dok	u->2	
d dom	s->3	
d dra	m->1	
d dro	g->2	
d dub	b->2	
d dyl	i->1	
d dys	t->1	
d där	 ->7	,->1	e->1	
d då 	d->1	p->1	v->2	
d eff	e->3	
d eft	e->8	
d eko	n->2	
d ele	k->1	
d ell	e->12	
d en 	"->1	a->3	b->8	c->1	d->3	e->11	f->10	g->6	h->3	i->2	j->1	k->3	l->4	m->8	n->5	o->2	p->2	r->6	s->11	t->1	u->1	v->8	ä->1	ö->1	
d ena	 ->1	
d enb	a->2	
d end	a->1	
d ene	r->4	
d enh	e->2	ä->2	
d enl	i->2	
d eno	r->1	
d ent	u->1	
d er 	o->3	r->1	s->4	å->1	
d er.	N->1	P->1	
d era	 ->3	
d erb	j->1	
d ert	,->1	
d ett	 ->42	
d eur	o->5	
d eve	n->1	
d exi	l->1	
d exk	l->1	
d exp	e->3	
d fal	l->1	
d fam	i->1	
d far	a->1	l->2	
d fas	t->1	
d fat	t->2	
d fed	e->2	
d fic	k->1	
d fin	n->5	s->1	
d fle	r->8	x->1	
d fly	g->1	
d fon	d->1	
d for	d->1	m->3	s->1	t->1	
d fra	m->7	n->2	
d fri	 ->1	g->1	h->11	v->1	
d fru	k->1	
d frå	g->14	n->26	
d ful	l->3	
d fun	k->7	n->1	
d fyr	t->1	
d fys	i->1	
d fäl	l->1	
d få 	t->1	
d får	 ->2	
d fåt	t->1	
d föl	j->2	
d för	 ->104	.->2	;->1	b->2	d->6	e->15	h->6	k->1	l->4	n->1	o->2	r->1	s->20	t->1	v->6	ö->1	
d föt	t->1	
d gam	l->1	
d gar	a->1	
d gem	e->6	
d gen	o->5	t->2	
d ger	 ->2	
d gig	a->1	
d gil	t->1	
d gjo	r->2	
d glä	d->2	
d god	 ->1	a->3	k->2	
d got	t->1	
d gra	n->3	
d gru	n->4	p->1	
d grä	n->1	
d grö	n->1	
d gäl	l->60	
d gör	 ->1	a->1	
d ha 	d->1	
d had	e->1	
d hal	v->1	
d ham	n->1	
d han	 ->4	d->5	s->1	t->2	
d har	 ->24	
d hel	t->1	
d hem	l->2	
d hen	n->1	
d hit	t->1	
d hjä	l->26	
d hoc	-->2	
d hon	o->1	
d hos	 ->1	
d hun	d->1	
d hur	 ->4	
d häl	s->1	
d hän	d->2	s->17	v->1	
d här	 ->1	
d häv	d->1	
d hål	l->1	
d hög	 ->2	
d höj	d->1	
d hön	a->1	
d hör	 ->1	t->1	
d i E	U->1	u->3	
d i F	ö->1	
d i L	i->1	
d i M	e->3	
d i S	r->1	
d i a	l->1	r->1	
d i b	e->4	
d i d	a->3	e->12	i->1	
d i e	k->1	n->4	t->4	
d i f	e->1	o->1	r->3	u->1	ö->1	
d i h	a->1	e->1	ä->2	
d i j	u->1	
d i k	a->2	o->2	
d i l	a->1	i->1	
d i m	a->1	e->2	i->1	
d i o	m->1	
d i p	a->1	e->1	r->1	
d i r	a->1	e->1	å->1	
d i s	a->3	t->2	y->2	å->1	
d i t	a->2	v->1	
d i u	n->2	t->2	
d i v	a->1	i->1	å->1	
d i ä	n->1	
d i å	t->1	
d ibl	a->1	
d idé	 ->1	,->1	n->1	
d ifr	å->1	
d imp	u->2	
d in 	n->1	
d inf	i->1	o->7	r->1	ö->1	
d ing	e->2	
d inh	ä->1	
d inn	e->2	
d ino	m->6	
d inr	i->3	
d ins	a->2	p->1	t->4	y->4	
d int	e->23	o->1	r->4	
d inv	ä->1	
d is 	j->2	
d ive	r->1	
d ivä	g->1	
d jag	 ->15	
d jor	d->3	
d jul	i->1	
d jur	i->1	
d jus	t->1	
d jäm	s->3	
d kam	p->1	
d kan	 ->17	o->1	
d kap	i->1	
d kat	a->1	e->1	
d kin	e->1	
d kla	r->1	u->1	
d kli	m->1	
d kna	p->1	
d kol	l->1	
d kom	 ->1	m->48	p->3	
d kon	c->1	f->1	k->10	s->4	t->4	
d kor	r->1	
d kos	t->1	
d kra	f->1	v->5	
d kri	g->1	n->1	s->1	t->1	
d krä	v->1	
d kul	t->3	
d kun	n->1	
d kus	t->1	
d kva	l->8	r->1	
d kvi	n->4	
d kän	n->1	
d kär	n->2	
d köp	s->1	
d lad	e->1	
d lag	e->1	s->1	t->1	
d lan	s->1	
d led	d->1	n->2	
d leg	a->1	
d lig	g->1	
d lik	a->2	n->1	
d lin	d->1	
d liv	s->4	
d lun	c->1	
d läg	g->2	
d läm	n->1	
d län	d->1	
d lät	t->1	
d löp	e->1	
d lös	n->3	
d mai	n->1	
d maj	o->7	
d mak	t->1	
d man	 ->10	,->1	d->1	
d mar	k->3	
d mat	e->1	t->1	
d med	 ->71	b->3	d->2	f->1	l->8	v->1	
d mel	l->8	
d men	 ->1	a->1	
d mer	 ->2	!->1	
d met	o->1	
d mig	 ->3	,->2	
d mik	r->2	
d mil	i->1	j->7	l->1	
d min	 ->11	a->1	i->2	o->5	s->4	u->1	
d mit	t->2	
d mod	e->1	
d mon	o->1	
d mor	a->1	d->1	
d mot	 ->12	s->1	t->1	
d myc	k->9	
d män	n->1	
d mål	 ->1	s->1	
d mån	g->4	
d mås	t->13	
d möj	l->3	
d möt	e->4	
d nam	n->5	
d nat	i->6	u->6	
d naz	i->1	
d neg	a->3	
d ni 	h->1	m->2	s->1	
d ni,	 ->1	
d not	e->1	
d nu 	f->1	s->1	
d num	m->1	
d nuv	a->1	
d nya	 ->1	
d nyf	a->1	
d nyk	t->1	
d nyl	i->2	
d nyp	l->1	
d nyt	t->1	
d näm	n->2	
d när	 ->7	
d näs	t->1	
d någ	o->6	r->5	
d nöd	v->5	
d nöj	e->2	
d nöt	k->1	
d och	 ->100	,->1	
d ock	s->6	
d oer	h->1	
d off	e->1	r->1	
d ojä	m->1	
d oli	k->5	
d om 	a->27	b->2	d->14	e->4	g->1	h->2	i->1	k->1	l->1	m->2	s->4	t->1	u->3	v->3	y->1	
d om.	M->1	
d omb	u->1	
d omf	a->2	
d omr	ö->5	
d oms	o->4	t->1	
d opt	i->1	
d ord	e->1	f->5	
d orm	e->1	
d oro	 ->1	
d oss	 ->5	,->1	.->6	?->1	
d osä	k->1	
d oti	l->1	
d pal	e->2	
d par	l->13	t->2	
d pas	s->1	
d pen	g->3	
d per	 ->1	f->1	s->3	
d pla	n->1	s->1	
d ple	n->1	
d pol	i->8	
d pre	m->1	
d pri	n->6	v->1	
d pro	b->3	d->1	g->3	s->1	
d prö	v->1	
d psy	k->1	
d pub	l->1	
d pun	k->5	
d på 	4->1	7->1	a->5	d->14	e->7	f->1	k->2	l->2	m->3	n->1	o->2	p->1	s->2	t->2	u->1	v->2	ö->1	
d påf	ö->1	
d pål	i->1	
d rad	i->1	
d rea	k->1	
d red	a->1	e->1	
d ref	o->3	
d reg	e->7	i->1	l->1	
d rek	o->1	
d ren	t->1	
d rep	r->2	u->1	
d res	e->1	o->1	p->3	t->2	u->4	
d rev	i->1	
d rik	t->3	
d rol	l->3	
d räd	s->1	
d rät	t->15	
d råd	a->1	e->6	
d rös	t->1	
d röt	t->1	
d s.k	.->1	
d sak	e->3	n->1	
d sam	m->9	o->3	t->3	
d se 	t->2	
d sed	a->6	
d sek	t->2	
d ser	v->1	
d sid	a->8	
d sif	f->1	
d sig	 ->9	
d sin	 ->5	a->6	
d sit	t->3	u->7	
d sju	n->1	
d sjä	l->3	
d sjö	t->1	
d ska	k->1	l->9	m->1	p->1	
d ske	r->1	
d skj	u->1	
d skr	i->1	o->1	
d sku	g->1	l->7	
d sky	l->1	
d sla	k->1	
d slu	t->2	
d slö	s->1	
d smä	r->1	
d små	 ->1	f->2	
d sne	d->2	
d soc	i->7	
d som	 ->138	
d spe	c->2	
d spä	n->3	
d sta	b->1	d->1	l->1	n->1	t->4	
d sti	g->1	
d sto	l->3	r->19	
d str	a->1	i->1	u->5	ö->2	
d sty	r->1	
d stä	n->1	
d stå	 ->1	r->2	
d stö	d->5	r->2	t->2	
d sub	s->3	
d svä	l->1	
d svå	r->1	
d syf	t->3	
d sym	b->1	
d sys	s->8	
d säg	a->4	e->4	
d säk	e->7	r->1	
d säl	l->1	
d sär	s->3	
d så 	a->4	h->1	l->2	m->1	
d så,	 ->1	
d såd	a->7	
d t.e	x->1	
d t.o	.->1	
d ta 	h->1	u->1	
d tac	k->1	
d tag	e->9	i->1	
d tal	a->3	
d tan	k->43	
d tar	 ->1	
d tek	n->1	
d tem	p->1	
d ter	a->1	
d tex	t->1	
d tid	 ->5	,->2	.->1	e->5	i->1	p->1	s->2	t->1	
d til	l->94	
d tjä	n->1	
d tol	v->1	
d ton	v->1	
d top	p->2	
d tra	n->5	
d tre	 ->3	d->3	
d tro	 ->1	r->1	
d tun	n->1	
d tur	i->1	
d tvi	v->1	
d två	 ->7	
d typ	f->1	
d täc	k->1	
d tän	k->2	
d tät	a->1	
d und	a->2	e->8	
d ung	d->1	
d uni	o->2	
d upp	d->2	f->3	m->5	n->1	r->3	s->1	
d urs	k->1	ä->1	
d urv	a->1	
d uta	n->2	r->9	
d utb	e->2	i->2	
d utf	o->1	
d utg	å->2	
d utn	y->1	
d uts	k->6	l->2	
d utv	e->4	i->5	ä->2	
d vac	k->1	
d vad	 ->7	
d val	e->2	u->1	
d van	 ->1	
d var	 ->6	a->3	f->1	i->1	j->3	s->2	
d ver	k->5	s->2	
d vet	e->8	
d vi 	a->1	b->1	d->2	e->2	f->2	g->1	h->3	i->1	j->1	k->2	l->1	m->2	n->1	s->7	t->2	u->1	v->4	
d vid	 ->4	
d vik	t->2	
d vil	j->3	k->5	l->7	
d vis	a->4	s->7	
d vit	b->2	
d von	 ->1	
d väl	 ->1	
d vär	d->1	
d vår	 ->5	a->9	t->8	
d yrk	a->1	e->2	
d ytt	e->5	
d ÖVP	 ->1	
d Öst	e->1	
d än 	d->2	i->1	k->1	m->1	
d änd	a->1	r->4	å->1	
d änn	u->2	
d är 	E->3	a->3	d->14	e->5	f->3	g->1	i->2	k->3	l->2	m->2	n->1	o->1	s->1	t->1	v->4	
d äre	n->2	
d äve	n->2	
d år 	2->1	
d åre	n->1	t->1	
d årt	u->1	
d åt 	a->1	f->1	i->1	t->1	
d åta	g->1	l->2	
d åte	r->3	
d åtg	ä->3	
d öka	t->1	
d ökn	i->1	
d öms	e->1	
d öpp	e->1	n->1	
d öst	e->1	
d öve	r->31	
d övr	i->2	
d! Li	k->1	
d! Ni	 ->1	
d) i 	ä->1	
d), o	c->1	
d), r	å->1	
d), s	o->1	
d, "a	f->1	
d, 56	 ->1	
d, Da	n->1	
d, EC	H->1	
d, Fi	n->1	
d, It	a->2	
d, No	r->1	
d, Sp	a->2	
d, am	b->1	
d, at	t->5	
d, bl	i->1	
d, bo	r->1	
d, bö	r->1	
d, de	 ->1	n->1	s->1	t->2	
d, dv	s->1	
d, dä	r->5	
d, då	 ->2	
d, ef	t->3	
d, ek	o->1	
d, en	 ->4	
d, et	t->1	
d, fa	k->1	
d, fr	i->1	
d, fö	r->5	
d, gö	r->1	
d, ha	f->1	r->3	
d, he	r->2	
d, hu	r->1	
d, hy	g->1	r->1	
d, i 	s->2	
d, in	f->1	n->1	
d, ka	n->1	
d, ko	m->1	
d, kr	ä->1	
d, lä	n->1	
d, ma	n->1	
d, me	d->3	n->14	
d, mi	l->1	n->1	
d, nä	m->2	
d, nå	g->1	
d, oc	h->23	k->2	
d, om	 ->4	
d, pl	u->1	
d, pr	a->1	
d, på	 ->1	
d, re	v->1	
d, rä	t->1	
d, sa	m->1	
d, sk	a->1	u->1	
d, so	c->2	m->8	
d, sp	a->1	e->1	
d, st	a->1	r->1	
d, sä	r->1	
d, så	 ->3	v->1	
d, ti	l->1	
d, to	t->1	
d, tr	o->2	
d, ty	d->1	
d, un	d->2	
d, up	p->1	
d, ut	n->1	
d, va	r->3	
d, vi	d->2	l->4	
d, är	 ->2	
d, äv	e->1	
d- (P	T->1	
d-aff	ä->1	
d-för	k->1	
d-kos	t->1	
d. Vi	 ->1	
d. Ös	t->1	
d. ös	t->1	
d."Ja	g->1	
d."Me	d->1	
d.(Sa	m->1	
d., f	r->1	
d.- (	P->1	
d.. (	F->1	
d..(D	E->1	
d.All	t->1	
d.And	r->1	
d.Att	 ->2	
d.Bed	ö->1	
d.De 	b->1	e->1	f->1	k->1	
d.Den	 ->6	n->2	
d.Des	s->1	
d.Det	 ->30	t->6	
d.Dir	e->2	
d.Där	e->1	f->2	
d.Då 	f->1	
d.Eff	e->1	
d.Eme	l->1	
d.En 	b->1	
d.Eur	o->3	
d.Fak	t->1	
d.Frå	g->2	
d.För	 ->5	
d.Gen	o->1	
d.Had	e->1	
d.Han	 ->1	
d.Her	r->13	
d.Hur	 ->1	
d.I T	i->1	
d.I d	e->1	
d.I k	l->1	
d.I s	t->2	
d.I v	i->1	
d.Inf	ö->1	
d.Ini	t->1	
d.Inn	e->1	
d.Irl	a->1	
d.Jag	 ->23	
d.Kan	 ->1	
d.Kom	 ->1	m->4	
d.Kon	s->1	
d.Låt	 ->2	
d.Man	 ->1	
d.Men	 ->7	t->1	
d.Mit	t->1	
d.Mot	 ->1	
d.Män	n->1	
d.Mån	g->1	
d.Nat	u->1	
d.Ni 	h->1	m->1	
d.Nu 	h->1	ä->1	
d.När	 ->2	
d.Om 	S->1	d->2	
d.Omr	ö->14	
d.Ord	e->1	
d.Par	l->1	
d.På 	s->1	
d.Reg	e->3	
d.Sav	e->1	
d.Som	 ->2	
d.Sub	v->1	
d.Så 	ä->1	
d.Tac	k->1	
d.Til	l->1	
d.Tro	t->1	
d.Und	e->1	
d.Upp	e->1	
d.Uta	n->1	
d.Utg	i->1	
d.Vad	 ->1	
d.Var	 ->1	
d.Vet	e->1	
d.Vi 	e->1	f->1	h->3	k->2	m->2	t->1	ä->1	
d.Vil	k->1	
d.Vis	s->1	
d.Änd	r->1	
d.Äve	n->1	
d.Å a	n->2	
d.År 	1->1	
d: "D	e->1	
d: "O	m->1	
d: de	l->1	
d: en	 ->1	
d; de	t->3	
d; in	s->1	t->1	
d? Ha	r->1	
d?- (	P->2	
d?. (	E->1	
d?Där	 ->1	
d?För	 ->1	
d?Her	r->1	
d?Jag	 ->1	
d?Vi 	h->1	
d?Är 	d->1	
da - 	ä->1	
da 12	5->1	
da 20	0->1	
da 60	 ->1	
da Co	s->5	
da EU	 ->1	-->1	
da Er	i->1	
da Eu	r->3	
da Fe	i->1	
da Go	l->1	
da ag	e->2	
da ak	t->1	
da al	l->6	
da an	a->1	l->1	p->1	s->1	t->1	
da ar	b->6	
da at	t->26	
da av	 ->8	,->1	s->3	t->1	
da ba	r->2	
da be	g->1	h->1	k->2	s->1	t->1	v->1	
da bi	l->2	
da bo	t->2	
da bå	d->1	
da ch	a->2	
da ci	v->1	
da de	 ->11	b->1	l->1	m->3	n->16	r->1	s->3	t->14	
da di	s->2	
da dj	u->2	
da do	k->2	m->3	
da dr	i->1	
da ef	f->1	t->1	
da ek	o->2	
da el	i->1	l->4	
da en	 ->18	g->1	
da er	 ->2	
da et	t->7	
da eu	r->3	
da ex	e->1	
da fa	l->3	
da fi	l->1	n->1	s->1	
da fo	l->2	n->1	r->1	
da fr	a->4	å->3	
da fö	l->2	r->41	
da ga	r->1	
da ge	m->2	
da gi	f->1	
da gr	u->2	ä->1	
da gä	l->1	
da gö	r->1	
da ha	n->2	r->3	
da hi	s->1	
da hu	m->1	r->1	
da hy	p->1	
da hä	n->2	
da hö	g->1	
da i 	K->1	L->1	d->3	f->3	k->8	n->1	s->1	v->1	
da id	é->1	
da ig	e->2	
da in	 ->5	d->2	f->1	o->1	s->3	t->5	
da ja	g->2	
da jo	r->2	
da ka	m->1	p->1	
da ko	l->1	m->5	n->7	r->1	
da kr	a->2	e->1	
da ku	s->1	
da kv	a->1	
da kä	r->1	
da la	b->1	g->1	n->2	
da le	d->1	
da li	v->1	
da lo	k->1	v->1	
da lu	c->1	
da lä	n->4	
da lö	n->1	
da ma	n->1	r->1	t->1	
da me	d->22	
da mi	l->5	t->1	
da mo	t->4	
da my	c->2	
da mä	n->1	t->1	
da må	l->3	
da mö	j->2	r->1	
da na	t->1	
da ne	d->1	
da ni	 ->2	
da ny	a->1	h->1	
da nä	r->1	
da nå	g->3	
da nö	j->1	t->1	
da oc	h->14	
da od	u->1	
da ol	j->1	
da om	 ->4	r->2	
da or	d->2	g->1	
da os	s->6	
da pa	r->7	t->1	
da pe	n->2	r->3	
da ph	t->1	
da pl	a->3	
da po	l->4	s->1	
da pr	o->7	
da pu	n->1	
da på	 ->4	,->1	
da ra	m->1	
da re	f->1	g->5	k->3	p->2	s->6	
da ri	s->2	
da ry	g->1	
da rä	t->3	
da rå	d->1	
da rö	s->3	
da sa	m->2	
da sc	e->1	
da se	d->3	k->1	t->1	
da si	d->3	g->11	m->1	n->4	t->1	
da sk	a->2	e->1	o->2	u->1	y->1	ä->1	
da sm	å->1	
da so	m->15	
da st	a->5	o->1	r->2	ä->1	ö->1	
da su	b->1	m->1	
da sy	f->1	
da sä	k->1	n->3	t->4	
da ta	n->1	
da te	n->1	
da ti	d->1	l->38	n->1	o->1	
da to	t->1	
da tr	a->3	ä->1	å->2	
da tu	n->1	
da tå	g->1	
da un	d->3	i->1	
da up	p->3	
da ur	 ->1	
da ut	 ->3	:->1	b->1	s->1	t->2	
da va	r->1	t->1	
da ve	r->2	
da vi	 ->2	c->1	d->2	l->5	
da vä	g->1	v->1	
da vå	l->1	r->1	
da än	d->3	
da är	 ->3	e->1	
da åt	a->4	g->4	
da öa	r->1	
da ör	e->1	
da öv	e->2	
da!De	n->1	
da" b	i->1	
da, J	a->1	
da, b	l->1	
da, d	ä->1	
da, e	f->1	x->1	
da, f	r->1	å->1	ö->3	
da, h	a->1	u->1	
da, i	 ->1	n->1	
da, k	o->1	
da, m	e->3	
da, n	ä->1	
da, o	c->1	m->2	
da, p	å->1	
da, r	e->1	ä->1	
da, s	e->1	k->1	o->4	ä->1	å->1	
da, t	y->1	
da, v	i->3	ä->1	
da, ä	r->1	
da. E	n->1	
da.Be	r->1	
da.De	s->1	t->4	
da.Då	 ->1	
da.Et	t->1	
da.Fr	u->2	
da.Fö	r->1	
da.Ha	n->1	
da.He	r->4	
da.I 	v->1	
da.Ib	l->1	
da.Ja	g->3	
da.Kä	r->1	
da.Me	n->2	
da.Mi	n->1	
da.Ni	 ->1	
da.Nä	r->1	
da.Oc	h->2	
da.Ru	m->1	
da.Va	d->1	
da.Vi	 ->3	d->1	
da.Är	 ->1	
da.Äv	e->1	
da?De	t->2	
da?Fr	u->1	
da?In	i->1	
daboc	k->2	
dac b	l->1	ö->1	
dac o	s->1	
dac",	 ->1	
dac-s	y->1	
dad a	v->1	
dad b	e->1	
dad i	 ->1	
dad p	å->3	
dad r	ä->1	
dad s	t->1	
dad.S	u->1	
dade 	H->2	f->1	h->1	i->3	k->1	o->2	p->5	s->5	t->1	v->2	
dade,	 ->1	
dade.	E->1	
dades	 ->2	,->1	.->3	
dafon	e->1	
dafri	k->2	
dag -	 ->3	
dag I	N->1	
dag a	l->1	n->2	t->5	v->3	
dag b	e->1	
dag d	e->2	r->1	ö->1	
dag e	m->1	n->3	t->1	
dag f	i->1	o->2	r->1	å->1	ö->10	
dag g	a->1	r->1	ä->1	
dag h	a->15	i->1	o->1	u->1	ä->2	ö->1	
dag i	 ->7	n->8	
dag j	u->1	
dag k	a->2	l->2	o->2	
dag l	a->1	ä->2	ö->1	
dag m	e->4	å->4	
dag n	o->1	ä->1	
dag o	c->7	m->2	
dag p	å->3	
dag r	e->1	i->1	å->1	ö->1	
dag s	a->1	e->1	k->1	o->5	t->2	
dag t	a->4	i->3	o->1	r->2	y->1	ä->1	
dag u	p->2	t->2	
dag v	a->2	i->2	ä->2	
dag Ö	s->1	
dag ä	g->1	n->1	r->14	
dag, 	a->3	b->2	d->2	e->3	f->3	h->1	i->1	l->1	m->2	n->1	o->2	p->1	s->3	t->2	v->2	ä->3	
dag. 	P->1	
dag.(	A->1	
dag.A	n->1	r->1	
dag.D	e->9	
dag.E	r->1	
dag.F	r->1	ö->1	
dag.G	e->1	
dag.H	e->1	u->1	y->1	
dag.I	 ->2	
dag.J	a->7	
dag.K	a->1	
dag.L	i->1	
dag.O	m->1	
dag.V	i->1	
dag: 	d->1	
dag:D	e->1	
dagar	 ->8	.->1	n->6	s->2	
dagas	k->1	
dagen	 ->8	,->1	.->3	s->24	
dagli	g->8	
dagog	i->1	
dagor	d->52	
dags 	a->8	d->1	f->5	m->1	o->2	
dags,	 ->2	
dags.	F->1	
dagsb	o->1	
dagsl	ä->2	
dagst	i->2	
dahål	l->43	
daire	.->1	
dakis	 ->2	b->1	
dakti	o->1	
daktö	r->2	
dal!H	ä->1	
dal, 	s->1	
dalag	 ->3	,->1	
dalan	k->1	
daler	 ->2	n->3	
dalyd	e->2	
dalös	a->1	
dam -	 ->1	
dam 1	9->1	
dam i	n->1	
dam o	c->1	
dam p	å->1	
dam s	k->1	o->1	
dam t	i->1	
dam v	a->1	
dam ä	r->1	
dam, 	a->1	b->1	v->1	
dam.N	ä->1	
damaf	f->1	
damen	t->1	
damer	 ->41	i->4	
damfö	r->27	
damm 	a->1	
damma	r->3	
damot	 ->25	!->7	,->16	e->26	
damre	s->1	
damål	 ->1	,->2	.->2	e->6	s->2	
damöt	e->84	
dan -	 ->1	
dan 1	9->15	
dan 4	 ->1	
dan A	m->1	
dan E	M->1	
dan F	l->1	
dan P	l->1	
dan S	h->1	
dan a	l->2	n->9	r->2	t->2	v->9	
dan b	e->9	l->1	o->1	r->1	ä->1	ö->3	
dan d	a->1	e->25	i->2	o->1	å->1	
dan e	f->2	n->12	r->1	t->3	x->2	
dan f	a->1	e->1	i->5	l->4	o->3	r->4	å->1	ö->13	
dan g	a->2	e->3	j->1	o->1	å->1	ö->2	
dan h	a->47	ä->3	
dan i	 ->16	n->9	s->1	
dan j	a->3	u->1	
dan k	a->6	o->6	v->2	y->1	
dan l	a->1	e->1	i->2	y->1	ä->1	å->1	
dan m	a->2	e->3	o->1	y->4	å->4	
dan n	u->4	y->1	ä->2	å->3	ö->1	
dan o	c->5	f->1	m->5	r->1	v->1	
dan p	o->2	r->1	å->8	
dan r	a->1	e->4	o->1	u->1	ö->1	
dan s	a->8	i->3	k->11	o->1	t->2	
dan t	a->11	e->1	i->8	y->1	
dan u	n->2	p->2	r->1	t->5	
dan v	a->2	e->4	i->11	ä->2	
dan ä	g->2	n->1	r->9	
dan å	r->1	
dan ö	k->1	v->2	
dan, 	f->1	g->1	h->1	i->1	j->1	k->1	m->2	n->2	o->1	s->3	u->1	v->2	
dan.A	l->1	
dan.D	e->7	ä->1	
dan.H	e->1	
dan.I	 ->1	
dan.J	a->5	
dan.S	k->1	o->1	
dan? 	2->1	
dan?H	u->1	
dan?S	e->1	
dana 	-->2	a->2	b->4	d->4	e->1	f->9	g->1	h->4	i->1	l->1	m->1	o->2	p->3	r->5	s->8	t->1	v->1	å->2	
danan	d->1	
danbe	r->2	
dande	 ->82	,->3	.->6	n->1	t->13	
dandr	a->1	
danfl	y->1	
dange	l->1	
danhå	l->1	
danie	n->1	
danma	n->1	
danor	d->1	
danrö	j->6	
dans 	v->1	
dansk	 ->2	a->23	
dansv	a->7	
dant 	-->1	E->2	a->2	b->3	c->1	f->9	i->2	k->4	m->1	n->2	o->2	p->2	s->18	t->1	u->2	ä->1	
dant,	 ->1	
danta	 ->1	g->36	s->2	
dapes	t->1	
dar a	l->2	t->7	
dar b	e->1	
dar d	e->5	ä->1	
dar e	l->1	n->1	
dar g	e->1	
dar h	a->1	
dar i	 ->1	h->1	n->1	
dar j	u->1	
dar m	e->3	i->1	ä->1	
dar n	i->1	
dar o	s->1	
dar r	e->3	
dar s	i->2	o->2	
dar, 	k->1	u->1	
dar.D	e->1	
dar.J	a->1	
darbe	t->2	
dard 	f->1	o->1	p->1	s->2	v->1	
dard,	 ->2	
dard.	D->1	
dard;	 ->1	
darde	n->3	r->2	
dardi	s->9	
dare 	D->1	a->5	b->3	d->3	e->1	f->25	h->2	i->3	k->3	l->1	m->4	n->1	o->5	p->6	s->5	t->8	u->5	v->2	ä->2	
dare,	 ->8	
dare.	A->1	B->1	D->2	J->3	M->1	V->1	
dare?	D->1	O->1	
dareb	e->3	
daren	 ->5	
dares	 ->3	,->1	
dareu	t->4	
darfö	r->1	
daris	k->2	
darit	e->29	
darna	 ->19	.->1	s->3	
dars 	d->1	
darsk	a->2	
darsy	d->1	
das a	v->2	
das d	e->1	
das f	ö->2	
das g	e->1	
das i	 ->4	n->3	
das m	e->2	
das n	u->1	
das o	c->1	
das p	o->1	å->9	
das r	ä->1	
das s	o->1	
das t	a->1	i->4	
das u	t->3	
das ö	v->1	
das, 	f->1	m->1	s->1	u->1	å->1	
das.A	l->1	
das.B	l->1	
das.D	e->2	ä->1	
das.H	e->2	
das.I	 ->2	n->1	
das.M	e->1	
das.T	i->1	
das.V	i->1	
das.Å	t->1	
das?H	a->1	
dast 	1->1	2->1	5->1	7->1	9->1	a->2	b->2	d->5	e->9	f->6	g->4	i->7	k->5	l->1	m->6	n->3	o->5	p->4	r->2	s->4	t->6	u->2	ä->4	å->1	ö->1	
dast.	E->1	
daste	 ->1	
dat a	t->5	v->1	
dat b	e->1	
dat d	e->1	
dat f	o->1	r->2	ö->1	
dat h	i->1	
dat k	o->1	
dat m	å->1	
dat n	å->1	
dat p	å->4	
dat s	i->1	o->1	å->1	
dat u	p->1	
dat, 	b->1	m->2	s->1	
dat.F	ö->1	
dat.T	a->1	
data 	o->1	
data,	 ->1	
datab	a->1	
datas	ä->1	
daten	 ->1	
dater	 ->2	a->2	i->1	n->1	
datet	 ->3	.->1	
datio	n->33	
datla	n->1	
datli	s->1	
datlä	n->10	
dato 	ö->1	
dator	b->1	s->1	
datpe	r->9	
dats 	a->1	i->2	o->1	
dats,	 ->2	
dats.	R->1	S->1	
datum	 ->8	,->2	.->1	e->2	
dbar 	s->1	
dbara	 ->3	
dbart	 ->4	,->1	
dbedd	 ->1	
dbelä	g->1	
dbesl	u->16	
dbest	ä->1	
dbetä	n->1	
dborg	a->167	e->3	
dbrot	t->1	
dbruk	 ->6	,->2	a->13	e->13	s->22	
dbrän	d->1	
dbult	e->1	
dbävn	i->10	
dd at	t->17	
dd av	 ->4	s->1	
dd ba	k->1	
dd bö	r->1	
dd el	l->1	
dd fö	r->18	
dd hä	r->1	
dd i 	l->1	
dd in	o->1	
dd me	d->1	
dd mo	d->1	t->2	
dd må	s->1	
dd oc	h->4	
dd sa	m->2	
dd so	m->1	
dd st	å->1	
dd ti	l->3	
dd ut	a->1	v->1	
dd vi	d->2	
dd än	 ->1	n->1	
dd öv	e->1	
dd), 	s->1	
dd, d	e->1	
dd, e	k->1	
dd, h	e->1	
dd, v	i->1	
dd.De	t->2	
dd.Ja	g->2	
dd.Me	n->1	
dd.Na	t->1	
dd.Re	g->1	
dd.Vi	 ->1	
dda 6	0->1	
dda a	l->1	r->1	t->13	v->1	
dda c	i->1	
dda d	e->5	j->1	
dda e	l->1	
dda f	ö->2	
dda g	e->2	r->1	
dda i	 ->2	
dda k	a->1	o->1	r->1	
dda l	e->1	ö->1	
dda m	a->1	e->1	i->3	ä->1	
dda o	l->1	
dda p	l->1	
dda r	e->2	ä->2	
dda s	i->4	k->1	
dda t	i->1	
dda u	p->1	t->1	
dda v	å->1	
dda. 	E->1	
dda.M	e->1	
ddad 	b->1	
ddade	 ->4	s->1	
ddag 	a->1	k->1	m->1	o->1	
ddag,	 ->2	
ddag.	D->1	
ddage	n->2	
ddags	 ->2	,->1	b->1	
ddand	e->1	
ddar 	r->1	
ddare	,->1	
ddars	y->1	
ddas.	D->1	I->1	
ddats	.->1	
dde "	a->1	
dde 4	1->1	
dde A	m->2	
dde V	e->1	
dde a	t->2	
dde d	e->2	o->1	ä->1	
dde e	r->1	
dde f	r->3	ö->2	
dde i	 ->6	
dde j	a->1	
dde m	i->1	
dde p	å->4	
dde t	i->7	
dde v	å->1	
dde, 	j->1	
ddel 	a->1	
ddela	 ->10	d->2	n->41	r->1	t->5	
ddele	n->2	
ddelh	o->1	
dden 	a->1	h->1	
dden,	 ->1	
dder 	t->1	
ddes 	1->1	a->1	d->1	i->3	m->1	u->3	
ddes.	R->1	
ddet 	a->12	i->1	m->1	o->1	ö->1	
ddet,	 ->2	
ddhis	t->1	
ddigh	e->1	
ddigt	 ->1	
dding	t->2	
dditi	o->1	
ddnin	g->4	
dds e	m->1	
ddsme	d->4	
ddsni	v->6	
ddsom	r->1	
ddsor	g->1	
ddspr	o->1	
ddsst	ö->1	
ddssä	l->1	
ddstu	l->1	
de "a	l->1	v->1	
de "d	e->1	
de "f	ö->1	
de "k	o->2	
de "l	ä->2	
de "s	v->1	
de (A	5->29	
de (m	a->1	
de - 	a->1	d->3	e->1	f->2	h->1	j->2	o->2	p->1	s->4	t->1	u->1	ä->1	
de 11	 ->1	
de 12	 ->1	
de 14	 ->3	
de 15	 ->1	
de 18	 ->1	
de 19	9->3	
de 20	 ->1	
de 25	 ->4	
de 26	 ->1	
de 40	 ->1	
de 41	 ->1	
de 8 	t->1	
de 9 	m->1	
de Ah	e->1	
de Al	t->2	
de Am	s->2	
de B 	t->1	
de Bu	s->1	
de Ce	n->2	
de Da	n->1	
de Du	i->1	
de EU	-->1	
de Eu	r->7	
de Fr	a->1	
de Ga	m->1	r->2	
de Gr	a->2	
de Ha	i->1	
de He	d->1	
de Ho	l->1	
de Im	b->1	
de Ir	l->1	
de Ja	c->1	
de Ka	r->2	
de Ki	n->1	
de Ko	c->2	u->1	
de La	n->1	
de Lo	y->1	
de Ma	r->4	
de Me	l->1	
de Na	p->1	t->1	
de OL	A->1	
de Oi	l->1	
de Pa	l->6	
de Pr	o->14	
de Ra	p->1	
de Ro	m->2	
de Sa	n->1	
de Sc	h->2	
de Se	i->1	
de Sv	e->1	
de Sw	o->1	
de Tr	i->1	
de Tu	r->1	
de Va	t->1	
de Ve	n->1	
de We	b->1	
de ab	s->1	
de ad	j->1	m->5	
de af	f->1	
de ag	e->2	
de ai	d->1	
de ak	t->5	
de al	b->2	l->24	
de am	b->1	e->3	
de an	a->2	b->1	d->9	f->1	g->5	l->2	m->4	o->1	s->27	t->6	v->2	
de ap	p->2	
de ar	a->3	b->15	g->1	t->1	
de as	p->1	y->1	
de at	t->69	
de av	 ->162	.->1	d->1	f->3	g->4	s->1	t->4	v->1	
de ba	k->1	n->3	r->5	s->2	
de be	d->2	f->6	g->6	h->10	k->1	l->3	r->7	s->20	t->24	v->4	
de bi	d->3	l->14	o->1	
de bl	a->3	i->5	
de bo	r->2	
de br	a->1	e->1	i->7	o->6	ä->1	
de bu	d->2	
de by	g->2	r->3	t->1	
de bä	s->4	t->1	
de bå	d->6	t->3	
de bö	r->3	
de ce	n->3	
de ch	a->1	
de da	g->4	m->3	n->2	t->1	
de de	 ->13	b->4	c->2	l->11	m->5	n->40	p->1	s->2	t->29	
de di	a->1	p->1	r->7	s->6	t->1	
de dj	ä->1	
de do	c->2	g->1	m->2	
de dr	a->11	o->1	y->1	
de dä	r->12	
de då	 ->3	.->1	
de dö	r->1	
de ef	f->2	t->9	
de eg	e->3	n->2	
de ej	 ->1	
de ek	o->22	
de el	e->3	l->5	m->1	
de em	o->2	
de en	 ->24	d->8	e->2	g->1	h->1	l->2	o->4	s->9	t->1	
de ep	o->1	
de er	 ->1	b->1	k->1	
de et	a->1	n->2	t->13	
de eu	r->55	
de ev	e->1	
de ex	a->3	p->16	t->2	
de fa	c->2	k->7	l->6	m->3	n->1	r->11	s->2	t->3	x->1	
de fe	l->1	m->8	
de fi	c->2	l->1	n->15	s->4	
de fj	o->3	
de fl	a->4	e->23	y->2	
de fo	l->2	n->1	r->11	
de fr	a->25	e->4	i->9	u->4	ä->5	å->52	
de fu	n->5	t->1	
de fy	r->8	
de fä	s->1	
de få	 ->8	r->6	t->3	
de fö	l->2	r->177	
de ga	m->6	n->1	r->3	v->2	
de ge	 ->2	m->7	n->11	o->1	r->2	
de gi	l->1	
de gj	o->3	
de gl	ö->1	
de go	d->9	t->1	
de gr	a->2	u->22	ä->5	å->1	ö->2	
de gä	l->2	
de gå	n->4	r->1	
de gö	r->5	
de ha	 ->11	d->3	f->1	n->12	r->40	
de he	l->5	m->5	r->2	t->1	
de hi	e->1	n->3	s->2	t->2	
de hj	ä->1	
de ho	n->1	p->1	r->1	s->2	t->2	
de hu	r->1	v->1	
de hy	c->1	s->1	
de hä	n->3	r->15	
de hå	l->3	r->2	
de hö	g->5	j->1	r->1	
de i 	A->1	E->5	F->1	H->1	I->1	K->1	S->1	a->4	b->3	d->20	e->5	f->9	g->5	h->4	k->9	l->2	m->3	n->3	o->1	p->2	r->3	s->17	t->1	u->8	v->1	y->2	z->1	Ö->2	ä->1	
de ic	k->8	
de id	e->1	é->2	
de if	r->1	
de ig	e->1	
de in	b->4	d->4	f->7	g->11	i->3	l->6	n->10	o->4	r->6	s->16	t->59	v->6	
de is	r->3	
de it	a->5	
de ja	g->17	
de jo	r->3	u->1	
de ju	 ->1	d->1	r->1	s->2	
de jä	m->1	
de ka	m->1	n->29	p->2	r->1	t->9	
de ke	m->1	
de ki	n->5	
de kl	a->3	i->1	
de kn	a->2	
de ko	l->12	m->67	n->26	s->8	
de kr	a->8	i->6	y->1	ä->3	
de ku	l->2	n->29	s->2	
de kv	a->7	ä->1	
de kä	l->1	n->1	r->1	
de la	 ->1	g->9	n->2	s->1	
de le	d->8	g->1	v->3	
de li	b->4	d->2	g->3	n->1	v->3	
de lo	g->3	k->7	
de ly	c->1	s->1	
de lä	c->1	g->4	m->1	n->8	t->1	
de lå	n->3	t->1	
de lö	f->1	
de ma	j->6	k->6	n->11	r->6	x->1	
de me	d->59	k->2	l->3	n->2	r->2	s->20	t->2	
de mi	g->4	l->11	n->11	s->6	t->1	
de mo	d->1	n->1	t->6	
de mu	l->4	
de my	c->14	l->1	n->3	
de mä	k->2	n->33	r->3	
de må	l->16	n->15	s->15	
de mö	j->4	r->1	
de na	t->49	
de ne	d->1	g->2	
de ni	 ->3	o->2	v->1	
de no	r->9	
de nu	 ->3	v->7	
de ny	a->20	h->2	l->1	s->4	t->1	
de nä	m->2	r->19	t->1	
de nå	g->7	
de nö	d->3	
de ob	e->3	
de oc	h->106	k->15	
de oe	r->1	
de of	a->1	f->9	t->1	
de ol	a->1	i->41	j->1	y->6	
de om	 ->65	,->3	e->1	f->4	k->1	r->28	s->3	
de on	s->2	
de op	e->1	i->1	
de or	d->10	g->6	k->1	o->3	s->3	
de os	s->5	
de ot	i->1	
de ov	a->1	i->1	ä->1	
de pa	l->2	r->24	
de pe	k->2	l->1	n->3	r->22	
de pl	a->4	i->1	
de po	l->29	p->1	r->2	s->3	t->1	
de pr	a->3	e->4	i->22	o->37	
de pu	b->1	n->7	
de på	 ->50	b->2	g->3	p->3	s->1	
de ra	d->1	m->2	p->4	s->1	
de re	a->2	d->6	f->15	g->54	k->1	l->1	n->3	s->17	v->3	
de ri	k->18	s->3	
de ro	l->7	
de ru	b->1	n->1	t->1	
de rä	k->2	t->39	
de rå	d->8	
de rö	r->1	s->1	
de sa	g->2	k->2	m->18	n->2	
de se	d->4	k->2	n->33	s->1	t->2	x->3	
de si	f->2	g->12	n->1	s->2	t->9	
de sj	u->1	ä->3	
de sk	a->26	e->1	i->1	j->3	o->2	r->2	u->9	y->2	ä->2	
de sl	a->1	u->3	
de sm	å->21	
de sn	a->2	
de so	c->10	m->91	r->1	
de sp	a->1	e->3	
de st	a->20	e->2	i->1	o->24	r->15	y->3	ä->5	å->4	ö->18	
de su	m->1	n->1	v->1	
de sv	a->6	å->6	
de sy	f->4	m->1	n->3	r->1	s->17	
de sä	g->4	k->7	m->4	n->1	t->11	
de så	 ->5	d->1	r->1	
de t.	o->1	
de ta	 ->1	g->1	l->13	n->4	r->2	x->2	
de te	k->3	r->1	x->3	
de ti	d->16	l->68	o->1	s->1	t->1	
de tj	ä->8	
de to	g->1	t->2	
de tr	a->7	e->11	o->2	ä->2	
de tu	n->1	r->1	s->1	
de tv	e->1	i->3	å->19	
de ty	d->2	s->2	
de tä	n->1	
de ul	t->1	
de un	d->16	i->1	
de up	p->23	
de ur	a->4	b->1	
de ut	a->9	b->4	g->5	k->1	l->2	m->2	o->1	r->1	s->2	t->12	v->15	ö->2	
de va	d->4	l->4	n->2	r->27	t->3	
de ve	c->3	l->1	r->15	t->12	
de vi	 ->23	d->5	k->20	l->9	r->1	s->6	t->1	
de vo	l->1	n->2	
de vr	a->1	
de vä	g->1	l->4	n->5	r->8	s->1	
de vå	r->4	
de yr	k->3	
de yt	t->11	
de Ös	t->1	
de äg	t->1	
de äl	d->1	
de äm	n->1	
de än	 ->2	d->13	n->3	
de är	 ->50	.->1	e->2	
de äv	e->2	
de å 	r->1	
de år	 ->7	.->1	e->10	h->1	
de ås	i->3	t->1	
de åt	 ->2	a->8	e->6	g->37	t->1	
de öa	r->1	
de ök	n->1	
de öm	m->1	
de ön	s->4	
de öp	p->3	
de ös	t->3	
de öv	e->20	n->1	r->12	
de! J	a->5	
de! N	i->1	
de!Al	l->1	
de!Ja	g->1	
de!Ni	 ->1	
de", 	o->1	
de(A5	-->1	
de, ,	 ->1	
de, D	i->1	
de, E	r->1	
de, F	r->1	
de, G	r->1	
de, L	e->1	
de, a	t->8	v->1	
de, b	e->1	o->3	y->1	ö->1	
de, d	e->7	v->1	ä->1	å->1	
de, e	f->4	m->1	n->1	
de, f	r->4	ö->5	
de, h	a->2	e->6	u->2	
de, i	 ->6	n->8	
de, j	a->2	
de, k	a->2	i->1	o->4	
de, l	i->1	
de, m	e->10	i->1	o->1	å->1	
de, n	a->2	ä->5	å->1	
de, o	c->22	m->3	
de, p	r->1	å->3	
de, s	a->1	k->3	o->8	ä->1	å->3	
de, t	a->1	i->1	o->1	r->1	y->1	ä->1	å->1	
de, u	t->3	
de, v	a->4	e->1	i->6	å->1	
de, ä	n->1	r->2	
de, ö	k->1	
de- o	c->1	
de-Fr	a->2	
de-Lo	i->1	
de-lä	n->1	
de. D	e->2	
de. M	e->1	
de. O	c->1	
de. V	i->2	
de.- 	F->1	
de.. 	(->1	
de.At	t->1	
de.Av	 ->1	s->2	
de.De	 ->1	n->4	s->2	t->32	
de.Dä	r->4	
de.Ef	t->2	
de.Em	e->1	
de.En	 ->4	d->1	
de.Eu	r->1	
de.FP	Ö->1	
de.Fr	u->2	
de.Fö	r->7	
de.Ge	n->1	
de.Gr	u->1	
de.Ha	n->2	
de.He	l->1	r->6	
de.Ho	n->1	
de.Hu	r->1	v->4	
de.I 	d->1	v->2	
de.Id	é->1	
de.In	f->1	o->1	
de.Ja	g->35	
de.Ka	n->2	
de.Ko	m->2	
de.Li	k->1	
de.Ly	c->1	
de.Lå	t->2	
de.Ma	n->4	
de.Me	d->1	n->9	
de.Mi	n->3	
de.Må	n->1	
de.Ni	 ->1	
de.Nu	 ->1	
de.Nä	r->2	
de.Oc	h->3	
de.Om	 ->3	
de.Pa	r->1	
de.Pl	a->1	
de.Po	r->1	
de.Pr	o->1	
de.Re	s->1	
de.Sa	v->1	
de.Sc	h->1	
de.Se	d->1	
de.Sl	u->2	
de.So	m->4	
de.St	ö->1	
de.Så	 ->2	
de.TV	-->1	
de.Ta	 ->1	c->3	
de.Ti	l->1	
de.To	p->1	
de.Tr	a->1	o->1	
de.Tv	ä->1	
de.Un	d->2	
de.Va	d->2	r->1	
de.Vi	 ->9	t->1	
de.Åt	e->1	
de: "	A->1	v->1	
de: A	n->1	r->2	
de: D	e->2	
de: F	l->1	r->1	ö->1	
de: G	e->2	r->1	
de: H	a->1	
de: I	 ->1	
de: J	a->1	o->1	
de: K	o->2	ä->1	
de: M	a->1	
de: N	y->1	ä->1	
de: P	o->1	
de: S	t->2	
de: T	u->1	
de: U	t->1	
de: V	a->2	i->1	
de: b	a->1	
de: f	ö->1	
de: h	u->1	
de: i	 ->1	
de: k	o->1	
de: t	o->1	
de: Å	t->2	
de; d	e->2	
de; h	ä->1	
de; m	i->1	
de; p	u->1	
de?De	n->1	
de?Fö	r->1	
de?He	m->1	r->2	
de?Ja	g->1	
de?Vi	l->1	
deHer	r->1	
dePro	t->1	
deadl	i->1	
deal,	 ->1	
deala	 ->1	
deale	n->1	t->1	
deali	s->1	
deaux	,->1	
debat	t->170	
debes	t->1	
debud	 ->6	,->2	e->1	
debän	k->1	
decem	b->19	
decen	n->7	t->15	
dedel	 ->1	a->1	
deell	a->2	
deers	ä->2	
defin	i->36	
defon	d->1	
defri	h->1	
deful	l->7	
deför	b->1	e->1	f->7	h->2	k->1	s->1	
degem	e->3	
degen	e->1	
degra	d->1	
dehöj	a->1	
deira	 ->1	.->1	
dekod	 ->5	e->3	
dekol	l->1	
dekri	s->1	
dekva	t->5	
del (	k->2	
del -	 ->1	
del K	o->1	
del a	n->2	t->3	v->79	
del b	e->1	ä->1	ö->1	
del d	e->1	
del f	a->1	o->1	r->4	ö->16	
del h	a->2	y->1	
del i	 ->12	n->1	
del k	a->1	o->2	v->1	
del l	i->1	
del m	a->1	e->6	å->1	
del n	ä->1	
del o	c->14	m->1	
del p	a->1	e->1	o->1	å->5	
del s	a->3	k->1	o->11	å->1	
del t	i->4	o->1	
del u	n->1	r->1	t->1	
del v	i->1	
del ä	n->1	r->7	
del ö	v->1	
del, 	a->1	d->2	e->1	f->2	i->1	k->2	l->1	m->3	n->1	o->6	s->1	v->2	
del.B	e->1	
del.D	e->5	
del.E	U->1	f->1	
del.J	a->2	
del.M	e->3	
del.N	ä->1	
del.S	å->1	
del.V	i->5	
del?J	a->1	
dela 	K->1	a->7	d->2	e->1	k->4	l->1	m->1	n->1	p->1	r->1	u->1	
delad	,->1	e->10	
delag	d->1	
delak	t->8	
delan	d->44	
delar	 ->52	,->3	.->7	:->1	e->1	n->9	
delas	 ->6	,->2	.->1	p->1	
delat	 ->7	,->1	.->1	s->8	
delay	e->2	
delba	r->19	
deleg	a->16	e->4	
delen	 ->25	,->7	.->2	F->2	
deles	 ->23	
delfr	å->1	
delgi	v->1	
delha	v->3	
delho	e->1	
dell 	m->1	s->2	
dell"	,->1	.->1	
dell.	D->1	
delle	n->3	r->3	
dellå	n->4	
dellö	s->1	
deln 	m->1	o->1	
delni	n->41	
delpu	n->2	
delra	p->1	
dels 	a->6	d->1	f->2	k->1	o->1	s->1	t->2	å->1	
dels-	 ->1	
delsd	r->1	
delse	 ->50	,->4	-->1	.->11	a->1	b->1	f->9	l->3	m->1	n->18	r->32	u->1	v->1	x->1	
delsf	l->2	r->2	
delsh	a->1	i->1	
delsi	n->2	
delsk	o->2	r->2	v->1	
delsl	a->5	o->1	
delsm	y->9	ä->2	
delsn	y->1	
delso	m->2	r->3	
delsp	l->2	o->2	r->2	
delss	e->1	j->1	t->1	ä->43	
delst	a->4	i->1	o->41	
delsv	a->1	
delta	 ->15	,->2	g->30	r->9	
delti	d->2	
delto	g->2	
delut	b->2	
delvi	s->11	
delös	a->1	
dem 2	0->1	
dem a	t->5	v->1	
dem d	e->4	ä->1	å->2	
dem e	f->1	n->3	t->2	
dem f	r->3	ö->5	
dem g	r->1	ö->1	
dem h	a->2	e->1	
dem i	 ->8	n->2	
dem j	a->1	
dem k	r->1	
dem l	ä->1	
dem m	e->3	y->1	ö->1	
dem n	å->1	
dem o	c->9	m->1	
dem p	å->7	
dem r	e->1	
dem s	e->1	o->59	å->1	
dem t	i->5	
dem u	t->4	
dem v	a->1	e->1	
dem ä	r->1	
dem, 	e->2	f->1	h->1	m->1	s->1	v->3	ä->1	å->1	
dem.(	A->1	
dem.A	v->1	
dem.B	e->1	u->1	
dem.D	e->4	ä->2	
dem.E	n->1	
dem.F	r->1	ö->1	
dem.H	e->1	
dem.J	a->4	
dem.K	o->1	
dem.M	e->3	
dem.N	e->1	å->1	
dem.O	m->1	
dem.R	e->1	
dem.V	i->6	
dem: 	d->2	
dem?D	e->1	
demag	o->4	
demar	k->1	
demas	k->1	
demen	i->5	
demi,	 ->1	
demin	s->1	
demis	k->1	
demog	r->3	
demok	r->136	
demon	s->6	t->8	
den "	d->1	e->1	n->1	
den (	E->1	
den ,	 ->1	
den -	 ->11	
den 1	 ->9	0->1	1->2	3->2	4->5	5->1	6->1	7->2	8->4	9->6	
den 2	 ->1	0->14	1->1	4->1	6->1	
den 3	 ->4	0->1	1->2	
den 4	 ->2	
den 5	 ->1	
den 6	 ->1	
den 7	 ->1	
den 9	 ->2	
den B	e->2	
den E	U->1	u->3	
den G	a->1	r->1	
den J	o->1	
den K	a->2	i->1	o->2	
den L	a->1	
den P	r->3	
den R	a->1	
den T	h->1	
den X	X->1	
den a	b->1	d->2	g->1	k->6	l->18	m->3	n->62	r->5	s->1	t->18	v->30	
den b	a->8	e->38	i->4	l->4	o->4	r->13	u->4	y->3	ä->5	ö->5	
den c	e->3	
den d	a->14	e->27	i->1	j->1	o->2	r->1	ä->11	å->2	ö->4	
den e	f->4	g->5	k->31	l->4	n->41	p->1	r->1	t->3	u->77	x->7	
den f	a->4	e->1	i->6	j->3	o->3	r->42	u->1	y->2	å->2	ö->127	
den g	a->7	e->53	i->1	j->3	l->7	o->6	r->13	y->1	ä->4	å->3	ö->2	
den h	a->36	e->3	i->2	j->2	o->3	u->1	y->1	ä->60	å->2	ö->8	
den i	 ->45	c->1	d->1	h->1	l->1	n->116	r->3	s->8	t->4	
den j	u->4	
den k	a->18	e->1	i->1	l->2	o->47	r->6	u->6	v->1	ä->2	
den l	a->4	e->3	i->5	o->3	ä->3	å->3	ö->3	
den m	a->4	e->32	i->12	o->11	u->3	y->7	ä->4	å->21	ö->2	
den n	a->5	e->1	i->1	o->5	u->15	y->36	ä->8	å->1	ö->5	
den o	a->2	b->13	c->73	f->9	k->1	l->1	m->11	p->1	r->16	s->1	t->1	u->1	v->1	
den p	a->7	e->8	l->6	o->24	r->17	u->18	å->26	
den r	a->4	e->27	i->8	o->2	y->1	ä->20	å->1	ö->1	
den s	a->6	e->18	i->14	j->14	k->37	l->10	n->4	o->104	p->9	r->1	t->45	u->1	v->4	y->6	ä->2	å->2	ö->1	
den t	a->2	e->6	i->47	j->1	o->9	r->6	u->3	y->16	
den u	n->6	p->11	r->3	t->19	
den v	a->8	e->10	i->27	o->2	ä->7	å->1	
den z	i->1	
den ä	g->1	n->10	r->39	v->2	
den å	 ->1	s->7	t->5	
den ö	k->4	n->3	p->2	s->15	v->7	
den" 	e->1	
den) 	f->1	
den)(	P->2	
den),	 ->1	
den).	D->1	
den, 	1->1	B->2	K->1	P->1	a->2	b->7	d->10	e->1	f->12	h->3	i->7	j->1	k->6	l->1	m->10	n->2	o->20	s->18	t->3	u->3	v->6	ä->4	
den. 	D->1	I->1	M->1	
den..	 ->2	(->1	
den.A	l->1	t->1	v->4	
den.D	e->37	ä->2	
den.E	U->1	n->3	r->1	t->2	
den.F	a->1	r->1	ö->10	
den.H	a->2	e->6	i->1	o->1	ä->1	
den.I	 ->9	
den.J	a->18	
den.K	o->6	u->1	
den.L	å->2	
den.M	a->2	e->7	i->1	
den.N	i->1	u->1	ä->1	
den.O	m->2	r->2	
den.P	å->4	
den.R	å->1	
den.S	e->1	i->1	l->3	o->1	y->1	å->1	
den.T	a->1	h->1	i->1	
den.U	n->2	
den.V	a->2	i->14	
den.Ä	v->1	
den: 	D->1	H->1	K->1	d->1	f->1	v->1	
den:F	ö->1	
den; 	d->4	
den?D	e->3	
den?N	ä->1	
den?V	a->1	e->1	
denNä	s->1	
dena 	-->1	B->1	a->4	e->2	f->9	i->9	k->3	l->1	m->2	o->10	p->2	r->1	s->3	t->1	u->1	v->1	ä->2	
dena,	 ->13	
dena.	 ->1	D->2	E->1	F->1	J->4	O->1	V->2	Ä->1	
dena;	 ->1	
dena?	P->1	
denas	 ->1	
denau	e->1	
denbu	r->2	
denie	d->2	
denna	 ->511	,->2	.->8	?->1	
denne	 ->2	s->3	
dens 	I->1	a->3	b->2	e->1	f->7	h->1	i->2	k->1	l->3	m->3	o->4	p->4	s->9	t->3	u->11	v->2	ä->1	
dens,	 ->2	
densa	m->4	
dense	n->2	r->5	
densi	s->2	
dent 	A->1	C->1	a->1	p->1	t->1	
dent,	 ->1	
dente	n->4	r->1	
denti	e->2	f->10	t->8	
dentl	i->25	
dents	k->1	
deolo	g->5	
depar	t->9	
der -	 ->4	
der 1	9->8	
der 2	0->2	
der 4	0->1	
der E	G->1	l->1	u->4	
der F	N->2	
der I	 ->1	I->1	
der L	a->7	
der N	i->2	
der U	N->1	S->1	
der a	l->13	n->2	t->15	u->1	v->9	
der b	a->1	e->10	i->2	l->1	o->2	r->3	u->2	ö->2	
der d	a->3	e->152	i->1	o->1	r->1	ä->5	å->2	
der e	c->1	d->1	f->6	k->1	l->4	m->3	n->18	r->2	t->7	u->8	x->2	
der f	a->2	e->1	i->1	l->2	o->2	r->10	u->2	y->1	å->2	ö->74	
der g	e->5	i->1	j->1	o->3	r->1	y->2	å->1	
der h	a->9	e->11	i->1	o->3	u->3	ä->2	
der i	 ->35	l->1	n->33	
der j	a->3	o->1	u->1	
der k	a->5	o->15	r->4	u->2	
der l	e->1	i->3	y->1	ä->1	å->2	ö->1	
der m	a->9	e->12	i->23	o->9	y->2	ä->1	å->12	ö->2	
der n	a->1	i->2	u->3	ä->7	å->6	
der o	c->44	f->2	m->4	s->14	u->1	
der p	a->1	e->2	l->3	o->1	r->6	u->2	å->19	
der r	a->1	e->11	i->1	o->1	u->1	ä->3	å->1	
der s	a->7	e->7	i->19	k->9	l->1	m->1	o->85	p->2	t->7	y->1	å->8	
der t	a->2	i->33	o->2	r->7	v->3	ä->1	
der u	n->5	p->4	r->1	t->11	
der v	a->10	i->21	ä->1	å->5	
der ä	m->2	n->2	r->7	
der å	r->9	t->2	
der ö	v->1	
der" 	h->1	
der) 	B->1	V->1	
der)F	r->2	
der)J	a->1	
der)K	o->1	
der)T	a->1	
der, 	a->2	b->1	d->4	e->1	f->5	h->4	i->2	j->1	k->1	l->1	m->7	o->15	p->2	s->12	t->1	u->1	v->5	ä->2	å->1	ö->1	
der-p	r->1	
der. 	D->2	S->1	V->1	
der..	V->1	
der.A	t->2	v->2	
der.B	a->1	l->1	
der.C	S->1	
der.D	a->1	e->22	ä->3	
der.E	n->2	x->1	
der.F	r->4	ö->1	
der.H	ä->1	
der.I	 ->6	n->1	
der.J	a->12	
der.K	o->3	
der.M	e->3	
der.N	a->1	ä->1	
der.O	m->1	
der.R	å->1	
der.S	o->1	t->1	
der.T	i->1	r->1	
der.U	n->4	
der.V	a->3	i->2	
der.Ä	r->2	v->1	
der: 	k->1	
der; 	v->1	
der?.	 ->1	
der?H	e->1	
der?Ä	v->1	
dera 	E->1	a->2	d->5	e->2	f->1	g->1	i->3	k->1	l->1	o->1	p->1	r->3	v->2	ö->6	
dera,	 ->1	
dera.	I->1	
derad	e->7	
deral	 ->2	i->6	t->2	
deran	d->1	
derar	 ->26	,->1	
deras	 ->91	,->2	
derat	 ->5	.->1	i->2	
derba	r->1	
derbl	å->2	
derbö	r->11	
derde	l->4	
derdo	m->2	
dereg	l->3	
dergr	ä->4	
dergä	l->1	
derhu	s->2	
derhå	l->3	
deri,	 ->1	
derie	r->2	
derin	g->59	
derka	s->2	t->2	
derku	r->1	
derla	g->7	
derle	v->2	
derli	g->10	
derlä	g->1	n->18	t->18	
derlå	t->3	
derma	n->2	t->1	
derme	n->1	
dermi	n->1	
dermå	l->1	
dern 	f->2	l->2	o->1	p->1	s->1	
dern,	 ->1	
derna	 ->170	!->1	,->29	.->36	/->1	?->4	r->1	s->18	
derne	a->1	
derni	s->24	
dernt	 ->1	
deror	d->4	
derre	p->2	
derrä	t->1	
ders 	a->2	b->2	e->1	f->1	i->1	l->2	n->1	o->2	p->6	r->2	s->3	t->1	v->1	å->1	
dersa	m->1	
dersk	a->3	o->1	r->2	
dersm	å->1	
dersp	e->2	
derst	r->30	ä->3	ö->6	
derså	t->1	
dersö	k->48	
derta	g->1	
derte	c->17	
derti	l->1	
derut	b->2	v->1	
dervi	s->1	
dervä	r->1	
derät	t->3	
derös	t->1	
des -	 ->2	
des 1	9->3	
des 2	 ->1	
des A	d->1	
des S	p->1	
des V	i->1	
des a	n->1	t->5	u->1	v->23	
des b	e->2	l->1	o->1	r->1	ä->1	
des d	e->9	ä->2	å->1	
des e	l->2	m->2	n->2	t->4	
des f	a->1	i->1	l->1	o->1	r->3	ö->12	
des g	e->1	ö->1	
des h	a->3	e->1	ä->1	å->1	ö->2	
des i	 ->25	g->1	n->7	
des j	u->1	
des k	l->2	o->3	r->1	u->1	
des l	e->1	
des m	a->2	e->3	ö->3	
des n	o->1	å->1	ö->2	
des o	c->9	m->3	
des p	o->1	r->1	å->3	
des r	e->2	
des s	a->1	e->1	k->1	o->4	t->2	
des t	i->9	v->1	y->3	
des u	n->3	p->4	r->1	t->1	
des v	i->4	o->1	ä->1	
des ä	n->1	r->1	
des, 	a->1	e->1	g->1	o->3	t->1	v->1	
des.)	Å->1	
des.D	e->1	ä->1	
des.I	 ->1	
des.J	a->1	
des.M	e->1	ä->1	
des.R	e->1	
des.U	n->1	
desam	m->2	
desbe	s->1	
desdi	g->2	
desge	m->1	
deska	p->113	
deski	f->1	
desky	l->1	
despe	r->7	
dess 	a->5	b->7	d->5	e->6	f->10	g->4	h->2	i->8	k->5	l->2	m->5	n->3	o->4	p->2	r->7	s->10	t->3	u->3	v->3	ä->2	å->3	ö->2	
dessa	 ->332	!->1	,->4	.->7	
dessk	a->1	
desst	r->1	
dessu	t->36	
dessv	ä->4	
desta	t->1	
desto	 ->2	
destr	u->1	
destå	n->1	
desvi	s->2	
det "	K->1	e->1	r->2	
det (	B->2	I->1	f->1	h->1	i->1	k->1	
det -	 ->8	
det 2	1->1	2->1	
det A	k->1	
det B	N->1	r->1	
det C	a->1	
det E	l->1	r->1	u->2	
det G	r->1	
det I	t->1	
det K	o->1	
det M	i->1	o->2	
det P	o->3	
det S	E->1	v->1	
det T	u->1	
det a	b->4	c->2	k->5	l->16	m->1	n->71	r->18	t->61	v->226	
det b	a->11	e->56	i->5	l->15	o->2	r->9	u->2	y->2	ä->5	ö->8	
det c	e->2	i->3	
det d	a->13	e->14	i->4	o->6	r->4	y->1	ä->10	å->9	ö->2	
det e	f->1	g->9	k->7	l->4	m->2	n->56	r->4	t->10	u->26	v->2	x->6	
det f	.->1	a->66	e->11	i->111	j->4	l->3	o->10	r->44	u->5	ä->1	å->13	ö->154	
det g	a->6	e->12	i->3	j->2	l->3	o->6	r->4	ä->185	å->11	ö->11	
det h	a->83	e->9	i->3	o->5	y->1	ä->56	å->1	ö->4	
det i	 ->74	b->2	d->1	g->1	l->1	n->127	r->2	t->3	
det j	a->7	o->1	u->7	ä->1	
det k	a->24	l->7	n->1	o->52	r->19	u->3	v->1	y->1	ä->2	ö->1	
det l	a->9	e->1	i->9	o->2	u->1	y->1	ä->12	å->3	ö->1	
det m	a->7	e->39	i->8	o->11	u->3	y->14	å->29	ö->28	
det n	a->6	e->1	i->4	o->2	u->28	y->19	ä->10	å->8	ö->12	
det o	a->5	b->1	c->81	e->1	f->7	l->1	m->30	n->2	r->2	s->1	t->1	
det p	a->4	e->6	l->2	o->61	r->11	å->15	
det r	a->2	e->15	i->4	y->1	ä->10	å->11	ö->9	
det s	a->24	e->12	i->6	j->5	k->83	l->8	o->119	p->8	t->48	u->3	v->5	y->6	ä->37	å->19	ö->1	
det t	a->5	i->46	j->1	o->3	r->24	v->2	y->10	ä->2	
det u	n->10	p->23	r->3	t->21	
det v	a->55	e->16	i->84	o->7	ä->11	å->2	
det y	t->6	
det ä	g->1	m->1	n->20	r->310	v->7	
det å	l->2	r->4	t->7	
det ö	g->1	k->3	n->2	p->2	s->14	v->7	
det!.	 ->1	(->1	
det) 	h->1	
det)N	ä->1	
det, 	I->1	a->5	b->1	d->5	e->4	f->9	g->4	h->6	i->3	j->2	k->4	l->2	m->12	n->2	o->15	p->5	r->2	s->21	t->3	u->3	v->8	ä->2	
det. 	(->1	D->3	S->1	V->1	
det.(	A->1	P->1	
det.-	 ->1	
det..	 ->2	
det.A	l->1	n->2	v->3	
det.B	l->1	
det.D	e->24	ä->2	
det.E	G->1	f->1	k->1	n->4	t->1	u->2	
det.F	l->1	ö->1	
det.H	e->9	u->1	ä->2	
det.I	 ->5	b->1	n->1	
det.J	a->20	
det.K	ä->1	
det.L	å->1	
det.M	a->3	e->8	i->2	
det.N	u->3	
det.O	c->2	
det.P	r->1	u->1	å->3	
det.S	k->1	l->1	å->3	
det.T	a->1	i->1	
det.U	r->1	t->1	
det.V	a->1	i->19	å->1	
det.Ä	n->1	
det.Å	 ->1	t->1	
det.Ö	s->1	
det: 	U->1	f->1	o->1	
det; 	d->1	
det?.	 ->1	(->1	
det?D	e->2	
det?H	u->1	
det?I	 ->1	
det?J	a->1	
det?N	i->1	
det?V	i->1	
detak	t->1	
detal	j->34	
dets 	a->2	b->15	d->11	e->1	f->19	g->15	h->3	k->1	l->1	m->7	n->2	o->18	p->4	r->6	s->9	v->1	
dets,	 ->1	
detsa	m->5	
detta	 ->717	!->1	,->36	.->73	:->1	?->1	
deuro	p->2	
deutr	o->1	
deval	d->6	
devis	 ->2	
dez, 	i->1	
dez-k	a->2	
dfilm	e->1	
dfina	n->2	
dfråg	a->9	o->1	
dfull	 ->1	
dfäll	e->4	
dfödd	.->1	
dför 	d->1	e->2	g->1	i->1	k->1	m->1	o->1	s->2	
dför,	 ->2	
dföra	 ->3	.->1	n->223	
dförd	e->1	r->1	
dföre	d->2	
dförs	l->1	
dfört	.->1	r->1	
dföru	t->2	
dga E	U->1	u->1	
dga d	a->2	e->2	
dga f	o->1	ö->4	
dga g	e->1	
dga k	o->2	
dga m	a->1	e->2	
dga o	c->1	m->2	
dga p	å->1	
dga s	o->2	
dga u	n->1	t->1	
dga ä	n->1	r->1	
dga ö	v->1	
dga, 	f->1	
dga?D	e->1	
dgad 	d->1	p->1	r->1	s->1	
dgade	 ->2	
dgan 	f->2	o->6	s->1	
dgan.	V->1	
dgar 	a->1	d->1	k->1	s->1	
dgar.	D->1	
dgas 	d->1	e->1	m->1	p->1	s->1	
dgas,	 ->2	
dgas.	D->1	E->1	N->1	R->1	V->2	
dgat 	E->2	f->1	
dge F	u->1	
dge a	t->3	
dger 	a->3	d->2	e->1	m->1	s->1	u->1	ö->1	
dges 	a->2	e->1	i->2	
dget 	f->3	i->1	k->1	o->1	s->2	ä->1	
dget,	 ->4	
dget.	 ->1	D->2	K->1	M->2	
dgeta	n->1	r->2	
dgetb	e->1	
dgete	n->15	r->1	
dgetf	r->2	ö->9	
dgetk	o->16	r->1	
dgetm	ä->1	
dgetp	l->3	o->11	
dgets	i->1	t->2	y->1	
dgett	 ->1	
dgetu	t->10	
dgetå	r->10	
dgetö	v->1	
dgiva	n->4	r->19	
dgivi	t->2	
dgivn	i->3	
dgnin	g->71	
dgor 	i->1	
dgrän	s->1	
dgrön	a->1	
dgäng	l->2	
dgång	 ->1	e->1	
dgård	 ->1	e->1	
dgått	 ->1	
dgör 	k->1	
dgörl	i->2	
dhet 	i->1	l->1	m->3	o->1	s->2	
dhet.	J->1	
dhete	n->3	
dhets	-->1	a->2	f->5	p->1	t->2	u->2	
dhist	i->1	
dhjäl	p->1	
dhåll	e->2	i->1	s->1	
dhöll	 ->1	
di - 	n->1	
di at	t->2	
di av	l->1	
di be	b->1	
di ha	r->2	
di in	g->1	
di lo	v->1	
di lä	m->1	
di oc	h->5	
di re	d->1	
di so	m->2	
di ta	l->2	
di, v	i->1	
di.De	t->1	
di.So	m->1	
di.Vi	l->1	
di: f	r->1	
di; m	a->1	
dia -	 ->1	
dia a	t->1	
dia h	a->1	
dia s	k->1	o->1	
dial 	b->1	
dialo	g->31	
diari	t->21	
dias 	o->1	
diatä	c->1	
dicap	 ->1	
dicer	a->1	
dicin	e->1	
didat	 ->1	e->1	l->12	
die R	e->1	
die a	v->1	
die o	c->1	
die, 	h->1	
diebe	s->1	
diekt	i->1	
dien 	h->1	o->3	
diens	 ->1	e->2	
diepr	o->1	
dier 	a->1	f->2	o->3	r->1	
dier,	 ->2	
dier.	D->1	K->1	M->1	
diern	a->2	
diet 	d->1	o->2	
diet.	V->1	
diffe	r->5	
difie	r->5	
dig a	t->1	
dig b	y->1	
dig d	a->1	e->2	i->1	
dig e	f->2	l->1	
dig f	u->1	ö->7	
dig g	e->1	
dig h	a->1	
dig i	 ->2	n->1	
dig j	u->1	
dig l	e->2	
dig m	e->2	o->1	
dig n	a->1	
dig o	c->6	
dig p	a->1	
dig r	e->3	ä->1	
dig s	l->1	t->1	
dig t	i->4	
dig, 	b->1	m->1	
dig.D	e->1	
dig.E	u->1	
dig.M	e->1	
dig.P	r->1	
dig.U	n->1	
diga 	-->1	E->1	H->1	a->5	b->3	d->5	e->1	f->5	g->4	i->3	k->4	m->4	n->1	o->4	r->5	s->5	t->1	u->2	v->1	ä->1	å->2	
diga,	 ->3	
diga.	D->1	H->1	I->1	M->1	
digan	d->4	
digar	 ->4	e->82	
digat	.->1	
digen	 ->1	
diges	 ->1	
dighe	t->250	
digna	 ->1	
digra	 ->2	
digst	ä->1	
digt 	-->3	a->40	b->4	d->7	e->7	f->20	g->2	h->6	i->4	k->7	l->5	m->17	o->17	p->3	r->6	s->33	t->5	u->4	v->10	ä->9	å->2	ö->1	
digt,	 ->10	
digt.	E->1	J->3	M->1	
digt?	A->1	
digtv	i->7	
dikal	 ->3	a->6	e->1	i->1	t->5	
dikap	p->4	
dikat	 ->2	,->1	i->1	o->5	
diken	,->1	
dikta	t->3	
dikte	r->2	
dikti	o->5	
dilem	m->3	
dimen	s->13	
dinav	i->1	
dinbu	r->1	
dinfl	y->1	
ding 	f->1	h->1	o->1	s->1	t->1	
ding,	 ->3	
dings	 ->1	
dingt	o->2	
dinsa	t->1	
dinsk	a->1	
dinst	r->1	
dinär	 ->1	
diolo	g->2	
dioxi	d->5	n->2	
diplo	m->11	
direk	t->248	
dirig	e->1	
dirlä	n->2	
dis B	a->1	
dis l	a->1	
dis p	o->1	r->1	
dis s	i->1	
dis u	p->1	
dis v	ä->2	
disci	p->14	
diser	i->9	
disk 	g->2	h->1	m->1	o->1	p->1	r->1	s->1	t->1	
diska	 ->32	
diskr	e->1	i->20	
diskt	 ->10	
disku	s->60	t->81	
dispe	n->1	
dispo	s->3	
dista	n->1	
disti	n->1	
distr	i->2	
dit F	P->1	
dit a	l->1	
dit d	ä->2	
dit f	i->1	ö->1	
dit h	ö->1	
dit l	e->1	
dit r	u->1	
dit s	i->3	
dit t	o->1	
dital	i->1	
diter	 ->1	,->1	
dithö	r->1	
ditio	 ->1	n->21	
dits 	o->1	
dium 	e->1	i->2	
dium.	Ä->1	
diver	s->4	
divid	 ->2	e->4	u->8	
diz e	l->1	
diz f	å->1	ö->1	
diz, 	G->1	
diz-k	a->1	
diär,	 ->1	
dja -	 ->1	
dja D	a->1	
dja H	a->1	
dja a	n->1	v->1	
dja d	e->28	
dja e	n->3	t->1	
dja f	o->1	ö->3	
dja i	n->1	
dja k	o->1	r->1	u->1	v->1	
dja l	o->1	
dja m	i->1	y->1	
dja o	c->1	l->1	s->3	
dja p	r->1	
dja r	e->1	
dja s	i->2	k->1	t->1	y->1	
dja t	i->2	
dja u	p->1	
dja v	å->1	
dja Ö	s->1	
dja å	t->3	
dja.H	e->1	
dja.J	a->1	
djan 	a->1	f->1	o->1	
djand	e->3	
djar 	d->1	o->2	p->1	t->1	å->1	
djas 	a->3	g->1	m->1	å->1	
djas,	 ->2	
dje -	 ->1	
dje a	s->1	t->1	
dje b	e->2	
dje d	e->2	
dje f	i->1	r->1	ö->1	
dje g	a->1	r->1	ä->1	
dje k	o->1	
dje l	a->22	ä->2	
dje m	i->2	å->2	
dje n	o->1	
dje o	c->2	
dje p	e->1	r->1	u->4	
dje r	i->2	
dje s	a->1	
dje v	i->2	ä->2	
dje ä	r->1	
dje å	r->1	
dje ö	v->3	
dje, 	a->3	v->1	
dje: 	u->1	
djede	l->6	
djekt	i->2	
djela	n->6	
djer 	m->1	
djorn	a->1	
djung	e->2	
djup 	ö->1	
djupa	 ->5	,->1	d->1	r->1	s->3	t->2	
djupe	t->5	
djupg	å->7	
djupn	i->5	
djups	i->1	
djupt	 ->7	
djur 	o->1	ä->1	
djur,	 ->2	
djur-	 ->2	
djur.	D->1	H->1	
djura	r->1	
djure	n->1	t->1	
djurf	o->4	
djurl	i->2	
djärv	 ->1	a->3	h->1	t->2	
djävu	l->2	
dkare	 ->1	
dkomm	a->15	e->5	i->4	
dkore	a->1	
dkurs	 ->1	
dkust	e->2	
dkvis	t->1	
dkänd	 ->1	,->1	a->5	e->18	
dkänn	a->32	e->13	s->1	
dkäns	l->5	
dkänt	 ->10	,->1	s->7	
dla d	e->7	
dla f	r->1	
dla g	e->1	
dla i	 ->1	g->1	
dla m	e->1	
dla o	m->7	
dla s	p->1	
dla u	n->1	
dla v	i->1	å->1	
dla.D	e->1	
dla.V	i->1	
dlad 	l->1	
dlade	 ->7	s->3	
dlag 	t->1	
dlagd	a->1	
dland	s->1	
dlar 	b->1	d->15	f->9	i->9	m->4	n->1	o->69	p->2	r->1	s->2	t->2	v->1	
dlare	 ->1	,->3	
dlarn	a->2	
dlas 	h->1	i->4	l->1	p->1	s->1	t->3	u->1	
dlas,	 ->1	
dlas.	B->1	
dlat 	a->1	e->1	f->1	k->1	s->2	
dlats	 ->1	
dlem 	a->1	i->2	o->1	u->1	
dlem,	 ->1	
dlemm	a->14	
dlems	k->2	l->36	r->1	s->284	
dlen 	a->1	b->1	f->3	i->1	k->1	m->1	s->2	
dlen,	 ->2	
dlet 	ä->1	
dlida	n->2	
dlig 	a->1	b->2	d->1	f->2	g->1	h->1	j->1	l->3	o->6	p->2	r->3	s->3	t->4	
dlig,	 ->1	
dlig:	 ->1	
dliga	 ->38	,->2	.->3	n->1	r->6	s->1	
dlige	n->16	
dligg	j->1	ö->3	
dligh	e->5	
dligt	 ->80	,->4	.->5	:->1	;->1	
dline	 ->1	
dling	 ->24	,->3	.->13	a->70	e->31	s->49	
dlinj	e->2	
dlist	a->1	
dlägg	a->74	n->5	
dlösa	 ->1	
dmakt	h->1	
dmede	l->3	
dmedl	e->1	
dmini	s->25	
dmium	 ->2	,->1	
dmont	e->3	
dmott	a->1	
dmän 	f->1	
dmåle	t->1	
dmåls	ä->1	
dmån 	d->1	
dna d	a->1	
dna e	t->1	
dna f	ö->1	
dna g	e->1	
dna k	o->1	
dna l	o->1	
dna m	e->1	
dna r	a->1	
dna s	t->2	
dna t	i->1	
dna u	p->1	
dna v	a->1	
dnack	a->2	
dnad 	f->1	i->2	j->1	o->1	r->1	
dnade	 ->4	
dnand	e->2	
dnapp	n->1	
dnar 	o->1	
dnare	 ->2	,->1	
dnarn	a->1	
dnas 	o->1	s->1	
dnat 	f->2	
dnats	.->1	
dning	 ->151	,->29	.->25	:->1	?->1	a->30	e->134	s->36	
dnivå	n->1	
do Ro	j->1	
do an	g->1	
do at	t->3	
do, a	t->1	
do.De	t->1	
do.Fö	r->1	
do.He	r->1	
do.Om	 ->1	
dock 	a->12	d->3	e->2	f->4	g->1	h->1	i->7	k->2	l->1	m->2	n->2	o->2	p->1	s->7	t->3	u->1	v->5	ä->1	å->2	
dock,	 ->2	
doeff	e->1	
dofil	s->1	
dog i	 ->1	
dog.D	e->1	
dog.S	a->1	
dogjo	r->1	
dogm 	e->1	
dogma	t->1	
dogör	 ->1	a->4	e->3	s->1	
dokum	e->45	
dolf 	H->2	
dolla	r->9	
dom a	v->4	
dom b	e->1	
dom d	e->1	
dom f	ö->1	
dom g	ä->1	
dom i	 ->1	
dom n	ä->1	
dom o	c->5	
dom p	å->1	
dom r	e->1	
dom ä	r->1	
dom, 	a->1	o->1	v->2	ä->1	
dom.D	e->1	
dom/r	i->1	
domar	 ->9	,->3	.->2	e->5	k->1	n->8	
domen	 ->9	,->1	
domin	a->1	e->7	
domli	g->3	
dområ	d->14	
doms 	s->1	
doms-	 ->2	,->1	
domsb	r->1	
domsf	r->3	u->1	
domsg	r->1	
domsh	e->1	
domsl	u->3	
domsr	ä->1	
domst	o->83	
don (	f->2	
don -	 ->1	
don b	ä->2	
don e	f->1	
don f	ö->1	
don i	 ->1	n->2	
don k	o->1	
don m	å->1	
don o	c->2	m->1	
don p	e->1	å->2	
don s	o->11	å->2	
don u	r->1	
don ä	r->1	
don, 	P->1	b->1	d->2	f->1	o->2	s->1	v->2	
don.D	e->3	
don.J	a->3	
don.L	å->1	
don.M	e->1	
don.O	m->1	
don.V	a->1	
don?V	i->1	
donNä	s->1	
donen	 ->5	.->1	
donet	.->1	
donsi	n->1	
donsp	a->1	
donst	i->3	
donsä	g->1	
donså	t->1	
dont 	a->1	
dor d	e->1	
dor f	ö->2	
dor h	a->1	
dor o	c->1	m->1	
dor p	å->2	
dor s	o->6	
dor u	p->1	
dor v	i->1	
dor, 	i->1	o->1	s->2	
dor.D	e->1	
dor.H	e->1	
dor.K	o->1	
dor.M	a->1	
dorde	t->1	
dorer	 ->1	n->1	
dorna	 ->8	,->3	
dorsa	k->1	
dosam	t->1	
dosed	d->1	
dosko	p->3	
dosta	s->1	
doste	u->1	
dou f	r->1	
dovis	a->3	n->1	
dox, 	s->1	
doxal	 ->2	a->1	t->2	
doämn	e->1	
dpela	r->1	
dpoli	t->1	
dprin	c->1	
dpunk	t->119	
dra -	 ->1	
dra E	E->1	U->1	u->1	
dra L	i->2	
dra R	i->1	
dra a	l->1	n->4	r->4	s->2	t->11	v->2	
dra b	a->2	e->10	i->2	ä->1	ö->2	
dra d	e->24	
dra e	f->2	l->2	n->6	t->3	u->1	
dra f	a->6	o->1	r->17	u->1	ö->8	
dra g	e->1	i->4	j->1	r->3	ä->2	å->2	ö->1	
dra h	a->3	e->1	o->1	u->1	ä->2	å->4	
dra i	 ->5	f->1	g->1	n->16	
dra k	a->1	o->10	u->1	ä->1	
dra l	a->2	e->1	o->1	ä->12	ö->1	
dra m	a->1	e->12	i->4	y->1	å->9	ö->3	
dra n	a->2	y->5	ä->1	å->2	
dra o	c->5	l->1	m->12	p->1	r->8	s->1	
dra p	a->1	l->1	o->3	r->3	u->9	å->8	
dra r	a->9	e->5	u->1	ä->1	å->2	
dra s	a->6	e->4	i->22	l->4	o->3	t->5	u->1	y->2	ä->2	å->3	
dra t	a->4	i->37	j->1	r->1	
dra u	n->1	p->2	t->1	
dra v	a->1	i->5	ä->7	
dra y	t->2	
dra ä	n->3	r->4	
dra å	r->2	t->1	
dra ö	v->1	
dra, 	a->4	d->2	g->1	i->3	k->1	m->2	o->1	p->1	s->3	u->2	v->2	ä->1	
dra.D	e->2	
dra.J	a->1	
dra.N	u->1	ä->1	
dra.U	n->1	
dra.V	i->1	
dra: 	I->1	g->1	u->1	Ä->1	
dra; 	f->2	
drabb	a->50	
drabe	h->5	
drad 	i->1	
drade	 ->13	,->2	.->3	s->3	t->3	
drag 	-->1	a->6	d->2	e->1	f->6	h->1	i->6	k->2	m->1	o->3	s->12	t->14	v->1	ä->3	å->2	
drag,	 ->2	
drag.	B->1	D->1	H->1	R->1	V->2	
drag:	 ->1	
draga	n->114	
drage	l->1	n->29	t->121	
dragi	t->12	
dragn	a->1	i->48	
drags	a->2	f->1	g->8	m->1	n->1	r->2	s->1	t->2	ä->3	
draha	n->1	
draka	m->1	
dram 	i->1	
drama	r->1	t->6	
dran 	o->3	s->1	t->2	ö->1	
dran,	 ->1	
dran.	N->1	
drand	e->5	
drar 	a->5	d->4	e->1	g->1	h->1	i->7	j->2	k->1	m->4	n->4	o->3	p->1	s->3	t->17	u->1	v->2	ä->2	å->1	
drar,	 ->1	
drare	 ->3	,->2	.->1	
drarn	a->3	
dras 	a->3	b->1	d->1	f->6	g->1	h->1	i->2	m->2	o->1	p->1	s->1	t->3	
dras,	 ->2	
dras.	D->1	E->1	S->2	V->1	
drast	i->3	
drat 	A->1	e->2	h->1	p->2	s->2	t->1	
drata	l->5	
drats	 ->5	,->1	.->4	
dratu	s->3	
dre a	k->1	v->1	
dre b	e->1	y->2	
dre d	e->1	
dre e	f->1	u->1	x->1	
dre f	a->3	o->1	r->1	ö->3	
dre g	e->1	
dre h	o->1	
dre i	 ->1	
dre k	o->2	r->1	ä->1	
dre l	e->1	ä->2	
dre m	e->1	
dre o	c->2	m->1	v->1	
dre p	e->1	u->1	å->2	
dre r	ä->1	
dre s	o->1	p->1	t->1	u->1	
dre t	i->1	y->1	
dre u	p->1	t->4	
dre v	i->1	
dre ä	n->9	r->1	
dre, 	h->1	v->1	
dre.D	e->2	
dre?V	i->1	
dreko	m->1	
dren 	f->3	
dresa	 ->2	
dret 	t->1	
drevs	 ->1	
driat	i->2	
drick	e->2	s->1	
drid 	i->1	
drid,	 ->1	
drid.	E->1	
drift	 ->2	.->1	e->1	i->1	s->3	
drig 	a->4	d->1	f->3	h->3	i->1	k->4	m->5	o->1	r->1	s->2	t->3	v->2	ä->1	å->1	
drikt	 ->1	,->1	i->1	
dring	 ->39	,->4	.->6	?->2	a->55	e->7	s->202	
driva	 ->22	n->1	s->2	
drive	n->5	r->8	t->5	
drivk	r->3	
drivn	a->1	
drivs	 ->5	,->1	.->1	
drog 	a->1	f->1	s->1	t->2	
drogb	e->1	
droge	r->1	
drogk	u->1	
drogs	 ->2	
droll	 ->1	,->1	
drome	t->1	
dron 	p->1	
dropp	e->1	
drott	 ->1	,->2	.->1	
druck	i->1	n->1	
drunk	n->3	
drust	n->1	
dryft	a->1	
drygt	 ->3	
dräge	r->36	
drägl	i->1	
dräng	 ->1	
dränk	t->2	
dråps	l->1	
dröja	 ->1	.->1	
dröjd	e->1	
dröje	r->3	
dröjs	m->2	
drömm	a->1	
ds al	d->1	
ds an	m->1	
ds at	t->1	
ds av	 ->6	
ds be	h->1	r->1	t->2	
ds bl	i->2	
ds bå	d->1	
ds de	m->1	n->1	
ds dä	r->1	
ds ef	t->1	
ds em	o->1	
ds en	d->1	
ds fe	l->1	
ds fö	r->4	
ds ge	n->1	
ds gr	ä->1	
ds i 	L->1	d->1	p->2	u->1	
ds in	o->2	t->2	
ds ju	 ->1	
ds la	g->1	
ds li	k->1	
ds me	d->5	
ds my	c->1	
ds ny	a->1	
ds ob	l->1	
ds oc	h->1	
ds om	 ->1	
ds pa	r->1	
ds på	 ->24	.->1	
ds re	g->2	t->1	
ds rå	d->1	
ds sa	m->1	
ds sk	a->2	u->2	
ds so	m->2	
ds ta	 ->1	
ds ti	l->1	
ds tr	e->1	
ds un	d->1	
ds ut	 ->1	
ds ve	r->1	
ds vi	d->1	
ds än	 ->1	
ds år	 ->1	
ds åt	 ->2	g->1	
ds ök	a->1	
ds öv	e->1	
ds, m	e->1	
ds, o	c->1	
ds, s	o->1	
ds, t	r->1	
ds- o	c->2	
ds-in	t->2	
ds-ny	t->1	
ds-si	t->1	
ds. D	e->1	
ds.Be	t->1	
ds.De	t->1	
ds.Ja	g->1	
ds.Un	d->1	
ds/in	t->1	
ds; b	)->1	
dsNäs	t->1	
dsak 	b->2	h->1	m->1	u->1	ä->1	
dsakl	i->10	
dsakt	ö->1	
dsam 	h->1	ö->1	
dsamm	a->1	
dsamt	 ->4	
dsand	e->3	
dsanm	ä->1	
dsans	t->1	
dsarb	e->5	
dsats	e->1	
dsavg	ö->3	
dsavt	a->3	
dsbed	ö->1	
dsbef	o->2	r->4	
dsbeh	a->1	
dsbes	k->1	l->1	t->1	
dsbev	a->1	
dsbus	s->1	
dsbyg	d->43	
dscen	t->1	
dsdel	 ->4	a->8	e->1	
dsdir	e->3	
dsdom	i->1	
dsdug	l->1	
dsdöm	d->1	
dseff	e->4	
dseko	n->15	
dsen 	m->1	
dsen,	 ->1	
dset 	f->1	
dsets	 ->1	
dsfal	l->1	
dsfri	 ->3	a->1	s->10	
dsfrå	n->1	
dsför	b->1	d->1	f->2	h->3	m->1	
dsgrä	n->1	
dshan	d->6	
dsinf	o->2	
dsinr	i->2	
dsins	t->2	
dsint	e->2	
dsitu	a->1	
dsjuk	a->1	
dsk a	n->1	
dsk k	a->3	
dsk t	e->1	
dsk-b	r->1	
dska 	a->1	b->1	e->1	f->3	i->1	k->1	l->1	m->2	o->4	p->1	r->1	s->1	t->1	
dska,	 ->2	
dskad	o->2	
dskal	v->1	
dskan	d->18	s->1	
dskap	 ->8	,->2	e->3	
dskar	.->1	
dskas	 ->8	
dskog	a->1	
dskom	m->1	
dskon	t->4	
dskra	f->1	
dskri	g->6	
dskrä	p->1	
dskt 	p->1	
dskär	n->3	
dsla 	h->1	m->1	o->2	
dsla,	 ->1	
dsla.	B->1	
dslag	 ->3	
dslan	 ->3	
dslib	e->1	
dslig	a->1	
dslis	t->1	
dslän	d->2	
dslån	g->1	
dslös	h->2	
dsman	n->10	
dsmar	k->1	
dsmed	b->6	e->3	l->2	
dsmin	i->1	
dsmyn	d->2	
dsmän	 ->3	
dsmäs	s->2	
dsmål	e->1	
dsmöj	l->1	
dsmöt	e->1	
dsniv	å->8	
dsomr	å->7	
dsoms	p->1	
dsord	f->20	
dsorg	a->2	
dsori	e->1	
dspak	e->2	
dspar	t->1	
dspat	i->2	
dspen	s->6	
dsper	i->4	
dspla	c->3	n->8	
dspol	i->3	
dspri	n->1	s->1	
dspro	b->3	c->22	d->1	g->5	j->1	
dspun	k->1	
dsram	,->1	a->4	
dsreg	e->1	i->2	
dsrep	u->4	
dsrym	d->2	
dsrät	t->1	
dsrör	e->1	
dssam	t->4	
dsski	l->1	
dsskä	l->1	
dssta	n->3	t->1	v->1	
dsstä	l->24	
dsstö	d->1	
dssys	s->1	t->1	
dssäl	l->1	
dstad	 ->1	,->1	
dstag	a->2	
dsten	a->1	
dstil	l->1	
dstjä	r->2	
dstop	p->1	
dstow	n->3	
dsträ	c->1	
dstul	l->1	
dstur	i->1	
dstäd	e->2	
dstäm	d->1	
dstän	g->2	
dsupp	g->1	s->1	
dsutt	r->1	
dsutv	e->1	ä->1	
dsver	k->1	
dsvil	l->2	
dsvin	s->1	
dsväg	,->1	
dsyft	e->1	
dsyst	e->4	
dsänd	a->1	
dsåld	e->2	
dsåtg	å->1	
dsöda	n->1	
dt fr	å->1	
dt ha	r->1	
dt oc	h->3	
dt sa	d->1	
dt ta	l->1	
dt ut	t->1	
dt, O	b->1	
dt, f	ö->2	
dt, i	 ->1	
dta a	t->1	
dta d	e->4	
dta e	n->5	r->1	
dta f	ö->10	
dta g	e->1	r->1	
dta j	o->1	
dta k	o->1	
dta l	ä->1	
dta m	e->3	
dta n	ä->1	å->1	
dta o	m->1	
dta p	o->1	å->1	
dta s	a->1	
dta u	p->1	
dta ä	n->3	
dta å	t->5	
dta.D	e->1	
dtabe	l->6	
dtagb	a->15	
dtagi	t->8	
dtagn	a->1	
dtala	t->1	
dtar 	g->1	i->2	k->1	n->1	o->3	s->1	v->1	y->1	
dtas 	d->1	f->2	i->1	m->1	n->3	o->1	s->2	t->1	v->1	ä->1	
dtas,	 ->2	
dtas.	D->1	J->1	P->2	Ä->1	
dter 	f->4	ä->1	
dter,	 ->1	
dterH	e->1	
dterb	e->2	
dters	 ->5	
dtes,	 ->1	
dtid.	V->1	
dtog 	i->1	r->1	
dtogs	 ->2	
dtyck	e->1	l->5	
dtysk	a->1	
du ba	i->1	
du be	r->1	
du co	m->1	
du mi	g->1	
du är	 ->2	
duali	t->1	
dubbe	l->6	
dubbl	a->11	
ducen	t->22	
ducer	a->12	i->1	
duell	a->6	t->1	
duer,	 ->1	
duga,	 ->1	
dugli	g->6	
dukar	 ->1	
dukt 	a->1	h->1	s->3	
dukt,	 ->1	
dukte	n->4	r->10	
dukti	g->1	n->1	o->21	v->9	
dukts	 ->2	
dumhe	t->3	
dumpa	n->1	
dumpn	i->3	
dumt 	a->1	
dunan	s->1	
dunkl	a->1	
duppb	y->1	
duppg	i->1	
duppr	ä->2	
durre	g->1	
dussi	n->1	
dustr	i->114	
dutsl	ä->1	
dutyp	,->1	
dvagn	e->1	
dval 	a->16	f->1	i->1	l->1	m->1	
dvala	r->3	
dvale	n->1	
dvatt	n->1	
dverk	a->19	
dveta	n->4	
dvete	n->14	t->7	
dvetn	a->17	
dvika	 ->27	s->4	
dvike	r->3	
dviki	t->1	
dvikl	i->4	
dvinn	i->2	
dvis 	a->1	u->1	ö->1	
dvoka	t->5	
dvrid	a->1	e->5	n->6	
dvrän	g->1	
dvs. 	1->2	E->1	W->1	a->11	d->4	e->3	f->3	g->1	h->2	i->5	j->1	m->4	n->1	o->2	p->1	s->1	v->2	
dvunn	a->1	
dvänd	i->125	n->1	
dvärd	e->1	
dväst	r->2	
dwill	 ->1	
dyka 	u->2	
dyker	 ->5	
dylik	a->2	t->1	
dynam	i->5	
dyr h	i->1	
dyra 	k->1	s->1	
dyrar	e->2	
dyrka	n->1	
dyrt 	o->1	
dyrt.	 ->1	
dystr	a->1	
dzio-	P->4	
dzjik	i->5	
däck 	o->1	
dämpa	 ->2	
där -	 ->1	
där 1	6->1	
där 2	9->1	
där 5	0->1	
där 8	0->1	
där E	U->2	u->2	
där F	P->1	
där L	u->1	
där a	l->3	n->2	r->3	v->1	
där b	e->4	r->2	å->1	
där d	e->43	
där e	l->1	n->5	r->1	t->1	
där f	i->3	l->1	r->1	ö->1	
där g	e->2	å->1	
där h	a->7	i->1	o->1	
där i	n->5	
där j	a->3	
där k	a->2	o->5	u->1	
där l	e->1	
där m	a->21	e->2	i->1	o->2	y->1	å->2	
där n	a->1	e->2	i->1	ä->1	
där o	c->3	
där p	r->2	å->2	
där r	e->1	i->1	
där s	a->2	e->1	i->1	j->1	k->2	o->2	p->1	t->5	å->1	
där t	i->1	j->2	v->1	
där u	n->1	t->4	
där v	a->1	e->2	i->24	
där Ö	s->1	
där ä	n->1	r->2	v->1	
där å	t->1	
där!D	e->1	
där, 	f->1	n->1	o->4	t->1	v->3	
där. 	D->1	
där.D	e->2	
där.F	ö->1	
där.I	 ->1	
där.J	a->3	
där.S	o->2	å->1	
där.V	a->1	i->2	
där?J	a->1	
därav	 ->2	
däref	t->7	
därem	o->13	
därfö	r->184	
därhä	n->1	
däri 	s->1	
därib	l->6	
därif	r->2	
därig	e->15	
därme	d->40	
därpå	 ->2	
därrä	t->1	
därti	l->1	
därva	 ->1	t->1	
därvb	r->1	
därvi	d->4	
därvl	i->1	
då 24	 ->1	
då As	s->1	
då Da	 ->1	
då EG	-->1	
då Er	i->1	
då Eu	r->1	
då ak	t->1	
då al	l->2	
då an	s->3	
då ar	b->1	t->1	
då at	t->11	
då ba	r->2	
då be	f->1	h->3	k->1	s->1	
då bl	i->3	
då bo	r->1	
då bö	r->4	
då de	 ->6	f->1	n->4	t->5	
då då	l->1	
då en	 ->6	
då fa	s->1	
då fi	n->2	
då fo	r->1	
då fr	a->2	å->2	
då få	r->2	
då fö	r->4	
då ge	n->3	
då gö	r->1	
då ha	d->2	n->1	r->3	
då he	l->1	
då i 	s->5	
då id	é->1	
då in	g->1	n->1	t->8	
då ja	g->2	
då ju	 ->1	
då ka	l->1	n->9	
då ko	m->4	
då kv	a->1	
då la	g->1	
då ma	n->2	
då me	d->1	n->2	
då my	c->1	
då må	s->2	
då mö	j->1	
då oc	h->1	k->6	
då oe	n->1	
då ol	j->1	
då om	 ->2	
då pe	s->1	
då po	l->1	
då pr	o->1	
då på	t->1	
då ri	s->1	
då rä	c->1	k->2	
då se	 ->1	
då sj	ä->1	
då sk	a->2	u->5	
då sn	a->1	
då so	c->1	m->2	
då sä	g->1	r->1	
då så	 ->1	
då ta	 ->1	l->3	
då ti	l->4	
då tr	a->1	
då tv	i->1	
då ty	c->1	
då tä	n->1	
då un	d->2	i->1	
då up	p->2	
då va	n->1	
då ve	r->2	t->1	
då vi	 ->5	d->1	k->1	l->1	s->1	
då vr	e->1	
då än	t->1	
då är	 ->2	
då äv	e->1	
då öv	e->1	
då, f	r->1	
då, m	e->1	
då, n	ä->1	
då...	.->1	
då.De	 ->1	
då?In	t->1	
dålig	 ->5	a->6	t->8	
dåtgä	r->6	
dåvar	a->1	
dé - 	f->1	
dé at	t->2	
dé ja	g->1	
dé ko	m->1	
dé om	 ->1	
dé so	m->3	
dé är	 ->1	
dé, m	e->1	
dée, 	v->1	
déer 	i->1	o->2	s->2	t->1	
déer,	 ->1	
déern	a->1	
dén a	t->6	
dén b	a->1	e->1	ö->1	
dén m	e->1	
dén o	m->3	
dén v	a->1	
dén, 	s->1	
dö i 	e->1	
död i	 ->1	
död o	c->2	
död v	a->1	i->1	
död.A	l->1	
död.J	a->1	
död.M	e->1	
döda 	o->1	
döda"	 ->1	
döda,	 ->1	
dödad	e->3	
dödan	d->1	
dödas	 ->1	,->1	
dödat	s->1	
dödfö	d->1	
dödsd	ö->1	
dödsf	a->1	
döend	e->1	
dölja	 ->5	.->1	
dölje	r->3	
döljs	 ->1	
döma 	H->2	a->3	d->4	e->2	f->2	h->2	i->1	o->3	p->1	r->1	s->2	t->1	v->2	
döma,	 ->1	
döma.	D->1	
döman	d->7	
dömas	 ->2	
dömba	r->1	
dömd,	 ->1	
dömde	.->1	s->1	
döme.	K->1	
dömer	 ->9	
dömes	g->1	
dömli	g->2	
dömni	n->28	
döms 	e->2	v->1	
dömt 	b->2	p->1	v->1	
dömts	 ->1	
döpa 	d->1	
döper	 ->2	
döpte	 ->1	
dör M	o->1	
dör e	l->1	
dör f	l->1	
dör m	ä->1	
dör u	t->1	
dörr 	ö->1	
dörr,	 ->1	
dörra	r->3	
dörre	n->4	
döstr	a->1	
dött.	D->1	J->1	
döttr	a->1	
dövt 	f->1	
e "al	d->1	
e "av	g->1	
e "de	n->1	
e "fö	r->1	
e "ko	l->2	
e "lä	s->2	
e "sv	a->1	
e (A5	-->29	
e (Be	n->1	
e (C5	-->2	
e (Ku	l->2	
e (ar	t->1	
e (fi	s->1	
e (ma	i->1	
e - ,	 ->1	
e - a	t->5	
e - d	e->4	
e - e	n->2	
e - f	å->1	ö->1	
e - h	a->2	
e - i	n->1	
e - j	a->3	
e - k	r->1	
e - m	i->1	
e - n	ä->1	å->2	
e - o	c->4	
e - p	å->2	
e - s	a->1	o->3	y->1	
e - t	e->1	
e - u	t->2	
e - v	i->1	
e - ä	v->2	
e -, 	i->1	
e 100	 ->1	
e 11 	s->1	
e 115	 ->1	
e 12 	m->1	
e 14 	m->4	
e 15 	o->1	p->1	r->1	
e 18 	m->1	
e 195	7->1	
e 199	2->1	6->1	8->1	9->1	
e 20 	å->1	
e 200	6->1	
e 21 	j->1	
e 25 	m->2	o->1	p->1	
e 26 	i->1	
e 35 	m->1	
e 4, 	o->1	
e 40 	p->1	
e 41 	p->1	
e 8 t	i->1	
e 9 m	i->1	
e Ahe	r->1	
e Alt	e->2	
e Ams	t->3	
e B t	a->1	
e BNP	,->1	
e Ban	k->1	
e Bar	n->1	
e Ber	n->1	
e Bes	q->1	
e Bus	q->1	
e Cen	t->2	
e Cur	i->1	
e Dan	m->1	
e De 	R->1	
e Dir	e->1	
e Dui	s->1	
e EMU	:->1	
e EU 	a->1	
e EU-	m->1	p->1	
e EU:	s->1	
e Eko	f->1	
e Eur	o->23	
e FN:	s->1	
e FoU	-->1	
e For	e->1	
e Fra	n->2	
e Fun	d->1	
e Gam	a->1	
e Gar	g->2	
e Gra	c->1	ç->1	
e Gro	s->1	
e Grö	n->1	
e Hai	d->1	
e Hed	g->1	
e Hit	l->1	
e Hol	z->1	
e Imb	e->1	
e Irl	a->1	
e Isr	a->1	
e Ita	l->1	
e Jac	q->1	
e Jon	c->1	
e Kar	a->1	l->1	
e Kin	n->3	
e Koc	h->2	
e Kou	c->1	
e Lan	g->1	
e Loy	o->1	
e Mar	i->3	t->1	
e Mel	l->1	
e Nap	o->1	
e Nat	o->1	
e OLA	F->1	
e Oil	 ->1	
e Ouv	r->1	
e Pal	a->7	
e Pla	n->1	
e Pro	d->13	v->2	
e Que	c->1	
e Rap	k->1	
e Rep	u->1	
e Rom	a->2	
e Roo	 ->1	
e Roy	a->1	
e San	t->1	
e Sch	e->1	r->1	
e Sei	x->1	
e Sve	r->1	
e Swo	b->1	
e Tri	t->1	
e Tur	k->1	
e Vat	a->1	
e Ven	s->1	
e Web	,->1	
e abs	o->2	
e acc	e->11	
e ad 	i->1	
e adj	e->1	
e adm	i->5	
e aff	ä->1	
e age	r->4	
e aid	s->1	
e akt	 ->2	i->1	u->5	ö->2	
e alb	a->2	
e all	 ->2	a->10	d->1	i->1	m->11	r->4	s->12	t->31	v->6	
e alt	e->1	
e amb	i->2	
e ame	r->3	
e an 	a->2	
e ana	l->7	
e anb	u->1	
e and	e->1	r->13	
e anf	ö->1	
e ang	e->3	r->2	å->2	
e ani	n->1	
e anl	e->5	ä->1	
e anm	ä->4	
e ann	a->1	
e ano	r->1	
e anp	a->3	
e ans	a->2	e->9	j->1	l->7	p->1	t->11	v->18	å->1	ö->1	
e ant	a->13	i->1	o->2	
e anv	ä->9	
e app	a->1	l->1	
e ara	b->3	
e arb	e->21	
e arg	u->2	
e art	i->3	
e asp	e->3	
e ast	r->1	
e asy	l->1	
e att	 ->241	
e aut	o->4	
e av 	E->4	F->1	L->1	S->2	a->19	b->4	d->31	e->18	f->16	g->5	h->4	i->5	j->1	k->11	l->2	m->6	n->1	o->8	p->5	r->6	s->16	t->24	u->6	v->5	y->1	å->1	
e av.	D->1	
e avd	e->1	
e avf	a->3	o->1	
e avg	e->1	i->1	ö->4	
e avr	e->1	
e avs	e->2	k->2	l->2	t->1	
e avt	a->6	
e avv	i->3	
e bak	o->2	
e bal	a->1	
e ban	d->3	
e bar	a->101	
e bas	 ->1	k->2	
e bea	k->2	r->1	
e bed	r->5	ö->4	
e bef	a->3	i->5	o->6	r->1	
e beg	a->1	r->7	ä->5	å->1	
e beh	a->7	o->5	å->2	ö->17	
e bei	v->1	
e bek	l->2	v->1	y->2	
e bel	g->2	o->1	
e ber	 ->1	e->1	o->1	ä->2	ö->8	
e bes	k->2	l->12	t->22	v->5	
e bet	a->7	e->1	j->1	o->2	r->11	y->11	ä->11	
e bev	a->3	e->1	i->5	
e bid	r->6	
e bif	a->1	
e bil	 ->1	a->11	d->2	i->1	k->1	p->1	t->1	
e bin	d->1	
e bio	 ->1	l->1	
e bis	t->2	
e bla	n->6	
e ble	v->1	
e bli	 ->25	r->13	v->2	
e blu	n->2	
e bok	s->1	
e bor	d->1	t->4	
e bov	a->1	
e bra	 ->2	
e bre	d->2	
e bri	n->1	s->6	t->1	
e bro	m->1	t->5	
e brä	n->1	
e bud	g->3	
e bur	i->1	
e byg	g->3	
e byr	å->7	
e byt	e->1	
e bär	a->2	
e bäs	t->5	
e bät	t->2	
e båd	a->4	e->3	
e båt	a->4	
e béb	é->1	
e bör	 ->7	d->1	j->10	
e cen	t->4	
e cha	p->1	
e che	f->3	
e civ	i->1	
e con	t->2	
e dag	 ->4	,->1	.->2	a->7	l->1	o->3	
e dam	e->3	
e dan	s->4	
e dat	u->1	
e de 	P->3	a->4	b->1	d->1	e->1	f->4	g->1	h->1	i->3	k->2	l->2	m->1	o->2	p->2	s->2	u->1	v->4	å->1	ö->1	
e deb	a->7	
e dec	e->4	
e def	i->1	
e deg	r->1	
e del	 ->3	a->6	e->9	s->1	t->6	v->2	
e dem	 ->8	,->1	.->1	o->6	
e den	 ->71	i->2	n->11	
e dep	a->1	
e der	a->1	
e des	s->12	
e det	 ->68	,->2	.->5	:->1	s->1	t->29	
e dia	l->1	
e die	 ->1	
e dip	l->1	
e dir	e->9	
e dis	c->3	k->9	p->1	
e dit	h->1	
e djä	r->1	
e doc	k->10	
e dog	 ->1	
e dom	a->1	s->3	
e dra	 ->1	b->12	
e dro	g->1	
e dry	g->1	
e drö	j->2	
e dus	s->1	
e dyk	e->2	
e där	 ->15	.->1	e->1	f->16	i->1	m->1	v->1	
e då 	a->1	d->3	f->1	g->1	m->2	o->1	t->1	v->1	
e då.	D->1	
e döl	j->1	
e döm	a->1	
e dör	r->1	
e eff	e->3	
e eft	e->12	
e ege	n->4	
e egn	a->2	
e ej 	ä->1	
e eko	n->27	
e el-	 ->1	
e ele	m->3	
e eli	m->1	
e ell	e->18	
e elm	a->1	
e eme	l->2	
e emo	t->3	
e en 	"->1	a->7	b->1	d->2	e->6	f->4	g->2	h->4	i->2	k->3	m->5	n->3	o->3	p->3	r->9	s->8	t->1	v->4	å->1	ö->1	
e enb	a->9	
e end	a->18	
e ene	r->4	
e eng	a->4	
e enh	e->2	ä->1	
e eni	g->1	
e enl	i->4	
e eno	r->4	
e ens	 ->7	a->1	k->14	
e ent	y->2	
e epo	k->2	
e er 	a->5	e->4	m->1	o->1	
e er.	B->1	
e era	 ->1	
e erb	j->2	
e erf	a->1	o->1	
e eri	n->1	
e erk	ä->4	
e ers	ä->1	
e eta	p->1	
e etn	i->2	
e ett	 ->49	
e eur	o->65	
e eve	n->3	
e ex 	p->1	
e exa	k->2	m->2	
e exe	m->3	
e exi	s->2	
e exp	e->16	
e ext	e->1	r->1	
e fac	k->2	
e fak	t->9	
e fal	l->19	
e fam	i->3	
e fan	n->5	t->2	
e far	h->1	l->1	o->2	t->9	
e fas	c->1	t->8	
e fat	t->7	
e fax	a->1	
e fel	a->1	
e fem	 ->7	,->1	t->4	
e fic	k->4	
e fil	o->1	
e fin	a->6	n->42	
e fis	k->4	
e fjo	r->3	
e fjä	r->1	
e fla	m->4	
e fle	r->5	s->24	
e fly	g->1	k->1	
e fol	k->5	
e fon	d->1	
e for	d->5	m->9	s->2	t->13	
e fra	m->38	n->6	
e fre	d->5	
e fri	-->6	a->1	h->3	s->1	t->1	
e fru	 ->4	k->1	
e frä	m->9	
e frå	g->49	n->49	
e ful	l->1	
e fun	g->10	n->2	
e fut	t->1	
e fyr	a->11	
e fäs	t->2	
e få 	E->1	a->2	b->1	e->8	f->2	l->1	m->1	n->1	o->3	p->1	r->1	s->1	t->2	v->3	
e får	 ->24	,->1	
e fåt	t->5	
e föl	j->5	
e för	 ->189	.->3	?->1	a->5	b->17	d->10	e->45	f->10	g->1	h->7	k->3	l->5	m->3	n->7	o->4	p->2	r->2	s->63	t->2	u->4	v->8	ä->9	ö->1	
e gam	l->6	
e gan	s->1	
e gar	a->10	
e gav	 ->3	
e ge 	a->1	d->3	e->2	i->1	o->1	r->2	s->1	v->1	
e gem	e->11	
e gen	a->1	d->1	e->4	o->27	t->3	
e geo	g->2	
e ger	 ->6	
e get	t->2	
e gil	t->1	
e giv	e->2	
e gjo	r->8	
e glö	m->11	
e god	a->4	k->3	s->3	t->11	
e got	t->1	
e gra	d->3	n->7	
e gru	n->22	p->5	
e grä	n->8	
e grå	 ->1	
e grö	d->1	n->7	v->1	
e gäl	l->11	
e gär	n->5	
e gå 	a->1	b->2	i->2	l->4	p->1	t->1	
e gån	g->11	
e går	 ->8	
e gåt	t->2	
e göm	m->1	
e gör	 ->7	a->34	
e ha 	a->1	b->2	d->3	e->6	f->1	g->3	h->1	k->3	m->1	n->3	s->4	t->2	v->5	ä->1	ö->1	
e had	e->13	
e haf	t->4	
e hal	t->1	v->3	
e ham	n->1	
e han	 ->7	d->20	s->2	t->2	
e har	 ->155	,->1	m->1	
e hel	a->2	l->42	t->11	
e hem	 ->1	f->1	l->2	m->1	s->1	
e hen	n->1	
e her	r->4	
e het	e->1	
e hie	r->1	
e hin	d->6	
e his	t->2	
e hit	t->4	
e hjä	l->5	r->1	
e hon	 ->3	o->2	
e hop	p->2	
e hor	d->1	
e hos	 ->4	
e hot	a->1	e->2	
e hur	 ->7	u->3	
e huv	u->1	
e hyc	k->1	
e hys	a->1	
e hän	d->4	g->1	s->1	t->1	v->1	
e här	 ->20	,->1	
e häv	d->1	
e hål	l->10	
e hår	d->1	t->1	
e hög	a->1	e->4	r->1	s->2	
e höj	n->1	
e höl	l->1	
e hör	 ->4	a->1	t->2	
e i A	f->1	
e i B	e->1	i->1	
e i D	a->2	
e i E	G->1	u->7	
e i F	i->1	r->1	
e i H	e->2	
e i I	r->1	t->1	
e i K	f->1	o->2	ö->1	
e i L	i->1	
e i S	h->1	t->1	
e i T	e->1	
e i a	k->1	l->6	r->1	t->2	v->1	
e i b	e->2	u->1	ö->1	
e i d	a->11	e->29	
e i e	f->1	g->2	n->3	t->4	u->1	
e i f	e->1	o->2	r->9	y->1	ö->8	
e i g	e->1	å->6	
e i h	a->2	e->2	u->2	
e i k	o->3	r->6	u->2	
e i l	a->2	
e i m	a->1	e->3	i->3	o->1	å->1	
e i n	a->1	o->2	ä->2	å->2	ö->1	
e i o	c->1	m->2	
e i p	l->1	o->1	r->3	
e i r	e->2	ä->1	å->1	
e i s	a->2	e->2	i->11	j->1	k->2	t->11	y->1	å->1	
e i t	i->7	r->2	
e i u	n->4	t->7	
e i v	a->1	e->1	i->1	å->3	
e i y	r->1	t->1	
e i z	o->1	
e i Ö	s->2	
e i ä	m->1	
e i å	r->5	
e iak	t->2	
e ick	e->8	
e ide	n->1	
e idé	 ->1	e->2	
e ifr	å->4	
e ige	n->1	
e ign	o->1	
e ill	a->1	
e imp	l->1	
e inb	e->2	j->1	l->4	
e ind	i->6	u->2	
e inf	l->2	o->7	r->1	ö->13	
e ing	a->2	e->9	r->1	å->3	
e ini	t->3	
e ink	r->1	
e inl	e->5	ä->3	ö->1	
e inn	a->3	e->20	
e ino	m->13	
e inr	e->3	i->3	ä->5	
e ins	a->4	e->4	i->1	k->2	l->1	t->17	
e int	a->1	e->81	r->9	y->1	
e inv	a->1	e->5	ä->2	
e iso	l->1	
e isr	a->3	
e ita	l->6	
e jag	 ->71	,->2	
e jet	t->1	
e jor	d->5	
e jou	r->2	
e ju 	a->1	m->1	o->1	
e jud	i->1	
e jur	i->1	
e jus	t->4	
e jäm	f->1	l->3	
e kam	p->3	
e kan	 ->110	d->1	s->4	
e kap	i->2	
e kar	g->1	
e kat	a->9	e->2	
e kem	i->1	
e kin	e->5	
e kla	r->7	s->2	
e kli	m->1	
e kna	p->2	
e knä	c->1	
e kol	d->1	l->18	
e kom	 ->2	m->143	p->7	
e kon	c->4	f->4	g->1	k->11	s->11	t->18	
e kor	r->1	t->2	
e kos	t->8	
e kra	f->1	v->10	
e kre	t->1	
e kri	n->2	s->3	t->5	
e kro	s->1	
e kry	p->1	
e krä	n->3	v->9	
e kul	t->5	
e kun	d->6	g->15	n->84	s->4	
e kus	t->2	
e kva	n->2	r->6	
e kvi	n->2	
e kvä	l->1	
e käl	l->1	
e kän	d->1	n->6	s->1	t->1	
e kär	l->1	
e kör	a->1	
e la 	L->1	
e lad	e->1	
e lag	a->2	r->1	s->11	t->1	
e lan	d->35	
e las	t->2	
e led	a->17	e->5	
e leg	a->2	
e let	t->1	
e lev	d->1	e->2	n->1	
e lib	a->1	e->4	
e lid	e->2	
e lig	g->7	
e lik	s->1	
e lin	j->1	
e liv	s->4	
e log	i->3	
e lok	a->8	
e lur	a->1	
e lyc	k->8	
e lys	s->2	
e läc	k->1	
e läg	e->1	g->5	r->2	
e läm	n->3	p->3	
e län	d->12	g->30	
e lär	a->1	t->1	
e lät	 ->3	t->2	
e lån	g->5	
e lås	t->1	
e låt	a->4	e->1	s->2	
e löf	t->1	
e lön	e->1	
e löp	e->1	
e lös	 ->1	a->4	n->1	t->1	
e maj	o->6	
e mak	r->1	t->8	
e man	 ->35	,->2	d->1	
e mar	k->74	s->1	
e mat	e->1	
e max	b->1	
e med	 ->111	b->6	d->1	e->11	f->3	g->3	i->1	k->1	l->19	v->2	
e mek	a->3	
e mel	l->14	
e men	 ->2	,->1	i->2	
e mer	 ->10	
e mes	t->22	
e met	o->3	
e mig	 ->6	r->1	
e mil	j->14	l->2	
e min	 ->2	a->1	d->7	i->3	s->20	u->1	
e mis	s->9	
e mit	t->1	
e mob	i->1	
e mod	e->2	
e mon	e->1	
e mot	 ->7	i->2	s->7	
e mul	t->4	
e myc	k->22	
e myl	l->1	
e myn	d->7	
e mäk	t->2	
e män	 ->1	g->1	n->10	s->21	
e mär	k->3	
e mål	 ->6	,->1	.->3	e->5	s->3	
e mån	a->23	g->16	
e mås	t->32	
e möj	l->12	
e mör	d->1	
e möt	e->1	
e nat	i->51	t->1	u->4	
e ned	e->1	v->1	
e neg	a->2	
e nek	a->1	
e ni 	a->1	d->1	e->1	g->1	h->1	i->1	s->1	
e nio	 ->7	
e niv	å->4	
e nog	 ->2	a->1	
e nor	d->5	m->6	r->1	
e not	e->4	
e nu 	-->1	b->1	f->3	i->1	k->1	l->1	o->1	p->1	s->1	ä->2	
e nuv	a->8	
e nya	 ->23	
e nyh	e->3	
e nyl	i->1	
e nys	s->4	
e nyt	t->1	
e näm	l->1	n->6	
e när	 ->21	a->2	m->11	v->1	
e näs	t->3	
e nät	.->1	
e nå 	e->1	
e någ	o->33	r->7	
e når	 ->1	
e nöd	v->7	
e nöj	a->5	d->2	t->1	
e oav	s->1	
e obe	g->1	h->1	r->2	
e och	 ->223	/->1	
e ock	s->57	u->1	
e oer	h->1	
e ofa	n->1	
e off	e->12	r->1	
e ofr	å->1	
e oft	a->1	
e ola	g->1	
e oli	k->45	
e olj	a->2	e->1	
e olo	g->1	
e oly	c->7	
e olä	m->1	
e om 	"->1	-->1	I->1	K->1	a->11	b->6	d->29	e->13	f->5	g->2	h->3	i->1	j->1	k->2	l->1	m->8	n->3	o->2	r->2	s->5	t->3	u->4	v->8	Ö->1	ö->2	
e om,	 ->3	
e om.	M->1	
e omb	u->2	
e ome	d->2	
e omf	a->7	
e omk	r->1	
e omp	r->1	
e omr	å->32	ö->4	
e oms	t->3	
e omö	j->1	
e ons	d->2	
e ope	r->1	
e opi	n->1	
e opp	o->1	
e opr	o->1	
e ord	 ->2	a->1	f->22	n->1	
e org	a->6	
e ori	m->1	
e ork	a->1	
e oro	 ->1	a->1	l->3	s->1	
e ors	a->3	
e orä	t->1	
e oss	 ->14	
e oti	l->1	
e ova	n->2	
e ove	r->1	
e ovi	s->1	
e ovä	d->1	
e pal	e->3	
e par	a->2	c->1	k->1	l->24	t->10	
e pas	s->1	
e pek	a->4	
e pel	a->2	
e pen	g->4	n->1	
e per	i->21	m->1	s->17	
e pes	s->1	
e pil	o->1	
e pla	c->1	n->7	t->1	
e pli	m->1	
e pol	i->35	
e pop	u->1	
e por	t->2	
e pos	i->5	
e pot	e->1	
e pra	k->3	
e pre	c->6	l->1	m->2	s->4	
e pri	m->1	n->19	o->3	s->1	v->2	
e pro	b->15	c->2	d->3	f->1	g->14	j->4	p->3	t->5	v->1	
e pub	l->2	
e pun	k->14	
e på 	8->1	E->3	F->1	T->1	a->29	b->3	d->35	e->16	f->6	g->11	h->3	i->2	j->1	k->4	l->6	m->10	n->14	o->3	p->1	r->6	s->7	t->3	u->4	v->4	ä->1	ö->1	
e på,	 ->2	
e påb	ö->2	
e påg	å->4	
e påm	i->1	
e påp	e->5	
e pås	k->2	t->1	
e qua	 ->2	
e rad	i->1	
e ram	a->2	p->6	
e rap	p->10	
e ras	i->3	
e rat	i->1	
e rea	g->5	k->3	l->1	
e red	a->8	e->1	o->1	
e ref	e->1	l->1	o->15	
e reg	e->25	i->40	l->16	
e rek	o->1	r->1	
e rel	a->1	e->1	
e ren	g->1	t->3	
e rep	r->1	
e res	a->2	e->1	o->3	p->8	t->2	u->15	
e rev	i->3	
e rik	a->5	e->4	t->15	
e ris	k->5	
e rol	l->9	
e ros	 ->1	
e rot	a->1	
e rub	b->2	
e rul	l->1	
e run	d->1	
e rut	i->1	
e ryk	t->1	
e räc	k->8	
e räd	d->1	
e räk	n->4	
e rät	t->50	
e råd	 ->2	,->1	a->4	e->8	f->1	g->2	s->5	
e rör	 ->2	l->1	
e rös	t->3	
e sad	e->2	
e sag	t->5	
e sak	 ->1	e->4	n->1	
e sam	a->6	b->1	h->1	m->10	o->2	r->1	s->1	t->9	
e san	k->3	n->2	t->1	
e sat	s->1	
e se 	a->2	m->1	o->1	p->2	t->9	ö->1	
e sed	a->14	
e sek	l->2	t->2	
e sen	 ->1	a->39	
e ser	 ->2	v->2	
e ses	 ->4	
e set	t->3	
e sex	 ->3	
e sif	f->2	
e sig	 ->30	n->1	
e sik	t->1	
e sin	 ->1	a->1	
e sis	t->4	
e sit	t->1	u->10	
e sju	 ->1	k->1	
e sjä	l->11	
e ska	d->13	l->48	p->7	r->1	t->2	
e ske	 ->5	,->1	d->1	r->2	t->1	
e ski	l->4	
e skj	u->5	
e sko	g->2	
e skr	i->1	o->1	
e sku	l->28	r->1	
e sky	d->5	l->2	
e skä	m->2	n->1	r->3	
e skå	d->2	
e skö	t->1	
e sla	g->1	
e sli	r->1	
e slu	t->8	
e slä	p->1	
e små	 ->22	
e sna	b->7	r->5	
e soc	i->13	
e som	 ->213	
e sop	a->1	
e sor	g->1	t->1	
e spa	n->1	
e spe	c->4	l->1	
e spr	i->1	å->1	
e spä	n->1	
e spå	r->2	
e sta	b->1	d->1	n->2	r->8	t->23	
e ste	g->3	
e sti	g->1	
e sto	d->1	p->1	r->27	
e str	a->6	i->2	u->7	y->2	ä->3	å->2	
e sty	r->4	
e stä	d->1	l->9	m->1	
e stå	 ->7	e->1	n->3	r->3	t->1	
e stö	d->20	r->8	
e sum	m->2	
e sun	d->1	
e suv	e->2	
e sva	g->3	r->6	
e sve	k->1	
e svå	r->7	
e syf	t->6	
e sym	p->1	
e syn	a->3	d->1	p->2	
e syr	i->1	
e sys	s->7	t->16	
e säg	a->13	e->5	
e säk	e->12	r->3	
e säl	l->1	
e säm	s->4	
e sän	d->2	
e sär	s->3	
e sät	t->29	
e så 	a->3	b->1	e->1	f->1	g->1	h->2	i->1	k->1	l->1	m->4	o->2	t->1	v->2	
e såd	a->1	
e sål	e->8	u->1	
e sår	b->1	
e sök	a->1	
e sön	d->1	
e sör	j->3	
e t.e	x->1	
e t.o	.->1	
e ta 	a->1	d->2	e->2	h->4	i->3	l->2	m->1	o->1	r->2	s->6	t->3	u->6	v->1	
e tac	k->2	
e tag	i->8	
e tak	t->1	
e tal	 ->2	a->21	e->2	m->3	r->1	
e tan	k->5	
e tar	 ->5	
e tas	 ->3	
e tax	-->2	
e tec	k->1	
e tek	n->6	
e ten	d->1	
e ter	r->1	
e tex	t->3	
e tid	 ->1	,->3	.->1	e->10	i->12	p->2	s->3	t->1	
e til	l->216	
e tio	 ->5	
e tis	d->1	
e tit	t->4	
e tja	t->1	
e tjä	n->12	
e tog	 ->2	
e tol	e->4	
e top	p->1	
e tot	a->3	
e tra	d->1	f->1	g->2	n->3	s->1	
e tre	 ->11	d->1	n->1	
e tro	 ->2	l->1	r->1	t->4	v->1	
e trä	f->1	t->1	
e tum	m->3	
e tun	g->1	
e tur	k->3	
e tus	e->1	
e tve	k->2	
e tvi	n->2	s->2	
e tvä	r->4	
e två	 ->21	.->1	
e tyc	k->3	
e tyd	l->4	
e tyn	g->1	
e tys	k->3	
e tyv	ä->1	
e täc	k->6	
e tän	k->3	
e ult	r->1	
e und	a->4	e->30	
e uni	k->1	o->3	
e upp	 ->4	,->3	b->2	e->1	f->19	g->15	h->1	l->1	m->7	n->8	r->8	s->11	
e ura	n->4	
e urb	a->1	
e urh	o->2	
e urs	ä->1	
e urv	a->1	
e ut 	1->1	d->3	e->1	i->1	k->1	p->1	r->1	
e ut,	 ->2	
e ut?	E->1	
e uta	n->15	r->2	
e utb	e->1	i->5	
e ute	l->1	s->2	
e utf	o->1	ä->2	ö->2	
e utg	i->1	j->1	å->6	ö->8	
e utk	a->1	r->1	
e utl	a->1	ä->1	å->1	
e utm	a->2	ä->1	
e utn	y->3	
e uto	m->1	
e utr	i->3	u->1	y->3	
e uts	a->1	e->1	i->1	k->1	l->1	t->5	
e utt	a->11	j->3	r->5	
e utv	e->12	i->15	ä->6	
e utö	k->2	v->3	
e vac	k->1	
e vad	 ->15	
e val	d->3	e->1	f->2	t->1	
e van	h->1	l->2	
e var	 ->17	a->99	f->1	i->7	j->3	k->1	s->1	t->1	v->1	
e vat	t->11	
e vec	k->11	
e vel	a->3	
e vem	 ->1	
e ver	k->19	s->2	t->2	
e vet	 ->1	a->1	e->13	
e vi 	-->2	5->1	a->6	b->2	d->1	e->2	f->6	g->7	h->8	i->11	j->1	k->5	l->3	m->1	n->4	o->6	p->1	r->1	s->15	t->6	u->4	v->6	
e vi,	 ->1	
e via	 ->1	
e vid	 ->6	a->1	h->1	t->7	
e vik	t->27	
e vil	j->72	k->12	l->20	
e vin	n->1	s->1	
e vir	k->1	r->1	
e vis	,->1	a->8	s->2	
e vit	b->1	
e vol	y->2	
e von	 ->2	
e vor	e->4	
e vra	k->1	
e väc	k->1	
e väg	a->1	e->1	l->1	
e väl	 ->2	d->1	f->1	j->1	
e vän	s->3	t->6	
e vär	d->8	l->4	n->2	s->1	
e väs	e->3	
e väx	e->1	
e vån	i->1	
e vår	 ->6	t->1	
e yrk	e->3	
e ytt	e->9	r->2	
e Öst	e->1	
e ägn	a->2	
e ägt	 ->2	
e äld	r->1	
e ämn	e->1	
e än 	1->2	2->2	3->1	E->1	W->1	a->4	d->6	e->1	f->4	i->4	j->1	k->2	l->1	m->1	n->4	r->1	s->3	t->2	v->7	ä->1	
e än.	J->1	
e änd	r->24	å->3	
e änn	u->5	
e änt	l->4	
e är 	E->1	a->13	b->9	d->13	e->20	f->13	g->1	h->6	i->14	j->4	k->8	l->3	m->11	n->4	o->2	p->3	r->5	s->8	t->10	u->3	v->4	y->2	ö->3	
e är.	J->1	
e äre	n->2	
e äve	n->9	
e å r	e->1	
e åkl	a->1	
e ålä	g->1	
e år 	1->3	2->1	a->1	i->1	k->1	p->1	s->5	å->1	
e år.	D->3	H->1	I->1	R->1	V->1	
e åre	n->26	t->2	
e årh	u->1	
e års	r->1	
e årt	u->1	
e åsi	k->3	
e åst	a->2	
e åt 	F->1	d->1	l->1	r->1	s->1	
e åta	g->5	l->2	r->1	
e åte	r->16	
e åtf	ö->3	
e åtg	ä->42	
e åtm	i->1	
e ått	a->1	
e öar	n->1	
e öka	 ->1	r->2	s->1	t->1	
e ökn	i->2	
e ömm	a->1	
e öns	k->11	
e öpp	e->8	n->3	
e öst	e->3	
e öve	r->52	
e övn	i->1	
e övr	i->12	
e! Ja	g->5	
e! Ni	 ->2	
e!All	t->1	
e!Det	 ->1	
e!Jag	 ->1	
e!Men	 ->1	
e!Ni 	h->1	
e!Ska	l->1	
e!Äve	n->1	
e" sk	a->1	
e" so	m->1	
e", i	 ->1	
e", o	c->2	
e(A5-	0->1	
e) fö	r->1	
e) i 	e->1	
e) oc	h->1	
e, , 	a->1	
e, Al	s->1	
e, Be	l->1	
e, Da	r->1	v->1	
e, Di	m->1	
e, Er	i->1	k->1	
e, Fr	a->1	
e, Fö	r->1	
e, Gr	a->1	
e, Ha	g->1	
e, Le	i->1	
e, Li	s->1	
e, Ra	f->1	
e, Sp	a->1	
e, al	l->1	
e, an	s->1	
e, ar	b->1	
e, at	t->15	
e, av	 ->1	f->1	
e, be	r->1	s->1	
e, bl	.->1	
e, bo	r->3	
e, br	o->1	
e, by	g->1	
e, bä	r->1	
e, bå	d->3	
e, bö	r->1	
e, de	 ->3	n->5	r->2	t->9	
e, dv	s->2	
e, dä	r->2	
e, då	 ->1	
e, ef	t->7	
e, em	e->1	
e, en	 ->3	
e, et	t->1	
e, ex	e->1	
e, fi	n->1	
e, fr	a->3	ä->1	
e, fö	r->10	
e, ga	v->1	
e, ge	n->1	
e, gö	r->1	
e, ha	n->2	r->5	
e, he	l->1	r->9	
e, hu	r->3	
e, hö	g->1	
e, i 	B->1	a->1	d->1	m->1	r->1	s->4	v->2	
e, in	f->2	k->2	o->2	t->5	v->2	
e, ja	g->4	
e, ka	n->5	
e, ki	d->1	
e, ko	f->1	m->4	r->1	
e, kr	i->1	
e, kä	r->1	
e, li	k->3	
e, me	d->4	l->1	n->16	r->4	
e, mi	n->1	
e, mo	t->1	
e, mu	s->1	
e, my	c->1	
e, må	s->1	
e, na	t->2	
e, ny	l->1	
e, nä	m->5	r->5	
e, nå	g->1	
e, nö	d->1	
e, oa	v->1	
e, oc	h->38	k->1	
e, om	 ->5	f->1	
e, os	t->1	v->1	
e, pr	e->2	o->3	
e, på	 ->5	
e, rö	r->1	
e, sa	l->1	m->1	
e, sk	a->2	e->1	u->1	y->1	
e, so	m->19	
e, sä	g->1	r->2	
e, så	 ->3	v->1	
e, ta	c->1	
e, ti	l->1	
e, to	g->1	
e, tr	o->1	
e, ty	 ->3	
e, tä	n->1	
e, tå	l->1	
e, un	d->2	
e, ur	 ->1	
e, ut	a->2	g->1	m->1	r->1	
e, va	r->6	
e, ve	t->1	
e, vi	 ->2	l->15	s->1	
e, vä	c->1	
e, vå	r->4	
e, än	d->1	
e, är	 ->9	a->1	
e, åt	e->4	
e, ök	a->1	
e- oc	h->6	
e- pr	o->1	
e-Alp	e->1	
e-Ard	e->1	
e-Atl	a->1	
e-Fra	n->2	
e-Le 	B->1	
e-Loi	r->1	
e-Man	n->1	
e-Nor	m->1	
e-alb	a->1	
e-avt	a->2	
e-avv	i->1	
e-dan	s->1	
e-de-	F->2	
e-dis	k->2	
e-fal	l->1	
e-fos	s->1	
e-för	s->1	
e-lob	b->1	
e-län	d->1	
e-mai	l->1	
e-met	a->1	
e-pro	g->2	
e-spr	i->3	
e-sta	t->9	
e-sti	p->1	
e-sto	p->1	
e. De	 ->1	t->4	
e. Dä	r->1	
e. Me	n->1	
e. Oc	h->1	
e. Om	 ->1	
e. Vi	 ->1	,->1	
e. Än	d->1	
e.- (	P->1	
e.- F	r->1	
e.. (	F->1	
e.. P	r->1	
e.. V	i->1	
e..(E	N->1	
e...)	.->1	
e.Akt	i->1	
e.All	t->2	
e.Ann	a->1	
e.Att	 ->2	
e.Av 	d->1	
e.Avs	l->2	
e.Bes	l->1	
e.Bet	ä->1	
e.Båd	a->1	
e.De 	e->1	
e.Den	 ->7	n->2	
e.Der	a->1	
e.Des	s->6	
e.Det	 ->55	t->11	
e.Där	e->1	f->7	
e.Då 	f->1	s->1	
e.Eft	e->5	
e.Eme	l->1	
e.En 	a->3	r->1	v->1	
e.End	a->1	
e.Enl	i->2	
e.Ett	 ->1	
e.Eur	o->4	
e.FPÖ	 ->1	
e.Fru	 ->4	
e.Frå	g->1	
e.För	 ->11	e->3	s->1	
e.Gen	o->2	
e.Gru	p->1	
e.Han	 ->2	
e.Hel	a->1	
e.Her	r->12	
e.Hon	 ->1	
e.Hur	 ->1	
e.Huv	u->4	
e.I E	u->1	
e.I d	a->2	e->1	
e.I o	c->1	
e.I s	i->1	t->1	
e.I v	a->1	i->1	
e.Idé	n->1	
e.Imm	i->1	
e.Inf	ö->1	
e.Ino	m->1	
e.Jag	 ->60	
e.Kan	 ->1	s->1	
e.Kom	m->7	
e.Lik	a->1	s->1	
e.Lyc	k->1	
e.Läg	g->1	
e.Låt	 ->4	
e.Mal	t->1	
e.Man	 ->6	n->1	
e.Med	 ->1	b->1	
e.Men	 ->16	
e.Mer	 ->1	
e.Min	 ->5	a->2	
e.Mån	g->1	
e.Ni 	k->3	s->1	
e.Nu 	b->1	f->1	
e.När	 ->3	
e.Och	 ->3	
e.Off	e->1	
e.Om 	d->2	k->1	n->1	r->1	v->2	
e.Par	a->1	
e.Pla	s->1	
e.Por	t->1	
e.Pro	b->1	d->1	
e.På 	d->2	
e.Ref	o->1	
e.Res	u->1	
e.Rot	h->1	
e.Råd	e->2	
e.Sam	t->1	
e.Sav	e->1	
e.Sch	u->1	
e.Sed	a->1	
e.Ska	l->1	
e.Slu	t->2	
e.Som	 ->7	l->1	
e.Stä	m->1	
e.Stö	r->1	
e.Så 	f->1	n->1	
e.Sål	e->1	
e.TV-	b->1	
e.Ta 	d->1	
e.Tac	k->3	
e.Til	l->3	
e.Top	p->1	
e.Tra	n->1	
e.Tro	t->1	v->1	
e.Tvä	r->1	
e.Und	a->1	e->1	
e.Upp	f->1	
e.Ur 	d->1	
e.Vad	 ->2	a->1	
e.Var	 ->1	e->1	f->1	
e.Vi 	a->1	b->2	f->3	h->2	i->1	k->4	m->3	r->1	s->2	v->2	ä->2	
e.Vid	 ->2	
e.Vin	d->1	
e.Vit	b->1	
e.Vår	 ->3	
e.d.,	 ->1	
e.Änd	r->2	
e.Är 	d->1	
e.Äve	n->2	
e.Å a	n->1	
e.År 	1->1	
e.Åte	r->1	
e.Åtg	ä->1	
e.Öst	e->1	
e: "A	t->1	
e: "v	a->1	
e: An	l->1	
e: Ar	b->1	t->1	
e: De	t->2	
e: Fl	o->1	
e: Fr	ä->1	
e: Fö	r->1	
e: Ge	m->1	n->1	
e: Gr	e->1	
e: Ha	n->1	
e: I 	m->1	
e: Ja	g->1	
e: Jo	r->1	
e: Ko	c->1	m->1	
e: Kä	r->1	
e: Ma	i->1	
e: Na	r->1	
e: Ny	t->1	
e: Nä	r->1	
e: Po	r->1	
e: St	a->1	ö->1	
e: Tu	r->1	
e: Ut	n->1	
e: Va	d->1	p->1	
e: Vi	 ->2	
e: ba	l->1	
e: be	s->1	
e: de	t->1	
e: fö	r->1	
e: hu	r->1	
e: i 	l->1	r->1	
e: ko	m->1	
e: to	l->1	
e: ut	v->1	
e: va	r->1	
e: Åt	g->2	
e; de	n->1	t->1	
e; hä	r->1	
e; ja	g->1	
e; mi	n->1	
e; pu	n->1	
e?Den	 ->1	
e?Det	 ->1	
e?Enl	i->1	
e?För	 ->2	
e?Hem	l->1	
e?Her	r->3	
e?Hur	 ->1	
e?Här	m->1	
e?I f	j->1	
e?Jag	 ->1	
e?Kan	s->1	
e?Och	 ->1	
e?Som	 ->1	
e?Vi 	ä->1	
e?Vil	k->1	
eEn v	ä->1	
eFru 	t->1	
eHerr	 ->1	
eNäst	a->2	
eProt	o->1	
ea be	h->1	
ea oc	h->3	
ead-k	o->1	
eader	 ->3	,->1	-->1	
eadin	g->1	
eadli	n->1	
eager	a->16	
eake,	 ->1	
eakt 	o->1	
eakta	 ->9	d->1	n->4	r->3	s->8	t->5	
eakti	o->12	
eakto	r->10	
eal p	r->1	
eal, 	a->1	h->1	
eala 	s->1	
ealen	 ->1	
ealet	 ->1	
ealis	m->1	t->9	
ealit	e->7	
eamin	g->8	
ean-C	l->1	
eanut	s->1	
earbe	t->3	
earve	t->1	
eater	g->1	
eativ	a->2	
eato 	-->1	f->2	h->1	o->1	s->2	t->1	
eato.	J->1	
eatob	e->1	
eaton	-->1	
eatos	 ->11	
eattl	e->4	
eatör	e->1	
eau d	u->1	
eau f	ö->1	
eau",	 ->1	
eau, 	a->1	o->1	
eaux,	 ->1	
eb, s	o->1	
eball	m->1	
ebano	r->1	
ebar 	f->1	
ebase	n->1	
ebast	i->1	
ebatt	 ->53	,->9	.->21	:->1	?->1	B->1	e->82	i->1	k->1	
ebbel	s->1	
ebbpl	a->1	
ebefo	r->2	
ebefr	a->1	
ebeha	n->1	
ebeng	a->1	
ebest	ä->3	
ebesö	k->1	
ebeta	l->12	
ebild	,->1	
eboar	d->1	
eboel	i->1	
eboen	d->1	
ebola	g->4	
eborg	 ->1	
ebrei	s->1	
ebron	-->1	
ebrua	r->16	
ebrås	 ->2	
ebröd	.->1	
ebud 	f->4	v->1	ä->1	
ebud,	 ->2	
ebude	t->1	
ebygd	 ->1	
ebygg	a->22	e->2	
ebält	e->10	
ebänk	e->1	
ebär 	a->46	b->1	d->4	e->15	f->3	i->9	m->2	n->1	o->4	p->1	s->2	ä->1	ö->1	
ebär,	 ->1	
ebär.	D->1	F->1	
ebära	 ->15	
ebåda	d->1	
ebörd	.->1	e->6	
ebörs	e->1	
ec l'	e->1	
ecedo	 ->1	
ecemb	e->19	
ecenn	i->7	
ecent	r->15	
ecial	b->2	d->1	f->2	i->7	p->1	u->1	
eciel	l->42	
ecifi	c->2	k->27	
ecirk	u->1	
ecis 	d->4	e->1	f->1	h->1	i->1	l->5	p->1	s->21	v->1	
ecisa	 ->1	
ecise	r->11	
ecist	 ->1	
eck h	a->1	
eck i	n->1	
eck ä	r->1	
ecka 	h->2	i->1	r->1	s->1	ä->1	
ecka.	(->1	
eckan	 ->17	
ecken	 ->13	.->2	
eckla	 ->31	d->10	n->3	r->2	s->21	t->6	
eckli	n->175	
eckna	 ->3	d->6	n->1	r->2	s->6	t->11	
eckni	n->3	
eckor	 ->8	,->1	.->1	n->7	
ecove	r->1	
ectne	s->1	
ecu m	e->1	
ecu, 	e->1	
ecycl	i->1	
ed "a	l->1	n->1	
ed "e	n->1	
ed (a	t->1	
ed - 	o->1	
ed 12	 ->1	
ed 13	 ->2	
ed 14	,->1	
ed 16	4->1	
ed 19	9->1	
ed 2 	m->1	p->1	
ed 20	 ->1	0->1	
ed 24	 ->1	
ed 27	 ->2	
ed 28	 ->1	
ed 30	 ->1	
ed 36	7->1	
ed 5 	0->1	
ed 80	 ->1	
ed A.	 ->1	
ed Am	o->1	s->1	
ed BS	E->1	
ed Ba	l->1	
ed Da	l->1	v->1	
ed E-	k->1	
ed ED	D->1	
ed EU	-->1	
ed Er	i->4	
ed Eu	r->12	
ed Fr	a->4	
ed GA	-->1	
ed Ha	a->1	i->3	
ed In	t->1	
ed Is	l->1	r->1	
ed Jö	r->1	
ed Ko	u->2	
ed Le	a->1	
ed Li	b->1	t->1	
ed Ma	a->1	d->1	l->1	
ed Mi	d->1	
ed OL	A->1	
ed Os	l->1	
ed Pa	t->1	
ed Ry	s->1	
ed Sa	v->1	
ed Sy	d->1	r->3	
ed Th	e->1	
ed Tu	r->2	
ed US	A->4	
ed Va	n->1	
ed Ve	r->1	
ed ad	m->1	
ed al	l->33	t->1	
ed an	d->13	g->1	k->1	l->4	n->1	s->6	t->1	v->1	
ed ar	b->4	g->1	t->7	
ed at	t->106	
ed au	t->2	
ed av	 ->1	s->15	t->1	
ed ba	l->1	r->1	s->1	
ed be	d->2	g->1	k->3	v->1	
ed bi	b->1	d->2	l->2	
ed br	a->1	i->3	o->1	y->1	å->1	
ed bu	d->1	
ed bå	d->1	
ed da	g->3	t->1	
ed de	 ->67	l->3	m->13	n->82	r->3	s->22	t->56	
ed di	r->7	s->1	
ed dr	a->1	o->1	
ed du	b->2	
ed dy	l->1	s->1	
ed ef	t->2	
ed ek	o->1	
ed el	l->1	
ed en	 ->81	a->1	b->1	h->4	o->1	t->1	
ed er	 ->7	.->2	a->3	b->1	
ed et	t->29	
ed eu	r->2	
ed ex	i->1	k->1	p->3	
ed fa	r->3	t->1	
ed fe	d->1	
ed fi	n->1	
ed fl	e->3	
ed fo	n->1	r->2	
ed fr	a->4	i->14	u->1	å->11	
ed fu	l->3	n->6	
ed få	 ->1	
ed fö	l->1	r->37	t->1	
ed ga	m->1	
ed ge	m->4	n->3	
ed gi	g->1	
ed gl	ä->2	
ed go	d->5	
ed gr	a->1	u->2	ö->1	
ed ha	m->1	n->2	
ed he	m->2	n->1	
ed hj	ä->25	
ed ho	n->1	
ed hu	n->1	r->4	
ed hä	n->18	
ed hå	l->1	
ed hö	g->2	
ed i 	M->3	b->2	d->8	e->2	k->1	m->2	p->1	r->1	s->2	t->1	u->3	ä->1	
ed if	r->1	
ed im	p->1	
ed in	f->3	h->1	n->1	o->1	r->2	s->5	t->10	
ed is	 ->2	
ed jo	r->1	
ed ju	l->1	
ed jä	m->1	
ed ka	n->3	p->1	t->1	
ed ki	n->1	
ed kl	a->1	
ed kn	a->1	
ed ko	l->1	m->22	n->7	s->1	
ed kr	a->5	i->2	
ed ku	n->1	
ed kv	a->8	i->1	
ed kä	r->1	
ed kö	p->1	
ed la	g->2	n->1	
ed le	d->1	g->1	
ed li	g->1	k->3	n->1	v->3	
ed lä	m->1	
ed lö	s->2	
ed ma	j->1	n->1	r->3	t->1	
ed me	d->12	l->1	r->2	
ed mi	g->5	k->2	l->5	n->17	t->1	
ed mo	n->1	r->2	t->2	
ed my	c->6	
ed må	l->2	n->3	s->2	
ed mö	j->3	t->1	
ed na	m->4	t->8	z->1	
ed ne	g->3	
ed nu	 ->2	m->1	
ed ny	a->1	f->1	k->1	t->1	
ed nä	r->1	
ed nå	g->8	
ed nö	d->4	j->2	t->1	
ed oc	h->14	k->4	
ed of	f->1	
ed oj	ä->1	
ed ol	i->2	
ed om	 ->17	.->1	b->1	s->4	
ed or	d->4	m->1	o->1	
ed os	s->7	ä->1	
ed pa	l->1	r->12	
ed pe	n->3	r->2	
ed pl	a->1	
ed po	l->3	
ed pr	i->3	o->5	
ed ps	y->1	
ed pu	n->2	
ed på	 ->18	l->1	
ed ra	d->1	
ed re	d->2	f->2	g->2	k->1	p->3	s->9	
ed ri	k->2	
ed rä	t->10	
ed rå	d->5	
ed rö	t->1	
ed s.	k->1	
ed sa	k->2	m->8	
ed se	k->1	
ed si	f->1	g->8	n->11	t->6	
ed sj	ä->1	
ed sk	a->3	j->1	u->2	y->1	
ed sl	a->1	u->1	
ed sm	å->1	
ed sn	e->1	
ed so	c->5	m->2	
ed sp	e->2	ä->3	
ed st	a->4	i->1	o->21	r->5	ö->6	
ed su	b->2	
ed sv	ä->1	å->1	
ed sy	f->2	
ed sä	g->1	k->4	l->1	r->3	
ed så	 ->3	,->1	d->7	
ed t.	e->1	
ed ta	c->1	n->42	
ed te	k->1	x->1	
ed ti	d->9	l->13	
ed to	l->1	
ed tr	a->1	e->5	
ed tu	n->1	r->1	
ed tv	i->1	å->4	
ed ty	p->1	
ed tä	t->1	
ed un	d->3	g->1	i->2	
ed up	p->6	
ed ur	s->1	
ed ut	a->4	b->2	g->1	s->7	v->3	
ed va	d->5	l->1	r->7	
ed ve	r->3	t->3	
ed vi	 ->1	l->8	s->6	t->2	
ed vä	l->1	
ed vå	r->17	
ed yr	k->1	
ed yt	t->4	
ed ÖV	P->1	
ed Ös	t->1	
ed än	d->4	
ed är	 ->4	e->1	
ed år	 ->1	e->1	
ed åt	a->2	g->2	
ed ök	n->1	
ed öm	s->1	
ed öp	p->1	
ed ös	t->1	
ed öv	e->9	r->2	
ed, a	t->1	
ed, d	e->1	ä->1	
ed, e	f->1	
ed, f	r->1	
ed, g	ö->1	
ed, m	e->2	
ed, n	ä->1	
ed, o	c->1	m->2	
ed, p	r->1	
ed, s	å->1	
ed, v	a->1	
ed.De	n->1	t->3	
ed.Dä	r->1	
ed.Ef	f->1	
ed.Fö	r->1	
ed.He	r->1	
ed.Hu	r->1	
ed.I 	T->1	
ed.Ja	g->1	
ed.Ko	m->1	
ed.Vi	 ->2	
eda E	u->1	
eda a	l->1	n->2	
eda d	e->4	i->1	
eda e	n->6	t->2	
eda f	o->1	r->1	ö->4	
eda h	u->1	
eda i	n->2	
eda m	e->1	i->1	y->1	ö->1	
eda o	c->1	d->1	s->2	
eda p	r->1	å->3	
eda s	i->2	
eda t	i->30	
eda u	t->3	
eda å	t->1	
eda, 	p->1	t->1	v->1	
edago	g->1	
edakt	i->1	
edamo	t->74	
edamö	t->84	
edan 	1->15	4->1	A->1	E->1	F->1	P->1	S->1	a->13	b->9	d->25	e->15	f->20	g->10	h->41	i->17	j->3	k->7	l->5	m->5	n->9	o->4	p->8	r->4	s->19	t->19	u->7	v->13	ä->7	å->1	ö->1	
edan,	 ->11	
edan.	D->4	H->1	I->1	J->3	S->1	
edan?	 ->1	S->1	
edand	e->18	
edans	v->3	
edarb	e->2	
edare	 ->8	,->1	n->2	s->2	
edarf	ö->1	
edarn	a->8	
edars	k->1	
edas 	a->2	d->1	m->1	t->1	u->1	
edas,	 ->1	
edast	 ->1	
edat 	f->1	
edbes	l->16	
edbor	g->170	
edbro	t->1	
edd a	t->16	
edd f	ö->2	
edd t	i->3	
edd u	t->2	
edd ä	n->1	
edda 	a->13	e->1	l->1	r->2	t->1	
edda.	M->1	
edde 	A->1	d->1	e->1	f->4	t->7	
edde,	 ->1	
eddel	a->59	
edden	 ->1	,->1	
eddes	 ->6	.->1	
ede g	e->1	
ede o	c->1	
ede ä	r->1	
ede.R	e->1	
edel 	(->2	K->1	a->10	b->2	f->15	m->1	n->1	o->9	p->1	s->11	t->3	u->2	ä->3	
edel,	 ->12	
edel.	D->3	J->1	N->1	S->1	V->3	
edel?	J->1	
edela	r->4	
edelb	a->18	
edelh	a->3	
edell	å->4	
edelp	u->2	
edels	-->1	e->6	f->2	h->1	i->2	k->5	l->5	m->9	n->1	p->2	s->45	t->42	
edelt	i->1	
eden 	a->1	
eden,	 ->1	
edens	 ->1	
edepa	r->2	
eder 	b->1	d->3	e->6	f->6	h->1	i->3	k->1	n->3	o->4	r->1	s->1	t->16	u->1	v->1	
eder,	 ->2	
edera	l->10	t->2	
ederb	ö->11	
ederg	ä->1	
ederi	e->2	
ederl	ä->18	
eders	a->1	
edert	a->1	
ederv	ä->1	
edes 	a->4	b->4	d->1	e->3	f->2	g->1	h->4	i->3	k->3	l->1	n->3	o->1	p->3	r->2	s->2	t->2	u->1	v->2	ä->2	
edet 	l->1	s->1	t->1	
edfin	a->2	
edför	 ->10	,->2	a->4	d->1	e->2	t->1	
edgat	 ->1	
edge 	F->1	a->3	
edger	 ->10	
edges	 ->5	
edget	t->1	
edgiv	i->2	
edgån	g->2	
edgör	l->2	
edhjä	l->1	
edi -	 ->1	
edi.D	e->1	
edia 	-->1	a->1	h->1	s->2	
edial	 ->1	
edias	 ->1	
ediat	ä->1	
edici	n->1	
edien	s->2	
edier	 ->3	.->2	n->2	
edige	n->1	
edigh	e->1	
edign	a->1	
edinf	l->1	
eding	 ->4	,->3	s->1	
edite	r->2	
editi	o->1	
edja 	a->1	
edjan	 ->2	
edje 	a->1	b->2	d->2	f->2	g->3	l->24	m->4	o->2	p->6	r->2	s->1	v->4	ä->1	å->1	ö->1	
edje,	 ->4	
edje:	 ->1	
edjed	e->6	
edjel	a->6	
edjor	n->1	
edkvi	s->1	
edkän	s->5	
edla 	v->2	
edlag	d->1	
edlar	 ->1	
edlem	 ->5	,->1	m->14	s->323	
edlen	 ->10	,->2	
edlet	 ->1	
edlid	a->2	
edlig	 ->5	a->2	h->2	t->1	
edlin	g->2	
edläg	g->4	
edmon	t->3	
ednin	g->83	
edo a	n->1	t->3	
edofi	l->1	
edogj	o->1	
edogö	r->9	
edom 	o->2	
edom,	 ->2	
edoma	r->4	
edome	n->4	
edovi	s->4	
edra 	a->2	d->1	o->2	
edrad	e->1	
edrag	,->1	a->110	i->1	n->48	
edran	d->3	
edrar	 ->3	
edrev	s->1	
edriv	a->6	e->3	s->6	
edrog	 ->1	
edrus	t->1	
edräg	e->36	l->1	
eds a	t->1	
eds b	l->1	
eds i	 ->1	
eds m	e->1	
eds r	e->1	
eds s	a->1	
eds u	n->1	
eds å	r->1	
eds, 	m->1	
eds.J	a->1	
edsan	s->1	
edsav	t->3	
edsbe	s->1	v->1	
edsen	 ->1	,->1	
edsfö	r->3	
edska	p->2	
edskr	ä->1	
edskä	r->3	
edspa	r->1	
edspr	o->22	
edssa	m->4	
edsst	ä->24	
edstj	ä->2	
edstä	m->1	n->2	
edsup	p->1	
edt o	c->2	
edt, 	f->1	i->1	
edter	 ->5	,->1	H->1	b->2	s->5	
educe	r->4	
edurr	e->1	
edver	k->19	
edvet	a->4	e->21	n->17	
edvri	d->12	
edvär	d->1	
edöma	 ->12	,->1	s->2	
edömb	a->1	
edömd	e->1	
edöme	r->4	
edöml	i->2	
edömn	i->28	
edöms	 ->3	
edömt	 ->1	
ee-fö	r->1	
ee-lo	b->1	
ee.De	t->1	
eelan	d->2	
eell 	r->1	
eell.	F->1	
eella	 ->4	
eende	 ->27	,->4	.->4	:->1	;->1	n->13	t->13	
eenhe	t->5	
eer o	m->1	
eer s	a->1	o->1	
eer, 	T->1	f->1	s->2	
eerJa	g->1	
eerbe	t->3	
eerin	g->1	
eers 	b->3	
eersä	t->2	
ees W	i->1	
eexem	p->1	
ef ha	r->1	
efade	r->1	
efall	e->20	
efant	 ->1	
efara	 ->2	r->3	
efatt	a->10	n->2	
efel 	o->1	
efen 	D->1	
efer 	o->3	p->1	
efer,	 ->2	
efer.	O->1	
efere	n->4	r->3	
efern	a->8	
effek	t->148	
effic	i->1	
efing	-->1	
efini	e->13	t->23	
efinn	a->3	e->28	
efint	l->10	
efit-	a->5	
eflek	t->7	
efläc	k->1	
efoga	d->2	t->3	
efoge	n->27	
efolk	a->1	n->42	
efon,	 ->1	
efond	e->1	
eford	r->8	
eform	 ->27	,->7	.->5	:->1	a->4	e->77	f->2	i->1	p->15	s->1	å->1	
efrak	t->10	
efria	 ->1	s->3	
efrie	l->6	
efrih	e->2	
efräm	j->1	
efråg	o->2	
efter	 ->145	,->1	.->2	;->1	b->1	f->11	g->8	h->5	l->6	m->9	s->177	t->6	å->1	
efull	 ->2	.->2	a->7	t->7	
efuse	"->1	
efusi	o->1	
efälh	a->1	
efäng	d->1	
efär 	1->3	7->1	l->1	s->2	t->2	
efärl	i->1	
efäst	 ->1	a->5	e->4	
eföll	 ->1	
eförb	e->1	
eföre	s->4	t->2	
eförf	a->8	
eförh	å->3	
eförk	l->1	
eföro	r->1	
eförs	k->1	
eförv	a->1	
eg at	t->1	
eg bo	r->1	
eg fr	a->5	å->1	
eg fö	r->5	
eg gj	o->1	
eg ha	r->1	
eg hä	r->1	
eg i 	M->1	a->1	d->1	f->2	k->1	r->3	s->2	u->1	v->1	
eg jä	m->1	
eg lä	n->2	
eg mo	t->4	
eg nä	r->2	
eg oc	h->2	
eg på	 ->3	
eg so	m->7	
eg te	r->1	
eg ti	l->3	
eg un	d->1	
eg vi	 ->1	
eg, d	ä->1	
eg, o	c->1	
eg, u	t->1	
eg.De	t->2	
ega B	e->2	o->1	
ega E	l->1	v->1	
ega F	i->1	l->3	r->2	
ega H	u->1	
ega J	a->1	e->1	o->1	
ega K	o->1	
ega L	i->1	
ega M	u->1	
ega N	a->1	i->1	
ega R	a->1	o->1	
ega S	a->1	
ega a	n->1	
ega b	e->1	
ega d	e->1	
ega f	r->2	
ega k	o->1	
ega s	a->1	o->1	
ega t	i->1	
ega v	a->4	
ega! 	V->1	
ega!D	e->1	
ega!J	a->1	
ega!Ä	v->1	
ega, 	E->1	a->2	
ega.J	a->1	
egad.	V->1	
egade	 ->1	
egagn	a->4	
egal 	i->1	p->2	s->1	
egala	 ->7	
egali	s->1	t->1	
egalt	 ->9	
egan 	B->2	D->1	J->1	K->2	L->1	N->1	P->1	S->1	W->3	f->1	v->2	
egapr	o->1	
egas 	i->1	k->1	
egat 	e->1	f->1	n->1	
egati	o->16	v->26	
egdra	g->1	
ege.O	m->1	
ege?H	e->1	
egel 	r->1	ä->2	
egelb	r->1	u->15	
egelm	ä->2	
egeln	 ->6	
egelr	ä->2	
egels	y->2	
egelv	e->19	
egeme	n->3	
egen 	b->1	d->5	f->1	g->2	h->2	i->2	k->4	o->3	p->2	r->4	s->4	u->1	v->1	ä->1	ö->1	
egena	n->1	
egend	o->5	
egene	r->1	
egenf	ö->5	
egens	k->22	
egent	l->43	
eger 	a->5	b->2	f->4	h->1	i->7	k->1	m->2	o->2	r->1	s->4	t->2	u->1	v->4	
eger!	 ->58	D->3	E->1	J->2	V->1	
eger,	 ->14	
eger.	A->1	D->1	H->1	J->2	
eger:	 ->1	
egera	 ->2	s->1	t->1	
egeri	n->288	
egern	 ->1	a->8	
egers	 ->1	
eget 	a->2	g->2	h->2	i->2	k->1	l->2	m->1	o->1	p->3	r->1	s->2	t->1	v->1	y->1	ä->1	ö->1	
eget,	 ->2	
eget.	D->1	
egi f	ö->5	
egi h	a->1	
egi i	 ->1	
egi k	a->1	
egi m	å->1	
egi o	c->2	
egi s	o->4	
egi t	i->2	
egi, 	d->1	e->1	i->1	m->1	
egi.D	e->1	
egi.F	r->1	
egi.J	a->1	
egick	 ->1	
egier	 ->11	,->4	.->1	n->1	
egiet	,->1	.->1	
egime	n->3	
egin 	f->1	k->1	m->1	o->1	s->1	
egin.	D->1	S->1	
egins	 ->1	
egion	 ->12	,->3	.->7	a->89	e->141	
egipl	a->1	
egisk	 ->3	a->10	t->4	
egist	e->10	r->10	
egiti	m->18	
egium	 ->2	.->1	
egla 	d->2	m->1	p->4	
eglad	e->2	
eglar	 ->11	,->1	.->1	
eglas	 ->2	
egler	 ->39	,->10	.->6	?->1	a->19	i->15	n->36	
eglin	g->1	
egna 	a->1	b->2	e->1	f->9	i->5	k->2	m->4	n->3	o->1	p->3	r->1	s->9	v->2	å->2	
egni,	 ->1	
egois	t->2	
egor 	F->1	
egori	 ->3	e->5	s->1	
egors	 ->2	
egrad	e->3	
egrat	 ->1	i->16	
egrav	a->1	
egrep	p->13	
egrer	a->17	i->6	
egrip	a->2	e->13	l->6	n->1	
egrit	e->3	
egrun	d->2	
egrän	s->68	
eguro	,->1	
egär 	a->3	b->1	d->1	e->3	o->1	s->1	ö->1	
egär.	V->1	
egära	 ->9	,->1	n->21	s->3	
egärd	e->3	
egärs	 ->1	
egärt	 ->7	,->2	.->1	
egå e	n->1	
egå s	å->1	
egåen	d->15	
egång	a->3	s->1	
egår 	b->3	
egås 	a->1	i->1	o->1	
egått	 ->2	s->1	
ehabi	l->1	
ehagl	i->2	
ehand	a->3	l->85	
ehar 	c->1	e->1	
ehava	n->1	r->1	
ehind	r->1	
ehov 	a->15	i->1	k->1	o->4	s->2	
ehov,	 ->2	
ehov.	A->1	H->1	U->1	
ehove	n->5	t->34	
ehren	d->7	
ehäft	a->1	
ehåll	 ->9	,->2	.->5	?->1	a->29	e->57	i->3	s->14	
ehöja	n->1	
ehöll	 ->4	s->1	
ehöri	g->18	
ehöva	 ->15	s->1	
ehövd	e->2	
ehöve	r->99	
ehövs	 ->20	,->2	.->5	
ehövt	 ->2	s->1	
eidos	k->2	
eijs 	o->1	
eijs.	(->1	
eik.D	e->1	
eikh 	h->1	
eikh-	a->1	
eikh.	D->1	F->1	
eille	 ->1	
ein.J	a->1	
einci	t->1	
eindr	ä->2	
eindu	s->1	
einen	 ->3	,->2	s->1	
einsp	e->1	
einst	e->2	
einz 	F->2	
eira 	R->1	ä->1	
eira,	 ->2	
eira.	J->1	
eiser	a->1	i->1	
eisk 	a->9	b->6	c->2	d->2	f->1	g->1	h->2	i->6	j->3	k->11	l->9	m->5	n->13	o->4	p->4	r->3	s->5	u->3	å->13	
eisk.	H->1	
eiska	 ->585	.->1	
eiske	 ->2	
eiskt	 ->20	
eismi	s->2	
eivra	s->1	
eixas	 ->5	
eiz, 	t->1	
ej an	g->1	
ej at	t->1	
ej av	g->1	
ej be	r->1	s->1	
ej bo	r->1	
ej i 	f->1	
ej ko	m->1	
ej lå	n->1	
ej lö	s->1	
ej nä	r->1	
ej ti	l->1	
ej är	 ->1	
ej, b	e->1	i->1	
ej, d	e->1	
ej, h	e->1	
ej, j	a->1	
ej, m	a->2	
ej, n	a->1	
ej, s	k->1	ä->1	
ej.(A	p->1	
ej.Ex	p->1	
ej.I 	s->1	
ej.Rå	d->1	
ejda 	m->1	
ejdas	 ->1	
ejdat	 ->1	
ejdos	k->1	
ejord	b->3	
ejudi	c->1	k->3	
ejält	 ->3	
ek ho	n->1	
ek os	s->1	
ek so	m->1	
eka B	a->1	
eka a	t->9	
eka d	e->4	
eka f	ö->5	
eka p	å->6	
eka r	å->1	
eka v	i->1	
eka, 	d->1	h->1	
eka.D	e->1	
eka.M	i->1	
ekad 	r->1	
ekade	 ->7	,->1	.->2	s->1	
ekan 	a->1	d->1	e->2	f->1	h->1	k->2	m->1	o->2	s->2	ä->1	
ekan,	 ->1	
ekand	e->11	
ekani	k->1	s->9	
ekant	 ->1	,->2	
ekar 	T->1	a->4	b->1	h->1	i->4	m->1	o->1	p->1	s->1	u->1	
ekar,	 ->1	
ekas 	a->2	k->1	o->1	t->1	
ekas,	 ->1	
ekast	e->1	
ekat 	-->1	a->2	f->1	h->1	o->1	p->4	u->1	
ekat,	 ->4	
ekat.	Ö->1	
ekel 	a->1	k->1	
ekel,	 ->1	
ekels	k->1	
eken 	i->1	v->1	
eken,	 ->1	
ekens	 ->1	
eker 	m->1	
ekern	a->1	
ekhet	 ->2	,->1	e->1	
eking	 ->1	
ekisk	a->6	
ekist	a->2	
eklag	a->34	l->8	
eklam	 ->2	
eklan	d->14	g->1	
ekler	n->1	
eklet	 ->1	
eklös	t->1	
eknik	 ->6	e->7	
eknis	k->36	
eknol	o->3	
ekod 	f->5	
ekode	n->1	r->2	
ekoka	 ->1	
ekoll	e->1	
ekolo	g->14	
ekom 	o->1	p->1	
ekomm	a->5	e->54	i->6	u->3	
ekomp	l->1	
ekoms	t->1	
ekon 	a->1	
ekonc	e->1	
ekonf	e->2	
ekono	m->283	
ekons	t->3	
ekonv	e->1	
ekord	 ->1	t->1	
ekort	 ->1	
ekost	n->1	
ekosy	s->4	
ekret	a->2	e->14	
ekris	 ->1	
ekryt	e->1	
ekräf	t->30	
eksak	e->1	
eksam	 ->1	h->2	m->1	t->1	
ekt a	n->1	t->5	v->2	
ekt b	a->1	e->3	i->1	y->1	
ekt d	r->1	
ekt e	l->1	r->2	
ekt f	a->1	r->1	å->1	ö->25	
ekt g	å->1	
ekt h	a->3	
ekt i	 ->1	n->2	
ekt k	a->1	l->1	o->2	
ekt l	ä->2	
ekt m	a->1	e->4	o->2	
ekt n	ä->1	
ekt o	c->4	m->1	
ekt p	o->1	å->2	
ekt s	a->2	k->1	m->1	o->13	t->2	v->1	ä->3	
ekt t	i->8	
ekt u	p->1	t->2	
ekt v	a->1	i->2	
ekt ä	r->1	
ekt",	 ->1	
ekt, 	e->2	f->1	n->1	u->1	v->3	
ekt.D	e->3	å->1	
ekt.F	e->1	ö->1	
ekt.I	 ->1	
ekt.J	a->1	
ekt.M	a->1	å->1	
ekt.S	l->1	
ekt.U	n->1	
ekt: 	u->1	
ekt; 	e->1	
ekt?T	ä->1	
ekt?U	t->1	
ekta 	a->1	b->2	e->1	g->1	s->4	v->1	
ekta.	J->1	
ektab	e->2	i->1	
ektad	m->2	
ektak	e->2	u->1	
ektar	 ->2	
ekten	 ->31	,->1	.->6	
ekter	 ->23	,->7	.->4	a->38	n->7	
ektet	 ->12	,->1	s->1	
ektin	v->1	
ektio	n->18	
ektiv	 ->114	,->15	.->13	:->2	?->2	a->41	e->109	f->3	i->26	t->29	
ektor	 ->8	,->4	.->3	a->18	e->19	i->1	n->49	p->1	s->4	
ektri	c->1	
ektro	n->9	
ektru	m->2	
ektue	l->3	
ektyr	.->1	
ektör	,->1	e->5	s->1	
ekula	t->4	
ekund	e->2	ä->1	
ekval	i->1	
ekvat	 ->3	a->2	i->1	
ekven	s->46	t->16	
ekvot	e->1	
ekväm	l->15	t->1	
ekymm	e->6	
ekymr	a->10	
ekämp	a->29	n->12	
ekänn	e->1	
el (k	o->2	
el - 	d->2	s->1	u->1	ö->1	
el 1 	i->1	u->1	
el 10	5->1	
el 11	0->1	
el 12	 ->1	,->1	
el 13	 ->4	.->1	
el 14	3->1	
el 15	8->3	
el 16	)->1	
el 2.	1->1	2->1	
el 22	6->1	
el 25	5->4	
el 28	0->5	
el 29	9->2	
el 3.	1->1	8->1	
el 30	 ->1	
el 33	 ->2	
el 37	 ->1	.->1	
el 39	 ->1	
el 4 	c->1	i->4	
el 4.	2->1	
el 42	 ->1	
el 48	 ->2	
el 5 	g->1	
el 5.	4->1	
el 50	 ->1	,->1	
el 52	 ->1	
el 56	,->1	
el 6 	i->6	o->3	
el 6.	S->1	
el 62	 ->1	
el 67	 ->1	
el 7 	i->6	n->1	
el 7,	 ->1	
el 81	 ->1	.->9	
el 82	,->1	.->1	
el 87	.->2	
el 88	 ->2	
el 9.	1->1	
el 94	 ->1	
el 95	 ->1	
el Ba	s->1	
el Hi	l->1	
el Ko	u->1	
el Ny	a->1	
el Pe	a->1	
el Ri	o->1	
el al	d->1	l->1	
el an	d->1	g->1	m->1	s->1	v->1	
el at	t->14	
el av	 ->81	,->1	s->1	
el be	f->1	g->1	r->1	v->1	
el bl	a->1	
el bä	s->1	
el bö	r->2	
el de	 ->1	l->6	t->1	
el dr	a->1	
el en	k->1	
el et	t->1	
el fa	l->2	r->1	s->1	
el fo	r->1	
el fr	i->1	ä->1	å->3	
el få	 ->1	
el fö	r->28	
el ga	n->1	
el ge	n->2	t->1	
el gö	r->1	
el ha	r->5	
el hi	n->1	
el hj	ä->1	
el hy	c->1	
el hä	l->1	n->1	
el i 	V->1	a->3	d->6	e->1	f->2	g->1	m->1	s->1	u->1	v->2	ä->1	
el in	o->1	s->2	t->2	
el ka	n->4	
el ko	m->3	
el kv	i->1	ä->1	
el le	t->1	
el li	g->1	
el lö	p->1	s->1	
el ma	k->1	
el me	d->5	n->1	r->2	
el må	s->2	
el ni	 ->1	v->1	
el nu	 ->1	
el ny	t->1	
el nä	r->3	
el oc	h->36	k->1	
el om	 ->10	,->1	
el pa	r->1	
el pe	l->1	n->1	
el po	s->1	
el på	 ->24	,->1	.->1	
el ra	d->1	
el re	t->1	
el ri	s->1	
el rä	c->1	
el rö	r->1	
el sa	k->1	m->2	
el se	t->1	
el si	g->1	
el sk	a->3	u->1	
el so	m->17	
el st	e->1	
el sä	k->2	t->1	
el så	 ->1	
el ti	l->7	
el to	l->1	
el tr	ä->1	
el un	d->3	
el up	p->1	
el ur	 ->1	
el ut	a->1	f->1	
el va	n->1	r->1	
el ve	r->1	t->1	
el vi	l->1	s->1	
el än	 ->1	d->1	
el är	 ->15	
el äv	e->1	
el åt	e->1	
el öv	e->1	
el! I	n->1	
el! J	a->1	
el!Me	n->1	
el!Ti	l->1	
el, A	n->1	
el, a	n->1	t->2	
el, d	e->1	ä->1	å->1	
el, e	f->1	l->2	t->1	
el, f	o->1	ö->1	
el, i	 ->2	
el, j	u->1	
el, k	o->3	
el, l	i->1	ä->1	
el, m	e->7	
el, n	i->1	ä->2	
el, o	c->9	m->1	
el, s	o->4	å->1	
el, u	t->1	
el, v	a->1	i->3	
el, ä	v->1	
el, å	n->1	
el, ö	v->1	
el- o	c->3	
el-I)	;->1	
el-II	)->1	
el-Sh	e->5	
el-Sy	r->1	
el.Be	t->1	
el.De	n->1	t->10	
el.Dä	r->1	
el.EU	-->1	
el.Ef	t->1	
el.Eu	r->1	
el.Fr	a->1	
el.Ge	n->1	
el.I 	s->1	
el.Ja	g->4	
el.Me	n->4	
el.Nä	r->2	
el.Sa	m->1	
el.Sc	h->1	
el.Så	 ->1	
el.Tv	å->1	
el.Vi	 ->10	
el.Än	d->1	
el.Är	 ->1	
el: E	u->1	
el: F	i->1	
el: U	n->1	
el: V	e->1	
el: d	e->1	
el; i	 ->1	
el?El	l->1	
el?Ja	g->1	
ela 9	0->1	
ela B	a->1	
ela E	U->2	u->17	
ela K	o->1	
ela M	e->1	
ela S	u->1	
ela a	n->1	r->1	t->6	
ela b	e->1	ö->1	
ela d	e->18	i->2	
ela e	l->3	n->9	r->1	
ela f	l->1	r->4	ö->3	
ela g	e->3	
ela h	a->2	
ela i	 ->2	d->1	n->3	
ela k	o->11	
ela l	i->1	ä->1	
ela m	a->1	e->1	
ela n	ä->1	
ela o	c->2	f->1	
ela p	l->1	å->1	
ela r	e->4	
ela s	i->1	k->2	p->1	t->1	y->1	
ela t	e->1	i->9	y->1	
ela u	n->6	t->3	
ela v	e->1	ä->4	å->1	
ela å	r->1	t->2	
ela, 	h->1	
ela?A	v->1	
elad,	 ->1	
elade	 ->7	s->4	
elag 	o->1	
elagd	 ->2	a->3	
elakt	i->24	
eland	 ->5	,->2	e->44	s->6	
elar 	-->2	a->17	d->7	e->3	f->4	h->4	i->4	j->2	k->2	m->3	n->2	o->5	p->1	s->4	u->1	v->2	ä->1	
elar,	 ->3	
elar.	B->1	D->4	I->1	J->1	
elar:	 ->1	
elare	 ->5	.->1	n->4	
elarn	a->12	
elas 	a->2	d->1	i->3	k->1	
elas,	 ->2	
elas.	T->1	
elasp	e->1	
elast	a->6	n->4	
elat 	B->1	a->5	e->3	f->1	g->2	h->3	i->2	u->2	
elat,	 ->1	
elat.	H->1	
elate	r->4	
elati	o->9	v->13	
elats	 ->7	.->1	
elaye	d->2	
elbar	 ->1	a->5	t->14	
elber	ä->1	
elbro	t->1	
elbun	d->15	
elbyr	å->1	
eleda	n->2	
elefa	n->1	
elefo	n->1	
elega	t->17	
elege	r->4	
eleko	m->3	
elekt	i->1	r->10	
eleme	n->9	
elen 	a->15	f->1	g->1	i->3	k->1	m->1	o->1	v->1	ä->1	
elen"	 ->1	
elen,	 ->8	
elen.	D->3	
elenF	r->2	
elenä	t->1	
eler 	i->1	
eler.	D->1	
elern	a->5	
elers	u->3	
eles 	a->1	f->7	k->1	n->4	r->5	s->3	t->1	u->1	
elet 	o->1	
eleva	n->9	
eleve	r->1	
elevi	s->1	
elfed	e->1	
elfrå	g->3	
elfte	 ->1	
elfun	k->1	
elgad	o->1	
elgen	 ->1	
elgie	n->9	
elgis	k->8	
elgiv	n->1	
elhav	e->1	s->2	
elhet	 ->10	,->5	.->1	?->1	e->1	s->3	
elhjä	r->8	
elhoe	k->1	
elig 	f->1	
elig?	H->1	
eliga	 ->2	
elige	n->1	
eligg	a->8	e->18	
eligh	e->2	
eligi	ö->4	
eligt	 ->4	,->1	
elike	n->1	
elill	i->1	
elimi	n->6	
elinj	e->1	
elisk	 ->1	a->12	e->1	t->1	
elkri	t->1	
elkur	s->1	
elkvo	t->1	
ell b	a->1	e->2	l->2	
ell d	e->3	i->1	u->1	
ell e	l->1	n->1	u->1	
ell f	e->1	o->1	r->2	ö->7	
ell g	e->2	
ell i	 ->1	n->1	
ell k	o->5	ä->1	
ell l	i->1	ä->1	
ell m	e->2	å->2	
ell n	a->3	i->7	
ell o	c->6	e->1	l->1	m->1	r->1	
ell p	l->1	o->4	r->1	
ell r	e->4	i->1	ä->7	
ell s	a->1	o->6	t->1	u->1	
ell t	e->1	i->1	r->1	v->1	
ell u	n->1	p->1	
ell v	e->3	
ell å	k->1	t->1	
ell ö	k->1	p->2	
ell",	 ->1	
ell".	I->1	
ell, 	e->1	m->1	s->1	u->1	
ell- 	o->3	
ell.A	n->1	
ell.D	e->3	
ell.F	i->1	
ell.J	a->1	
ell.M	e->1	
ell.S	å->1	
ell.V	o->1	
ell.Ä	n->1	
ella 	E->1	F->1	a->11	b->22	d->15	e->6	f->32	g->5	h->8	i->13	j->5	k->16	l->5	m->25	n->7	o->30	p->27	r->32	s->35	t->9	u->13	v->4	ä->1	å->8	ö->1	
ella,	 ->3	
ella.	D->1	
ellam	t->1	
ellan	 ->192	"->1	,->3	.->2	l->1	n->1	s->7	t->1	ö->19	
ellbe	s->1	
ellbi	l->1	
ellek	t->3	
ellen	 ->2	,->1	
eller	 ->375	.->1	t->67	
ellfö	r->3	
elli 	h->1	
ellig	e->5	
ellis	e->2	
ellit	 ->1	
elliv	e->1	
ellmy	n->1	
ellre	 ->6	
ellrä	t->4	
ellsk	t->1	
ellt 	a->9	b->4	d->2	e->2	f->12	g->3	h->1	i->8	k->2	l->1	m->6	n->1	o->7	p->4	r->2	s->30	t->2	u->2	v->4	y->1	ä->2	å->1	ö->2	
ellt,	 ->6	
ellt.	D->1	
ellt;	 ->1	
ellån	g->4	
ellös	a->1	n->1	
elmaj	o->1	
elmas	t->1	
elmed	e->1	
elmsh	a->1	
elmäs	s->2	
eln "	u->1	
eln f	ö->3	
eln i	 ->1	
eln k	o->1	
eln m	e->1	
eln o	c->1	m->1	
eln t	i->5	
eln ä	r->2	
eln, 	d->1	h->1	
eln.D	e->1	
elnin	g->42	
elns 	l->2	
elodl	a->1	
eloge	 ->1	,->1	
elona	p->2	
elopp	 ->4	.->1	e->11	
elors	 ->2	.->1	
elpla	n->1	
elpro	b->1	
elpun	k->2	
elrap	p->1	
elreg	l->4	
elrik	t->1	
elrol	l->1	
elrum	 ->1	
elryc	k->1	
elräk	n->1	
elrät	t->2	
els a	l->1	t->3	v->3	
els d	ä->1	
els e	x->1	
els f	ö->2	
els i	n->1	
els k	o->1	
els o	c->1	
els p	r->2	
els s	k->1	t->1	
els t	i->2	
els v	a->1	ä->1	
els å	t->2	
els- 	o->1	
elsat	t->1	
elsdr	ä->1	
else 	-->3	a->14	b->1	d->2	e->1	f->16	g->2	h->3	i->5	j->3	k->5	m->15	n->4	o->17	p->2	r->1	s->20	t->2	u->1	v->1	ä->3	ö->4	
else,	 ->12	
else-	 ->1	
else.	B->1	D->5	E->2	J->3	K->1	L->1	M->2	N->1	S->2	V->2	
elsea	k->1	
elseb	y->1	
elsef	u->11	
elseh	i->1	
elsek	o->2	
elsel	ö->3	
elsem	ö->1	
elsen	 ->41	,->3	.->5	s->4	
elseo	m->1	
elser	 ->84	!->1	,->19	.->13	:->1	i->1	n->52	s->1	
elseu	t->1	
elsev	i->2	
elsex	p->1	
elsfl	o->2	
elsfr	å->2	
elsha	n->1	
elshi	n->1	
elsik	e->1	
elsin	d->2	g->20	
elsk-	f->1	
elska	 ->6	:->1	
elski	f->1	
elsko	n->2	
elskr	i->2	o->2	
elskt	 ->1	
elskv	a->1	
elsky	d->1	
elsla	g->5	
elslo	g->1	
elsmy	n->9	
elsmä	n->1	s->2	
elsny	h->1	
elsom	r->2	
elson	 ->4	.->1	
elsor	g->3	
elspl	a->2	
elspo	l->2	
elspr	o->2	
elsse	k->1	
elssj	ö->1	
elsst	ö->1	
elssä	k->43	
elst 	a->2	b->1	f->1	h->1	i->6	k->1	l->1	m->3	n->1	p->2	r->1	s->7	t->2	u->1	v->4	ä->1	
elst,	 ->7	
elst.	 ->1	A->1	F->1	V->1	
elsta	t->4	
elsti	l->1	
elsto	r->41	
elsut	a->3	
elsva	r->1	
elsyn	.->1	
elsys	t->2	
elsät	t->102	
elt -	 ->1	
elt E	U->1	
elt a	b->1	d->1	n->2	t->7	v->1	
elt b	e->1	
elt d	e->1	i->1	ä->1	
elt e	l->1	n->22	r->1	t->3	
elt f	l->1	r->2	ö->9	
elt g	o->3	
elt h	a->2	
elt i	 ->6	n->4	
elt k	l->16	o->8	
elt l	i->1	o->1	
elt m	e->3	o->1	
elt n	o->2	y->3	å->1	ö->1	
elt o	a->3	c->16	l->1	m->3	r->2	s->1	t->1	v->1	
elt p	a->1	å->2	
elt r	a->1	i->4	ä->6	
elt s	a->1	j->1	k->1	n->1	o->2	t->1	ä->8	
elt t	i->4	y->1	
elt u	p->2	t->2	
elt v	a->1	i->2	
elt ä	r->1	
elt å	t->1	v->1	
elt ö	v->3	
elt, 	o->1	
elt. 	D->1	
elt.D	e->3	
elt.E	n->1	
elt.H	e->1	ä->1	
elt.I	 ->1	
elt.J	a->1	
elt.U	n->1	
elt.V	a->2	
elt; 	d->1	
elt?J	a->1	
elta 	f->1	i->12	p->2	
elta,	 ->2	
eltag	a->24	i->6	
eltar	 ->9	
eltid	a->1	s->1	
eltis	k->1	
eltog	 ->2	
eltra	f->1	
eltäc	k->4	
elutb	e->2	
elux,	 ->1	
elva 	a->1	å->2	
elver	k->21	
elvis	 ->38	,->2	
elväg	g->3	
elvän	n->1	
elysa	 ->1	
elyse	r->1	
elysn	i->1	
elyst	 ->1	
elzen	.->1	
eläge	n->15	t->5	
elägg	a->2	e->1	n->1	s->1	
elägn	a->6	
elämn	a->3	
eländ	e->1	
elätt	n->1	
elöna	r->1	s->1	
elös 	-->1	
elösa	.->1	
elöst	 ->2	
em - 	a->1	s->1	
em 20	 ->1	
em al	l->2	
em an	d->1	
em at	t->5	
em av	 ->6	
em be	t->3	
em da	g->1	
em de	 ->2	l->1	n->1	r->1	t->1	
em di	k->1	
em dä	r->4	
em då	 ->1	l->1	
em ef	t->4	
em en	 ->4	l->1	
em et	t->2	
em fa	t->1	
em fr	å->3	
em fu	n->1	
em fö	r->29	
em gr	u->2	
em gå	n->1	
em gö	r->1	
em ha	r->4	
em he	l->1	
em hä	r->1	
em i 	E->1	T->1	b->2	d->6	f->5	h->1	n->1	o->1	s->1	u->1	v->1	Ö->1	
em in	f->1	o->4	t->2	
em ja	g->1	
em ka	n->2	
em ko	m->5	
em kr	ä->1	
em lä	m->1	n->1	
em me	d->20	n->1	r->2	
em mo	t->1	
em my	c->1	
em må	n->1	s->1	
em mö	j->1	
em ni	 ->1	
em nä	r->3	
em nå	g->1	
em oc	h->22	k->1	
em om	 ->3	
em pu	n->2	
em på	 ->11	
em re	l->1	
em se	g->1	
em sk	a->5	
em so	m->101	
em st	ö->1	
em så	 ->1	
em ti	l->6	
em ur	 ->1	
em ut	 ->1	a->1	v->2	
em va	r->2	
em ve	r->1	t->1	
em vi	 ->2	k->1	l->1	
em är	 ->8	
em år	 ->8	,->1	.->2	e->2	s->1	
em åt	g->1	
em öv	e->2	
em, a	n->1	
em, b	å->1	
em, d	ä->1	
em, e	f->2	x->1	
em, f	ö->2	
em, g	e->1	
em, h	a->1	u->1	
em, i	n->1	
em, k	a->1	
em, m	e->5	
em, o	c->4	
em, p	å->2	
em, s	e->1	o->1	å->1	
em, u	t->1	
em, v	a->2	i->3	
em, ä	n->1	
em, å	t->1	
em. D	e->1	
em. H	o->1	
em. M	a->1	
em.(A	p->1	
em.. 	F->1	
em.Al	l->1	
em.Av	b->1	
em.Be	t->1	
em.Bu	d->1	
em.De	 ->4	n->1	t->7	
em.Dä	r->3	
em.En	 ->1	
em.Eu	r->1	
em.Fr	u->1	
em.Fö	r->2	
em.Ge	n->1	
em.He	r->5	
em.In	o->1	
em.Ja	g->7	
em.Ko	m->1	
em.Ma	n->1	
em.Me	d->1	n->2	
em.Må	n->1	
em.Ne	j->1	
em.Ni	 ->1	
em.Nå	g->1	
em.Om	 ->1	
em.Pr	o->1	
em.Re	s->1	
em.Sl	u->1	
em.So	m->1	
em.Ty	v->1	
em.Ur	 ->1	
em.Ve	m->1	
em.Vi	 ->6	d->2	
em: A	s->1	
em: d	e->2	u->1	
em: p	a->1	
em; d	e->2	
em?De	t->1	
em?Me	n->1	
ema f	ö->1	
ema g	å->1	
ema h	ö->1	
ema, 	f->1	
emago	g->4	
emala	 ->1	
eman 	h->1	s->1	v->1	
eman.	H->1	
emang	 ->10	,->1	.->4	e->2	
emann	a->1	i->2	
emark	 ->1	
emask	e->1	
emat 	s->1	
emati	k->4	s->12	
embar	g->1	
ember	 ->30	,->8	.->6	v->1	
emble	m->1	
embry	o->1	
embur	g->6	
embyg	d->1	
emeda	n->1	
emede	l->1	
emell	a->7	e->59	i->1	
emen 	-->1	b->1	e->1	f->3	i->6	m->5	o->1	p->2	r->1	s->1	t->1	v->1	ä->1	
emen,	 ->4	
emen.	U->1	
emeni	n->5	
emens	a->196	k->194	
ement	 ->13	,->2	.->1	a->4	e->10	ä->2	
emest	e->4	
emet 	-->3	a->2	b->3	f->15	g->2	h->2	i->9	l->2	m->24	n->1	p->4	s->3	t->3	v->2	ä->15	
emet)	.->1	
emet,	 ->9	
emet.	B->1	D->1	E->1	H->2	I->2	J->2	M->2	N->1	P->1	V->2	
emet?	K->1	
emets	 ->1	
emför	d->1	
emhög	e->14	
emi, 	v->1	
emigr	a->1	e->1	
emik 	o->1	
emika	l->5	
emina	r->1	
emini	m->1	s->3	
emins	k->1	
emis-	f->1	
emisk	 ->1	.->1	
emism	 ->3	e->2	
emiss	 ->1	
emist	e->2	i->4	
emiti	s->3	
emiär	m->10	
emlan	d->3	
emlig	a->2	h->4	
emlän	d->1	
emläs	t->1	
emläx	o->1	
emlös	a->2	h->3	
emma 	h->1	i->4	o->1	s->1	ä->2	
emma,	 ->1	
emma:	 ->1	
emmap	l->1	
emmar	 ->7	!->1	,->5	.->1	
emmet	 ->1	
emogr	a->3	
emokr	a->137	
emomr	å->3	
emons	t->6	
emont	e->8	
emot 	-->2	E->1	I->1	J->1	T->2	U->1	a->8	b->3	d->20	e->8	f->3	h->4	i->5	k->2	l->1	m->4	n->3	o->1	p->2	s->9	t->2	v->7	y->1	Ö->1	ä->2	ö->2	
emot.	 ->1	F->2	V->1	
emoti	o->1	
empel	 ->71	,->5	.->3	:->3	v->28	
emper	a->4	
empla	r->2	
emple	n->3	t->3	
empor	ä->2	
empun	k->1	
ems a	n->2	
ems t	u->1	
ems- 	o->1	
emsan	 ->1	.->1	
emsk 	k->1	
emska	 ->3	p->2	s->1	
emsla	n->9	
emslä	n->27	
emsre	g->1	
emsst	a->284	
emt h	å->2	
emt r	a->1	
emt s	t->1	
emte 	F->1	b->1	d->1	h->1	k->1	p->2	r->6	v->1	
emted	e->2	
emtie	l->1	
emtio	 ->1	e->1	
emton	 ->5	
emvis	t->1	
emynd	i->1	
emän 	g->1	h->1	i->2	l->1	o->4	s->4	t->2	u->2	
emän,	 ->1	
emän.	I->1	
emänd	r->3	
emänn	e->12	
emäns	 ->3	
emärk	e->5	
emäss	i->1	
emål 	f->13	o->1	s->2	
emåna	d->1	
emåri	g->1	
emårs	p->2	
emöda	 ->3	
emöjl	i->4	
emöns	t->1	
emöta	 ->4	
emöte	r->1	
emöts	 ->2	
en "E	u->1	
en "L	o->1	
en "T	i->2	
en "d	e->1	ö->1	
en "e	u->2	
en "h	e->1	
en "n	o->1	
en "r	e->2	
en "s	p->1	
en "å	t->1	
en (1	4->2	9->1	
en (B	5->2	
en (E	I->1	
en (F	U->1	
en (I	M->1	
en (K	O->1	
en (e	l->1	
en (i	n->1	
en (m	a->1	
en (o	c->1	
en (s	å->1	
en , 	b->1	
en - 	"->1	2->1	6->1	A->1	R->1	a->3	b->2	d->7	e->5	f->2	h->5	i->3	j->2	l->2	m->1	o->6	s->4	u->2	v->3	ä->1	
en 1 	j->6	m->2	o->2	s->1	
en 1,	 ->1	
en 10	 ->1	
en 11	 ->2	
en 12	6->1	
en 13	 ->3	,->1	
en 14	 ->7	
en 15	 ->1	
en 16	 ->1	
en 17	 ->2	,->1	
en 18	 ->5	
en 19	 ->1	1->1	9->11	
en 2 	d->1	o->1	
en 2,	 ->1	
en 20	0->16	
en 21	 ->1	
en 23	 ->1	
en 24	 ->1	
en 26	 ->2	
en 29	,->1	
en 3 	f->1	j->1	m->1	o->1	
en 3,	 ->1	
en 30	 ->1	
en 31	 ->3	
en 38	 ->1	
en 39	,->1	
en 4 	j->2	
en 4,	 ->2	
en 5 	o->1	
en 6 	d->1	
en 7 	d->1	o->1	
en 79	/->1	
en 9 	d->1	f->1	
en 90	 ->1	
en AB	B->1	C->1	
en AD	R->1	
en Am	s->1	
en An	n->1	
en Ar	i->1	
en Ba	r->2	
en Be	l->1	r->3	
en Br	u->1	
en CE	N->1	
en Ca	s->1	
en Ch	a->1	
en De	 ->4	
en Du	i->1	
en EU	 ->1	-->1	:->2	
en En	 ->1	l->2	
en Er	i->1	
en Eu	r->11	
en FE	O->1	
en FN	,->1	
en Fö	r->1	
en Ga	r->1	
en Gr	a->1	e->1	u->1	
en Ha	i->1	
en I 	-->1	
en IM	O->1	
en IX	,->1	
en Is	a->1	r->1	
en Ja	c->2	
en Jo	r->1	
en Ju	g->1	
en Ka	l->2	r->3	
en Ki	n->4	
en Ko	c->2	m->1	
en La	n->1	
en Le	a->1	
en Lo	y->1	
en Mi	n->1	
en Na	t->2	
en PR	-->1	
en Pa	l->1	
en Pr	o->4	
en Ra	n->2	
en Re	d->2	
en Ro	v->1	
en SS	 ->1	
en Sc	h->1	
en So	l->1	
en Sy	r->1	
en Sã	o->1	
en Th	e->1	
en To	t->1	
en Ty	s->3	
en Un	i->2	
en Vi	v->1	
en Wo	g->1	
en XX	V->1	
en ab	s->2	
en ac	c->4	
en ad	e->1	m->5	r->1	v->1	
en ag	e->1	r->1	
en ak	t->10	
en al	b->2	d->2	l->44	
en am	b->1	e->3	
en an	 ->1	a->9	b->1	d->57	g->9	i->3	l->21	m->5	n->28	o->2	p->1	s->31	t->6	v->5	
en ar	a->1	b->13	t->5	
en as	p->6	y->1	
en at	t->270	
en au	k->2	t->1	
en av	 ->412	.->2	b->7	f->3	g->13	i->2	l->3	s->35	t->1	v->4	
en ax	e->1	
en ba	k->2	l->8	n->3	r->10	
en be	a->2	d->9	f->9	g->21	h->18	k->10	l->7	m->6	r->15	s->25	t->29	v->2	
en bi	b->1	d->3	l->12	n->1	o->2	t->1	
en bl	a->5	e->1	i->16	o->3	
en bo	k->3	r->12	s->1	t->3	
en br	a->14	e->7	i->14	o->4	u->1	ä->1	
en bu	d->9	
en by	g->2	r->6	
en bä	r->2	s->6	t->15	
en bå	d->3	
en bö	r->28	
en ce	n->8	r->1	
en ch	a->4	e->2	o->1	
en co	n->1	r->1	s->4	
en da	g->14	m->1	n->7	
en de	 ->24	a->1	b->21	c->3	f->5	g->1	l->55	m->15	n->29	r->1	s->2	t->126	
en di	a->7	k->1	r->3	s->12	v->1	
en dj	u->5	ä->1	
en do	c->1	g->1	k->2	m->6	
en dr	a->2	i->1	o->1	u->2	y->1	
en du	b->1	m->1	n->1	
en dy	n->1	
en dä	r->34	
en då	 ->7	v->1	
en dö	d->2	l->1	m->2	p->1	r->3	
en ef	f->19	t->23	
en eg	e->12	n->4	
en ej	 ->1	
en ek	o->49	
en el	e->2	l->28	o->2	
en en	 ->39	a->12	b->2	d->25	e->1	g->7	h->16	k->3	l->7	o->9	s->10	t->1	
en ep	o->1	
en er	b->2	h->1	i->1	k->3	t->1	
en et	n->3	t->18	
en eu	r->142	
en ev	e->4	
en ex	a->2	i->2	k->1	p->10	t->4	
en fa	k->5	l->3	n->1	r->4	s->7	t->4	
en fe	d->1	l->3	m->4	
en fi	c->2	l->1	n->24	
en fj	o->1	ä->6	
en fl	a->2	e->3	i->1	y->1	
en fo	k->1	l->2	n->4	r->18	
en fr	a->38	e->7	i->12	u->3	y->1	ä->2	å->115	
en fu	l->10	n->9	s->1	
en fy	s->2	
en fä	l->1	r->1	s->2	
en få	 ->5	n->1	r->19	t->1	
en fö	l->6	r->570	
en ga	m->7	n->6	r->12	v->1	
en ge	 ->2	d->1	m->95	n->35	o->1	r->4	s->1	
en gi	c->2	g->2	v->2	
en gj	o->11	
en gl	a->1	e->1	o->3	ä->6	
en gn	u->2	
en go	d->24	
en gr	a->13	e->5	u->25	ä->2	ö->1	
en gu	m->1	
en gy	n->1	
en gä	l->21	r->1	
en gå	 ->1	n->49	r->5	
en gö	r->14	
en ha	 ->5	d->7	f->4	l->8	m->3	n->22	r->201	
en he	b->1	j->1	l->26	m->2	r->1	
en hi	s->3	t->2	
en hj	ä->5	
en ho	n->1	p->7	r->1	s->8	t->6	
en hu	n->1	r->4	v->6	
en hy	p->1	s->1	
en hä	m->2	n->12	r->69	v->2	
en hå	l->15	r->4	
en hö	g->22	j->2	r->3	
en i 	A->5	B->7	C->1	D->2	E->22	F->4	G->4	H->2	I->4	K->9	L->6	M->7	N->2	O->1	R->2	S->11	T->9	V->1	W->2	a->11	b->5	c->2	d->68	e->19	f->42	g->6	h->7	i->3	k->8	l->4	m->21	n->1	o->6	p->9	r->10	s->42	t->2	u->16	v->18	z->1	Ö->14	å->1	ö->1	
en ic	k->4	
en id	e->3	é->3	
en if	r->1	
en ih	ä->1	å->1	
en il	l->3	
en im	p->1	
en in	 ->1	b->2	c->1	d->6	e->2	f->20	g->5	h->2	l->5	n->19	o->37	r->68	s->20	t->131	v->3	
en ir	a->1	l->2	
en is	r->10	
en it	a->4	
en ja	g->87	k->2	
en ju	 ->1	b->1	r->5	s->9	
en jä	m->6	
en ka	l->2	m->4	n->87	r->1	s->2	t->12	
en ke	d->1	l->1	
en ki	n->1	
en kl	a->17	
en kn	a->1	
en ko	a->4	l->2	m->152	n->59	p->3	r->4	s->10	
en kr	a->11	i->11	ä->13	
en ku	l->10	n->13	r->1	
en kv	a->3	o->4	
en kä	l->3	n->15	r->1	
en la	d->2	g->11	r->1	
en le	d->7	g->2	
en li	b->3	g->7	k->6	n->3	t->10	v->1	
en lo	g->1	k->5	v->2	
en lu	c->1	
en ly	c->2	d->1	s->1	
en lä	g->12	m->4	n->3	r->1	t->2	
en lå	g->3	n->19	t->2	
en lö	j->1	k->1	s->15	
en ma	g->1	j->3	k->2	l->1	n->11	r->13	s->5	x->2	
en me	d->143	l->33	n->14	r->21	s->2	t->5	
en mi	l->12	n->31	s->12	t->1	
en mo	d->13	n->3	t->36	
en mu	l->1	n->3	
en my	c->64	n->8	
en mä	n->14	r->3	t->1	
en må	 ->1	h->1	l->1	n->10	s->94	
en mö	j->17	r->2	t->3	
en na	t->19	
en ne	d->7	g->4	u->1	
en ni	 ->4	o->1	v->2	
en no	g->1	l->1	m->1	r->5	t->3	
en nu	 ->14	,->1	m->1	v->14	
en ny	 ->24	a->38	c->2	e->1	l->3	s->2	t->4	
en nä	m->7	r->34	s->1	
en nå	b->2	g->16	
en nö	d->14	j->1	t->1	
en oa	c->2	n->2	v->2	
en ob	a->1	e->19	l->5	
en oc	h->399	k->43	
en oe	g->1	n->1	r->2	
en of	a->1	f->23	t->1	ö->5	
en oh	ä->1	
en ok	l->2	o->1	ä->2	
en ol	j->1	y->6	
en om	 ->230	,->2	.->1	I->1	b->1	e->4	f->13	i->1	m->1	o->1	p->2	r->5	s->3	v->6	ö->1	
en on	d->1	e->1	ö->2	
en op	e->1	t->2	
en or	d->10	g->5	i->1	k->1	m->1	o->22	t->1	ä->1	
en os	s->2	
en ot	a->1	i->2	j->1	
en ou	m->2	n->1	
en ov	a->1	i->1	
en oä	n->1	
en oö	n->1	v->2	
en pa	l->4	r->14	s->2	
en pe	k->2	r->20	t->1	
en pl	a->15	u->1	ö->1	
en po	e->1	l->50	r->5	s->15	
en pr	a->1	e->8	i->10	o->23	
en pu	n->27	r->1	
en py	r->1	
en på	 ->147	?->1	f->1	g->5	m->1	p->2	s->1	t->1	v->3	
en ra	d->20	m->1	p->7	s->3	t->1	
en re	a->1	d->17	e->2	f->17	g->46	k->3	l->4	n->8	s->27	v->7	
en ri	k->15	m->3	s->10	
en ro	l->4	
en ru	n->2	
en ry	s->1	
en rä	c->2	d->3	k->5	t->38	
en rå	d->8	g->1	
en ré	f->1	
en rö	d->2	r->2	s->7	
en sa	d->5	k->16	m->33	n->3	t->6	
en sc	e->1	o->1	
en se	 ->5	d->5	g->2	k->2	n->12	p->1	r->12	t->1	x->1	
en si	f->1	g->3	n->4	s->16	t->13	
en sj	u->5	ä->26	
en sk	a->127	e->3	i->7	j->2	o->2	r->7	u->46	y->9	ä->2	ö->2	
en sl	a->4	o->1	u->15	
en sm	i->1	u->1	ä->2	å->1	
en sn	a->12	e->2	
en so	c->39	l->2	m->233	r->5	
en sp	a->3	e->11	l->1	r->3	ä->1	
en sr	i->1	
en st	a->43	i->4	o->52	r->34	u->7	y->2	ä->13	å->19	ö->36	
en su	b->2	c->1	m->1	n->2	p->1	
en sv	a->4	e->1	å->2	
en sy	f->3	m->3	n->6	r->2	s->3	
en sä	g->7	k->4	l->2	r->10	t->2	
en så	 ->27	,->1	d->41	g->1	s->2	v->1	
en sö	d->1	k->1	
en ta	 ->4	c->8	g->1	l->6	n->2	r->6	
en te	c->1	k->8	r->4	x->2	
en ti	b->3	d->37	l->166	m->1	t->3	
en tj	ä->5	
en to	g->2	l->2	m->1	n->2	t->11	
en tr	a->5	e->15	o->10	ä->2	ö->1	
en tu	f->1	n->4	r->3	
en tv	e->6	i->5	ä->2	å->3	
en ty	c->3	d->14	g->1	n->2	p->5	s->12	v->4	
en tä	n->4	
en un	d->54	g->1	i->9	
en up	p->50	
en ur	 ->3	s->5	v->1	
en ut	a->14	b->2	e->2	f->4	g->10	i->1	j->1	l->1	m->7	n->2	p->1	s->10	t->6	v->27	ö->2	
en va	d->6	l->7	n->4	r->42	t->1	
en ve	c->2	d->2	m->2	r->27	t->10	
en vi	 ->72	d->39	k->50	l->36	n->1	s->39	t->3	
en vo	l->1	r->2	
en vä	c->1	d->2	g->2	l->10	n->7	r->8	s->4	v->1	x->6	
en vå	l->3	
en wa	l->1	
en yt	t->5	
en zi	g->2	
en Ös	t->1	
en äg	a->1	n->1	
en äl	s->1	
en än	 ->6	d->27	n->9	t->1	
en är	 ->207	,->1	.->2	a->1	l->1	
en äv	e->16	
en å 	a->1	d->3	e->2	
en åb	e->1	
en åk	l->2	
en ål	a->1	d->2	
en år	 ->2	
en ås	i->9	t->1	y->1	
en åt	 ->7	a->1	e->13	f->2	g->9	s->1	t->1	
en öd	e->1	
en ök	a->21	n->9	
en öm	 ->1	
en ön	s->4	
en öp	p->6	
en ör	e->1	
en ös	t->18	
en öv	e->53	n->2	
en! E	r->1	
en! J	a->1	
en! M	i->1	
en! N	i->1	
en!Nä	r->2	
en!Rö	s->1	
en" a	l->1	
en" e	t->1	
en" i	 ->1	
en" o	c->1	
en" s	o->1	
en", 	"->1	o->1	s->1	
en".D	e->3	
en".O	r->1	
en) (	S->1	
en) f	ö->1	
en) h	a->1	
en) z	o->1	
en)(P	a->2	
en), 	o->1	
en).D	e->1	
en).H	e->1	
en)Ja	g->1	
en)Nä	s->1	
en, "	o->1	
en, 1	 ->1	0->1	5->1	9->1	
en, 8	,->1	
en, A	m->2	
en, B	N->1	e->3	
en, C	u->1	
en, E	u->2	
en, I	V->1	r->1	
en, J	o->1	
en, K	a->1	o->1	
en, L	o->1	
en, N	e->1	
en, P	a->2	e->1	
en, R	a->1	
en, S	l->1	v->1	
en, T	o->1	y->1	
en, V	 ->1	l->1	
en, W	i->1	
en, a	l->4	n->2	t->10	v->2	
en, b	a->2	l->5	o->1	r->1	å->3	ö->5	
en, d	e->31	v->5	ä->11	å->2	
en, e	f->12	k->1	l->3	n->10	t->6	x->1	
en, f	a->1	i->2	r->18	å->2	ö->42	
en, g	e->3	r->1	
en, h	a->8	e->15	ä->1	ö->1	
en, i	 ->15	n->20	
en, j	a->3	u->4	
en, k	a->5	o->8	u->1	v->1	ä->3	
en, l	i->5	ä->2	å->1	
en, m	a->1	e->36	i->3	ä->1	å->7	
en, n	a->1	ä->14	å->5	
en, o	c->84	m->10	s->1	
en, p	a->3	r->1	å->6	
en, r	ä->1	å->3	
en, s	a->6	e->1	k->9	l->2	n->2	o->58	t->3	ä->6	å->18	
en, t	.->2	a->3	i->11	r->3	v->3	y->4	
en, u	n->1	p->1	t->21	
en, v	a->8	i->31	o->1	ä->1	
en, y	t->1	
en, Î	l->1	
en, ä	g->1	n->1	r->13	v->12	
en, å	t->1	
en, ö	p->1	
en-SS	:->1	
en. D	e->4	ä->1	
en. F	o->1	
en. H	a->1	ä->1	
en. I	n->1	
en. J	a->3	
en. L	å->1	
en. M	e->2	
en. N	ä->1	
en. O	c->2	
en. V	i->2	
en." 	Ä->1	
en.(E	L->1	
en.(I	T->1	
en.).	H->1	
en.)A	n->1	
en.)B	e->4	
en.)F	r->3	
en.)G	e->1	
en.)H	e->1	
en.. 	(->9	
en..(	E->2	N->1	
en..H	e->1	
en.15	 ->1	
en.Al	l->9	
en.An	d->1	n->1	
en.Ar	b->1	t->1	
en.At	t->3	
en.Av	 ->6	
en.Be	t->2	
en.Bi	l->1	
en.Br	y->1	
en.Cu	n->1	
en.De	 ->15	n->37	s->10	t->138	
en.Dä	r->20	
en.Då	 ->1	
en.EU	 ->2	
en.Ef	f->1	t->2	
en.Em	e->1	
en.En	 ->7	d->2	l->4	
en.Er	 ->1	i->1	
en.Et	t->9	
en.Eu	r->5	
en.FE	O->1	
en.Fa	k->1	r->1	
en.Fi	n->1	
en.Fo	r->1	
en.Fr	u->3	å->3	
en.Fy	r->1	
en.Fö	l->1	r->32	
en.Ge	n->1	
en.Go	l->1	
en.Gå	 ->1	
en.Ha	d->1	n->4	r->2	
en.He	r->44	
en.Hi	t->2	
en.Ho	n->2	
en.Hu	r->2	
en.Hä	r->6	
en.I 	E->1	T->1	d->9	e->5	m->3	r->2	s->6	v->1	
en.In	g->1	o->1	r->1	s->1	
en.Ja	,->1	g->99	
en.Jo	r->1	
en.Ju	s->1	
en.Ka	n->5	
en.Ko	c->1	m->15	n->3	
en.Kr	a->1	
en.Ku	l->1	
en.Kv	a->1	
en.Le	d->1	
en.Li	k->1	
en.Lå	n->1	t->6	
en.Ma	n->5	r->1	x->1	
en.Me	d->5	n->28	
en.Mi	n->3	t->1	
en.Mo	t->4	
en.My	n->1	
en.Mä	n->1	r->1	
en.Må	n->1	
en.Na	t->2	
en.Ni	 ->6	
en.Nu	 ->4	
en.Ny	l->1	
en.Nä	r->7	
en.Oc	h->9	k->1	
en.Om	 ->12	
en.Or	d->4	s->1	
en.Oz	 ->1	
en.Pa	r->4	
en.Pe	r->1	
en.Pl	a->1	
en.Pr	e->1	o->2	
en.På	 ->9	
en.Re	f->1	n->1	
en.Ri	k->1	
en.Ro	t->1	
en.Rä	t->1	
en.Rå	d->4	
en.Sa	m->3	n->2	
en.Se	d->1	t->1	
en.Si	s->1	t->1	
en.Sk	a->1	
en.Sl	u->8	
en.Sn	a->1	
en.So	m->8	
en.St	a->1	ö->2	
en.Su	b->1	
en.Sy	f->2	
en.Sä	k->1	r->2	
en.Så	 ->4	
en.Ta	c->4	
en.Th	e->1	y->1	
en.Ti	d->1	l->4	
en.To	r->2	
en.Tr	o->2	
en.Tv	ä->1	
en.Ty	 ->1	v->2	
en.Un	d->5	i->1	
en.Up	p->1	
en.Ut	a->1	i->1	v->1	
en.Va	d->7	r->1	
en.Ve	t->1	
en.Vi	 ->69	d->3	l->2	s->1	t->1	
en.Vå	r->2	
en.Än	 ->1	d->1	
en.Är	a->2	
en.Äv	e->4	
en.Å 	E->1	a->1	
en.Ög	o->1	
en.Öv	e->1	
en: "	d->1	
en: D	e->1	
en: E	r->1	
en: H	a->1	
en: J	a->2	
en: K	o->2	
en: R	e->1	
en: T	å->1	
en: d	e->2	ä->1	
en: f	o->1	ö->2	
en: i	n->1	
en: j	a->1	
en: m	e->2	
en: v	a->3	i->1	
en:Fö	r->1	
en; a	v->1	
en; d	e->6	ä->1	
en; e	n->1	
en; f	i->1	ö->1	
en; i	n->1	
en; m	e->1	
en; o	c->1	
en; p	u->1	
en; s	a->1	
en; ä	n->1	
en?. 	(->1	
en?De	n->2	s->1	t->4	
en?Ef	t->1	
en?Fo	l->1	
en?Fr	u->1	
en?Fö	r->2	
en?He	r->2	
en?I 	d->1	
en?Ja	g->2	
en?Ka	n->1	
en?Ko	m->1	
en?Nä	r->1	
en?Va	d->1	
en?Ve	m->1	
en?Vi	 ->3	l->3	
en?Är	 ->3	
enFrå	g->3	
enHer	r->2	
enI d	e->1	
enJag	 ->2	
enNäs	t->5	
ena -	 ->1	
ena B	 ->1	
ena a	l->1	v->4	
ena d	e->3	
ena e	f->1	l->5	n->2	t->1	
ena f	a->2	r->3	u->1	å->1	ö->6	
ena g	a->1	ä->3	å->1	
ena h	a->1	
ena i	 ->15	n->1	
ena k	o->3	u->1	v->1	
ena l	a->1	ä->1	
ena m	e->5	i->1	o->1	
ena o	c->10	m->2	
ena p	a->1	å->2	
ena r	e->2	ö->1	
ena s	i->16	k->2	o->1	t->1	
ena t	a->1	
ena u	p->1	t->2	
ena v	o->1	å->1	
ena y	t->1	
ena ä	r->4	
ena ö	g->1	s->1	
ena, 	d->2	f->1	m->1	n->1	o->4	s->3	t->3	v->1	
ena. 	H->1	
ena.D	e->2	
ena.E	t->1	
ena.F	ö->1	
ena.J	a->3	u->1	
ena.O	m->1	
ena.V	a->1	i->1	
ena.Ä	v->1	
ena; 	p->1	
ena?P	å->1	
enad 	i->1	n->1	r->1	u->2	
enad,	 ->1	
enad?	H->1	
enade	 ->22	,->1	.->1	s->2	
enand	e->7	
enans	v->1	
enant	 ->1	
enar 	a->7	b->1	d->5	e->1	h->1	i->1	j->6	k->1	n->3	o->1	p->1	s->5	v->1	
enar,	 ->2	
enar.	D->1	V->1	
enar:	 ->1	
enare	 ->24	,->4	.->2	l->1	n->4	
enari	e->1	o->4	
enarn	a->5	
enars	a->4	
enarå	d->1	
enas 	h->1	i->1	m->4	n->1	o->2	t->1	
enast	 ->13	?->1	e->63	å->2	
enat.	 ->1	
enate	n->1	
enats	 ->1	
enaue	r->1	
enavt	a->3	
enbar	 ->1	.->2	a->1	l->12	t->50	
enber	g->3	
enbet	ä->5	
enbur	g->2	
encer	,->1	
end f	ö->1	
end i	 ->1	
end j	u->1	
end o	c->2	
end u	n->1	
end! 	L->1	N->1	
end, 	f->1	t->1	
end- 	(->1	
enda 	2->1	E->1	a->1	c->1	d->3	e->2	f->2	i->1	j->2	l->3	m->4	n->1	o->1	p->6	r->3	s->16	v->3	ö->1	
enda.	R->1	
endai	r->1	
endas	t->71	
endat	i->33	
endbe	t->1	
ende 	"->1	-->4	A->1	B->1	K->1	M->1	a->28	b->9	d->8	e->23	f->27	g->1	h->6	i->7	j->1	k->6	l->1	m->5	n->4	o->13	p->24	r->14	s->15	t->12	u->3	v->7	ä->3	å->2	ö->2	
ende"	,->1	
ende,	 ->11	
ende.	D->5	F->1	H->3	J->3	M->4	O->1	S->3	V->1	
ende:	 ->22	
ende;	 ->1	
endef	ö->2	
endek	r->1	
endel	a->1	
endem	i->1	
enden	 ->18	,->1	.->3	a->3	s->11	
ender	 ->4	a->19	k->1	u->2	ö->1	
endes	 ->1	k->1	
endet	 ->33	.->4	s->1	
endev	a->6	
endie	r->1	
endom	 ->2	l->2	s->1	
endra	g->1	
ends 	b->2	
endt 	f->1	h->1	o->1	s->1	t->1	u->1	
endt,	 ->1	
endée	,->1	
endöv	t->1	
enefi	t->5	
enelu	x->1	
enema	n->1	
enen 	f->2	
enen.	J->1	
ener 	(->2	I->4	i->1	
ener-	p->10	
enerN	ä->1	
enera	 ->1	d->1	l->20	r->1	t->4	
enere	l->16	r->3	
energ	i->109	
enerö	s->4	
enet 	a->1	p->1	
eneti	s->1	
enezu	e->1	
enfrå	g->1	
enfär	d->1	
enför	d->1	e->5	s->1	
enga 	k->1	
engag	e->18	
engar	 ->28	,->5	.->6	?->1	n->15	
engel	s->10	
engen	 ->2	,->1	a->3	k->1	o->1	r->1	s->1	
engue	r->2	
engäl	d->1	
engör	 ->1	i->2	
enham	n->1	
enhan	d->1	
enhet	 ->41	"->2	,->11	.->17	e->76	l->36	s->10	
enhäl	l->32	
enhår	d->1	
eni f	ö->1	
eni s	a->1	
eni.A	l->1	
enied	 ->1	.->1	
enig 	i->1	
eniga	 ->2	,->1	.->1	
enigh	e->9	
enind	u->1	
ening	 ->35	,->2	.->1	a->17	e->17	s->16	
enist	a->2	
enjör	 ->2	
enkel	 ->3	:->2	m->1	r->1	t->27	v->2	
enkla	 ->10	d->1	r->4	s->3	
enkli	n->1	
enkol	e->1	
enkon	v->1	
enkän	n->1	
enlig	 ->4	a->3	h->34	t->93	
enlös	 ->1	
enna 	-->1	E->1	a->17	b->25	c->2	d->33	e->9	f->94	g->21	h->6	i->14	j->1	k->51	l->9	m->25	n->2	o->10	p->37	r->65	s->58	t->27	u->18	v->24	y->1	ä->3	å->5	ö->8	
enna,	 ->2	
enna.	-->1	D->1	J->3	O->1	V->1	Ä->1	
enna?	S->1	
enndr	a->1	
enne 	F->1	a->2	f->2	h->3	t->1	ä->2	
enne.	J->1	
ennes	 ->21	,->1	
ennie	f->1	r->5	s->2	t->3	
ennin	g->10	
enniu	m->3	
enom 	A->1	D->1	E->5	S->1	W->1	a->109	b->5	d->23	e->20	f->5	g->1	h->3	i->6	k->3	l->2	m->5	n->2	o->2	p->5	r->1	s->7	t->4	u->5	v->5	y->1	ä->2	å->3	ö->2	
enom,	 ->1	
enom.	H->1	V->1	
enoma	r->2	
enomb	l->5	r->2	
enomd	r->6	
enome	n->3	
enomf	ö->161	
enomg	i->1	r->4	å->11	
enoml	ä->2	
enomr	å->1	
enoms	k->1	l->3	n->11	y->3	
enomt	ä->1	
enorm	 ->7	a->18	t->7	
enove	r->3	
enpro	b->1	
enreg	e->1	
enren	i->1	
enres	u->1	
enry 	F->1	
enröt	t->1	
ens 2	8->1	
ens B	N->3	
ens E	U->1	u->2	
ens I	s->1	
ens V	D->1	
ens X	X->1	
ens a	d->1	g->1	l->4	n->17	r->8	t->2	v->8	
ens b	a->1	e->28	i->1	l->2	r->1	u->7	y->1	ä->1	å->2	
ens c	e->1	
ens d	a->9	e->13	i->5	o->5	ä->1	
ens e	f->5	g->4	k->17	l->1	m->1	n->4	x->3	
ens f	a->5	e->2	i->3	o->5	r->12	u->2	ö->52	
ens g	a->1	e->5	o->2	r->8	å->1	
ens h	a->7	e->1	i->3	o->1	u->1	ä->4	
ens i	 ->5	d->1	k->1	m->1	n->40	
ens j	o->2	u->2	
ens k	a->2	o->23	r->4	u->4	v->3	ä->2	
ens l	a->9	e->2	i->3	j->1	o->2	ä->7	ö->1	
ens m	a->3	e->34	i->5	o->4	y->1	å->6	ö->3	
ens n	a->4	e->1	i->2	u->6	ä->1	å->1	ö->1	
ens o	b->2	c->20	d->1	i->2	l->1	m->31	r->14	t->2	
ens p	a->7	e->2	l->2	o->10	r->7	å->3	
ens r	a->13	e->34	i->4	o->8	u->1	ä->17	å->1	ö->1	
ens s	a->11	e->3	i->16	j->1	k->7	l->3	n->2	o->11	p->3	t->33	v->1	y->3	ä->7	
ens t	a->4	e->8	i->5	j->7	o->1	r->4	u->1	
ens u	n->1	p->7	r->5	t->35	
ens v	a->2	e->7	i->16	ä->11	
ens y	t->7	
ens ä	g->4	n->3	r->5	
ens å	l->2	r->3	s->2	t->3	
ens ö	d->3	k->1	r->1	v->8	
ens!V	i->1	
ens, 	b->1	d->3	f->3	m->3	n->1	o->7	p->1	s->2	v->1	
ens- 	o->2	
ens.D	e->6	
ens.F	ö->1	
ens.I	 ->1	
ens.J	a->2	
ens.M	a->1	
ens.O	a->1	
ens.S	o->1	
ens/d	e->1	
ens: 	h->1	
ens?E	t->1	
ens?J	a->1	
ensa 	u->2	
ensam	 ->48	,->1	m->131	r->1	t->26	
ensar	 ->1	
ensat	i->3	t->1	
ensav	g->1	
ensbe	g->3	r->1	s->6	v->2	
ensde	b->2	
ensdo	m->1	
ensdu	g->2	
ense 	m->4	o->1	v->1	
ense,	 ->1	
ensen	 ->102	,->13	.->36	?->1	N->1	s->17	
enser	 ->27	,->1	.->7	a->7	n->18	
ensfr	i->1	ä->1	å->3	
ensfö	r->3	
enshi	n->2	
enshä	m->2	
ensib	i->1	
ensid	i->4	
ensif	i->3	
ensin	 ->1	i->1	n->1	r->1	
ensio	n->26	
ensis	k->2	
ensit	e->1	
ensiv	 ->3	a->3	t->6	
ensk 	T->1	k->1	
enska	 ->15	p->298	
enske	 ->2	
enski	l->28	
ensko	m->18	
enskr	a->35	i->3	
enskt	 ->2	
ensku	l->5	
ensme	d->1	
ensmi	n->1	
ensmy	n->8	
ensmå	l->1	
ensna	c->2	
ensni	n->7	
ensom	r->2	
ensor	d->1	
enspo	l->76	
enspr	i->5	
ensra	m->1	
ensre	g->9	l->1	
ensrä	t->9	
enssi	t->1	
enssk	a->1	y->2	
ensst	ä->20	ö->1	
enssv	å->1	
enssy	s->1	
ensta	k->5	t->1	
enstr	e->2	
ensut	s->2	
ensva	r->1	
ensve	r->1	
ensvi	l->9	
ensvä	n->1	
ensär	e->2	
ent (	t->1	
ent -	 ->3	
ent 1	9->2	
ent A	s->1	
ent C	l->1	
ent a	l->5	n->2	t->2	v->50	
ent b	a->1	o->1	r->1	u->1	ö->1	
ent e	k->1	l->3	n->2	
ent f	r->3	y->1	ö->33	
ent g	e->4	r->1	
ent h	a->7	e->1	o->1	u->2	
ent i	 ->14	d->1	g->1	n->8	
ent k	a->4	o->5	r->1	u->1	v->1	
ent l	e->1	
ent m	e->7	o->2	å->1	
ent o	c->24	m->4	
ent p	å->4	
ent r	e->2	
ent s	a->1	e->2	j->1	k->3	o->28	t->1	ä->4	å->1	
ent t	a->1	e->2	i->12	
ent u	n->2	p->2	t->2	
ent v	a->2	e->1	ä->1	
ent ä	n->1	r->4	
ent å	t->1	
ent ö	n->1	v->2	
ent, 	L->1	S->1	a->1	b->1	d->2	e->2	f->2	g->1	i->4	k->1	m->2	o->4	r->2	s->2	u->1	v->1	
ent. 	V->1	
ent.D	e->8	
ent.E	n->1	u->1	
ent.F	r->1	ö->3	
ent.H	e->2	
ent.I	 ->4	
ent.J	a->5	
ent.L	å->1	
ent.M	a->1	e->2	
ent.N	ä->1	
ent.O	K->1	
ent.P	l->1	
ent.S	a->1	
ent.V	i->1	
enta 	N->1	S->1	a->1	b->1	f->1	h->1	i->1	m->1	n->10	p->1	r->1	s->17	
enta,	 ->1	
entab	l->1	
ental	 ->1	a->2	i->1	s->10	
entan	d->2	s->6	t->10	
entar	 ->2	,->1	e->21	i->27	
entat	 ->4	e->1	i->16	
entav	 ->1	
entek	n->1	
entem	o->27	
enten	 ->23	,->5	.->4	s->4	
enter	 ->15	,->1	.->4	a->45	i->3	n->34	
entet	 ->306	,->37	-->1	.->29	:->1	?->1	s->103	
entfr	å->6	
entia	l->3	
entie	l->6	r->5	
entif	i->11	
entil	 ->1	e->1	i->1	
entim	e->1	
entin	g->22	s->1	
entio	n->41	
entit	e->8	
entka	t->1	
entli	g->207	
entor	g->1	
entpo	l->2	
entra	 ->4	,->1	l->76	t->16	
entre	l->1	p->5	r->15	t->1	
entru	m->9	
ents 	a->1	b->1	h->1	i->1	m->1	t->1	
entsa	t->1	
entsb	e->1	
entsf	o->1	
entsi	f->1	
entsk	a->1	o->1	y->5	
entsl	e->28	
entsu	t->2	
entti	l->1	
entue	l->21	
entur	e->1	
entus	i->3	
entva	r->1	
entvä	n->1	
entyd	i->4	
entyr	a->9	
entär	a->2	
enum 	f->1	h->1	i->1	ä->1	
enum.	D->1	
enusd	i->1	
enutv	e->1	
envet	e->1	
envis	a->1	h->3	t->1	
enväg	a->8	
enz b	e->1	
enz e	t->1	
enz f	r->1	ö->1	
enz o	c->6	m->1	
enz t	o->1	
enz)(	T->1	
enz).	H->1	
enz, 	L->3	
enzFr	u->1	
enzbe	t->1	
enÄra	d->1	
enägn	a->1	
enämt	 ->1	
enät 	k->1	
enåda	 ->1	
enève	 ->1	,->1	k->1	
enör 	t->1	
enörs	k->2	
eogra	f->8	
eolog	,->1	i->4	
eområ	d->3	
eonaz	i->1	
eoni 	s->1	
eonla	m->1	
eordr	a->1	
eoret	i->2	
eostr	a->2	
eote 	Q->1	
ep at	t->1	
ep ma	n->1	
epa a	t->1	
epa d	e->6	
epa m	i->4	
epa n	å->2	
epa p	a->1	
epa v	å->1	
epa, 	o->1	
epade	 ->8	
epar 	-->1	a->2	d->5	h->1	j->1	m->2	o->1	r->1	s->1	
epara	b->1	t->2	
epare	r->4	
epart	e->9	
epas 	d->1	i->2	n->1	o->1	
epas.	J->1	V->1	
epat 	-->1	s->1	
epat:	 ->1	
epats	 ->2	
epesk	å->1	
epher	d->3	
epnin	g->1	
epok 	i->1	
epok,	 ->1	
epoke	n->2	
epoli	s->1	t->1	
eposi	t->1	
epoti	s->5	
epp a	l->1	
epp i	 ->4	n->1	
epp o	c->1	m->1	
epp p	å->3	
epp s	o->1	
epp, 	b->1	
eppa 	s->1	
eppen	 ->1	
eppet	 ->10	
eppsb	r->1	y->1	
eppsr	e->2	
eppss	ä->2	
eppsv	a->2	
epren	ö->3	
epres	e->19	s->2	
epris	e->2	
eprod	u->1	
eprog	r->1	
epsis	 ->1	
epskä	l->1	
ept i	 ->1	
ept k	o->1	
ept.D	e->1	
ept.H	a->1	
eptab	e->27	l->10	
eptan	s->7	
epte 	f->1	
eptem	b->15	
epter	a->45	
eptet	 ->3	
eptik	e->3	
eptio	n->6	
eptis	k->5	
epubl	i->19	
er (C	5->2	
er (a	r->1	
er (i	 ->1	
er - 	1->2	a->6	c->1	d->8	e->3	g->1	h->1	i->6	k->3	m->1	n->1	o->3	s->5	t->1	v->1	ä->5	
er 1 	4->1	
er 10	 ->1	
er 19	3->1	8->1	9->27	
er 2 	b->1	
er 20	 ->2	0->3	
er 27	 ->1	
er 32	 ->1	
er 35	 ->1	
er 4 	0->1	
er 40	 ->2	
er 5 	å->1	
er 50	 ->1	
er 60	 ->1	
er 7 	g->1	
er 73	,->1	
er 80	 ->3	
er 90	 ->2	
er 97	/->1	
er Al	s->1	t->1	
er Am	o->2	
er Ar	a->1	
er Az	o->1	
er BN	I->1	
er BS	E->1	
er Ba	r->2	
er Br	y->1	
er Co	c->1	n->1	
er Da	n->1	
er Du	h->1	
er EG	-->1	.->1	
er EM	U->2	
er EU	:->3	
er Eh	u->1	
er Ek	o->1	
er El	s->1	
er Er	i->2	
er Eu	r->23	
er Ex	x->1	
er FN	:->2	
er Fa	r->1	
er Fi	n->1	
er Fö	r->3	
er GA	S->1	
er Ga	m->2	
er Go	m->1	
er Gr	e->1	
er Gu	s->1	t->1	
er He	l->1	
er Hi	m->1	
er I 	o->1	
er I-	p->1	
er II	 ->1	-->2	I->1	
er Is	r->3	
er It	a->1	
er Ja	p->1	
er Jo	n->1	s->1	
er Jö	r->2	
er Ki	n->2	
er Kv	i->1	
er La	a->7	
er Li	s->1	
er Ly	n->1	
er Ma	a->2	
er Me	l->1	
er Na	t->1	
er Ne	d->1	
er Ni	k->2	
er OF	S->1	
er Or	a->1	
er Os	l->1	
er PV	C->1	
er Pa	l->1	
er Ra	s->1	
er Ru	s->1	
er Sc	h->3	
er Se	a->1	i->1	
er Sh	a->1	
er Sk	o->1	
er Sy	r->2	
er Ta	m->1	n->1	
er To	r->1	
er Tu	r->3	
er UN	M->1	
er US	A->1	D->1	
er Ur	q->1	
er Vi	t->1	
er [S	E->1	
er ab	s->1	
er ac	c->1	
er ak	t->3	
er al	d->3	l->46	
er am	e->1	
er an	a->2	b->1	d->17	f->2	h->1	l->1	m->1	n->4	o->1	s->12	t->3	v->5	
er ar	b->10	t->4	
er as	y->1	
er at	t->785	
er au	c->1	
er av	 ->74	b->2	d->1	f->1	g->2	s->8	t->1	v->1	
er ba	k->7	r->5	s->1	
er be	a->2	d->3	f->2	g->4	h->9	k->4	r->3	s->8	t->11	v->5	
er bi	d->5	l->14	
er bl	.->1	a->1	i->7	o->1	y->1	
er bo	m->1	r->7	
er br	i->6	o->1	y->1	ö->1	
er bu	d->3	
er by	g->2	r->1	
er bä	s->2	t->1	
er bå	d->1	
er bö	r->10	
er ca	p->10	
er ci	r->1	t->1	
er da	g->4	n->1	t->1	
er de	 ->129	b->5	c->2	f->1	l->6	m->19	n->123	r->8	s->33	t->169	
er di	r->3	s->1	t->1	v->1	
er dj	u->2	ä->1	
er do	c->9	k->1	l->6	m->2	
er dr	a->3	
er du	b->2	m->1	
er dy	k->1	n->1	
er dä	r->23	
er då	 ->10	l->2	
er dö	d->1	l->1	
er ec	u->2	
er ed	 ->1	
er ef	f->6	t->14	
er eg	e->2	n->1	o->1	
er ej	 ->5	,->1	.->2	
er ek	o->7	
er el	l->36	v->1	
er em	e->12	o->2	
er en	 ->103	.->1	b->1	d->3	e->2	h->3	i->1	k->1	l->3	o->2	
er er	 ->11	,->1	a->1	t->1	
er et	n->1	t->58	
er eu	r->26	
er ex	a->1	e->3	p->2	t->2	
er fa	k->4	l->1	r->3	s->5	t->2	
er fe	d->1	m->2	
er fi	n->10	
er fl	e->8	y->2	
er fo	l->3	r->16	
er fr	a->47	i->2	ä->4	å->77	
er fu	l->4	
er fy	r->2	
er få	 ->4	r->11	
er fö	l->4	r->303	
er ga	m->1	r->2	
er ge	 ->1	m->10	n->21	r->1	s->2	
er gi	v->3	
er gj	o->1	
er gl	o->1	ö->1	
er go	d->7	l->1	
er gr	a->4	u->4	ä->10	
er gy	n->3	
er gä	l->3	
er gå	r->8	
er gö	r->12	
er ha	 ->5	l->2	m->2	n->9	r->61	
er he	l->35	r->1	
er hi	n->1	s->2	t->1	
er hj	ä->1	
er ho	n->6	s->4	
er hu	n->1	r->18	v->10	
er hy	s->1	
er hä	m->1	n->4	r->11	
er hå	l->2	
er hö	g->3	r->2	
er i 	-->1	A->1	B->3	C->1	D->1	E->12	F->3	K->4	M->1	S->3	U->2	a->10	b->6	d->49	e->10	f->23	g->6	h->4	i->1	j->1	k->7	l->2	m->11	n->3	o->6	p->4	r->5	s->18	t->1	u->5	v->14	Ö->4	ö->2	
er ic	k->1	
er if	r->3	
er ig	e->5	n->1	
er ih	o->1	
er il	l->2	
er im	m->1	
er in	 ->6	b->2	c->1	d->2	f->4	g->16	i->2	k->2	l->1	n->7	o->38	r->9	s->4	t->134	v->3	
er ir	l->1	
er ja	,->1	g->103	
er jo	r->3	
er ju	 ->6	,->1	d->1	l->1	s->1	
er jä	m->2	r->2	
er ka	l->1	m->2	n->23	r->1	t->5	
er ke	m->1	
er kl	a->2	i->1	
er kn	a->2	
er ko	l->2	m->70	n->31	r->3	s->4	
er kr	a->8	i->6	y->1	ä->3	
er ku	b->1	l->2	n->2	r->1	s->1	
er kv	a->2	i->3	
er kä	m->1	n->5	r->2	
er kö	l->1	
er la	g->6	n->1	s->1	
er le	d->8	g->1	v->1	
er li	g->3	k->10	v->2	
er lo	k->1	v->1	
er lu	g->2	
er ly	c->2	
er lä	g->3	k->1	m->3	n->4	s->2	t->1	
er lå	n->12	t->2	
er lö	n->2	s->1	
er ma	i->3	k->1	l->2	n->35	r->3	t->2	
er me	d->110	k->1	l->11	n->7	r->9	t->2	
er mi	g->51	l->7	n->18	s->1	t->3	
er mo	b->1	d->1	r->1	t->18	
er mu	t->1	
er my	c->13	n->2	
er mä	n->9	
er må	l->2	n->9	s->22	
er mö	j->7	t->2	
er na	t->8	
er ne	d->2	j->2	r->1	
er ni	 ->25	v->1	
er no	g->1	r->1	
er nu	 ->8	,->1	m->1	
er ny	 ->1	a->2	h->1	
er nä	m->2	r->20	s->6	
er nå	g->24	
er oa	c->1	v->1	
er ob	a->1	e->1	
er oc	h->352	k->55	
er of	f->1	r->1	t->3	
er ok	l->1	
er ol	a->1	i->2	j->1	y->1	
er om	 ->102	f->4	k->9	l->1	r->3	s->1	
er or	d->5	i->1	o->7	s->1	ä->1	
er os	s->52	
er ou	n->1	
er oö	v->1	
er pa	r->9	s->1	
er pe	n->2	r->5	
er pl	a->2	e->1	u->1	
er po	l->4	s->3	
er pr	a->2	e->1	i->3	o->18	ä->1	ö->1	
er pu	n->3	
er på	 ->151	,->3	.->3	b->1	l->1	m->2	v->1	
er ra	d->2	k->2	p->3	s->2	t->1	
er re	a->2	c->1	d->3	f->4	g->17	j->1	k->2	l->1	n->1	s->6	
er ri	g->1	k->2	m->1	s->6	
er ro	p->1	
er ru	m->2	t->1	
er rä	k->2	t->9	
er rå	d->12	
er rö	r->5	s->2	
er sa	d->1	g->2	k->3	m->32	
er se	 ->1	d->4	k->3	n->6	r->1	s->1	x->1	
er si	d->1	g->60	n->19	t->10	
er sj	u->1	ä->10	
er sk	a->39	i->1	j->1	r->1	u->7	y->3	ä->1	
er sl	u->5	ä->1	
er sm	å->2	
er sn	a->2	e->1	
er so	c->1	m->392	v->1	
er sp	e->7	i->1	o->1	r->1	
er st	a->21	e->1	o->14	r->4	ä->3	å->6	ö->4	
er su	b->1	
er sv	a->2	å->2	
er sy	f->1	m->3	n->5	s->2	
er sä	k->7	r->5	t->1	
er så	 ->26	,->1	d->2	l->4	s->3	v->1	
er sö	n->3	
er t.	e->1	
er ta	 ->1	g->2	l->10	n->2	r->1	
er ti	d->6	l->154	o->2	t->1	
er tj	ä->2	
er to	g->2	l->4	n->2	p->1	r->2	t->2	
er tr	a->3	e->9	o->5	y->2	ä->6	
er tu	n->1	r->1	
er tv	e->2	i->5	ä->1	å->4	
er ty	d->1	n->1	v->1	
er tä	n->1	
er un	d->28	g->2	i->6	
er up	p->35	
er ur	 ->3	s->1	
er ut	 ->12	,->2	.->2	?->1	a->28	b->3	e->2	f->5	g->1	i->1	k->1	n->1	r->1	s->2	t->2	v->4	ö->2	
er va	d->14	k->1	l->4	r->39	t->1	
er ve	d->1	k->1	m->1	r->5	t->8	
er vi	 ->109	,->1	d->14	k->2	l->16	s->14	t->3	
er vo	l->1	n->1	
er vä	g->1	l->7	n->2	r->4	
er vå	l->1	r->21	
er yt	t->1	
er Ös	t->4	
er äl	d->1	
er äm	n->2	
er än	 ->49	d->13	n->4	
er är	 ->57	e->1	
er äv	e->13	
er år	 ->14	,->1	e->3	t->1	
er åt	 ->4	a->2	e->6	f->1	m->3	t->1	
er ök	a->3	
er ön	s->1	
er öp	p->5	
er ör	e->1	
er öv	e->23	r->1	
er! D	e->15	i->1	
er! E	f->2	u->4	
er! F	ö->4	
er! G	o->1	r->1	
er! I	 ->7	
er! J	a->15	ä->1	
er! K	a->1	
er! L	å->2	
er! M	e->1	
er! N	ä->1	
er! P	å->1	
er! S	o->1	
er! T	a->1	i->2	
er! U	n->1	
er! V	i->5	å->1	
er! Ä	v->2	
er! Å	r->1	
er!"D	e->1	
er!"O	m->1	
er!De	 ->3	t->2	
er!Ef	t->1	
er!Ja	g->3	
er!My	c->1	
er!Vi	 ->2	
er" h	a->1	
er" m	å->1	
er" s	o->2	
er"),	 ->1	
er", 	s->1	
er".D	e->1	
er) B	o->1	
er) V	i->1	
er) o	c->2	
er)Fr	u->2	
er)Ja	g->1	
er)Ko	n->1	
er)Ta	c->1	
er, "	n->1	
er, M	a->1	
er, T	h->1	
er, a	c->1	d->1	l->4	n->2	t->13	v->3	
er, b	a->1	e->5	l->3	o->1	r->1	å->2	
er, d	e->10	i->1	j->1	v->4	ä->9	å->4	ö->1	
er, e	f->5	l->2	n->11	t->2	x->2	
er, f	i->1	r->8	ö->17	
er, g	e->5	å->1	ö->1	
er, h	a->9	e->10	o->1	u->2	ä->1	
er, i	 ->9	b->1	n->14	
er, j	a->4	
er, k	a->2	o->5	r->2	u->1	ä->2	
er, l	a->1	e->2	i->2	o->1	
er, m	a->1	e->37	i->2	o->2	y->1	ä->2	å->3	
er, n	e->1	o->1	y->1	ä->4	å->5	
er, o	c->54	m->7	r->2	
er, p	l->1	r->3	å->3	
er, r	e->2	o->1	å->1	ö->1	
er, s	a->2	e->1	k->5	m->1	n->2	o->41	p->1	t->2	v->1	ä->5	å->11	
er, t	a->2	i->11	j->3	r->2	u->1	
er, u	n->2	p->3	t->14	
er, v	a->3	e->2	i->16	ä->1	å->1	
er, ä	n->1	r->7	v->2	
er, å	t->3	
er, ö	v->1	
er-bi	l->1	
er-ko	m->1	
er-na	t->1	
er-pr	o->11	
er-re	g->1	
er. (	F->1	
er. D	e->4	
er. E	n->1	u->1	
er. F	r->1	
er. H	e->1	
er. J	a->1	
er. M	a->1	e->1	
er. S	y->1	å->1	
er. T	i->1	
er. V	i->1	
er. Ä	n->1	
er.(A	p->1	
er.(I	T->1	
er.) 	H->1	
er.- 	(->2	H->1	
er.. 	(->1	
er..(	E->1	N->1	
er..H	e->1	
er..V	i->1	
er.90	 ->1	
er.Al	l->2	t->1	
er.An	t->1	
er.At	t->3	
er.Av	 ->4	
er.Ba	r->1	
er.Be	d->2	t->4	
er.Bl	a->1	
er.CS	U->1	
er.Da	g->1	
er.De	 ->11	n->23	s->5	t->75	
er.Do	m->1	
er.Dä	r->7	
er.Då	 ->1	
er.EU	-->2	
er.Ef	t->1	
er.En	 ->8	l->2	
er.Et	t->4	
er.Eu	r->5	
er.Ex	e->1	
er.Fr	a->1	i->1	u->5	å->2	
er.Få	r->1	
er.Fö	r->16	
er.Ge	n->3	
er.Ha	n->1	
er.He	r->11	
er.Hä	n->1	r->5	
er.I 	E->1	H->1	I->1	b->1	d->5	e->2	f->1	j->1	m->1	r->2	v->1	
er.In	g->2	o->3	
er.It	a->1	
er.Ja	g->59	
er.Ka	n->1	r->1	
er.Ki	n->1	
er.Ko	d->1	m->14	n->4	
er.Kv	i->1	
er.Li	k->1	
er.Lå	t->4	
er.Ma	n->1	
er.Me	d->5	n->11	r->1	
er.Mi	n->3	
er.Mä	n->1	
er.Na	t->2	
er.Nu	 ->1	
er.Nä	r->9	
er.Oc	h->3	k->1	
er.Om	 ->8	r->1	
er.Or	d->1	o->1	
er.Pa	r->2	
er.Pl	a->1	
er.Pr	o->3	
er.Pu	n->1	
er.På	 ->1	
er.Re	d->1	v->1	
er.Rå	d->1	
er.Sa	m->2	
er.Sl	u->2	
er.So	m->4	
er.St	a->1	o->1	r->1	ö->1	
er.Så	d->1	l->1	
er.Ta	c->3	
er.Te	r->1	
er.Ti	l->11	
er.Tr	o->1	
er.Un	d->5	i->1	
er.Va	d->7	l->1	r->4	
er.Vi	 ->34	s->1	
er.Vå	r->1	
er.Än	d->2	
er.Är	 ->3	
er.Äv	e->4	
er.Å 	a->2	
er: "	J->1	
er: A	n->1	
er: D	e->1	
er: I	n->1	
er: K	ä->1	
er: V	i->2	
er: a	t->1	
er: d	e->4	
er: e	n->2	
er: f	ö->1	
er: i	n->1	
er: k	o->1	
er: v	i->2	
er; a	t->1	
er; d	e->2	å->1	
er; e	n->1	
er; o	c->1	
er; v	i->1	
er?- 	(->1	
er?. 	(->1	
er?Bo	r->1	
er?De	t->1	
er?Eu	r->1	
er?He	r->3	
er?Ja	g->1	
er?Ko	m->1	
er?Me	n->1	
er?På	 ->1	
er?Ta	c->1	
er?Ve	m->1	
er?Vi	 ->1	
er?Äv	e->1	
erHer	r->1	
erJag	 ->1	
erMed	 ->1	
erNäs	t->2	
era -	 ->3	
era 2	5->1	
era E	U->2	u->5	
era F	N->1	
era I	n->1	s->1	
era L	o->1	
era a	l->5	n->5	r->2	s->1	t->38	v->11	
era b	e->4	i->1	o->1	r->1	u->1	ä->2	å->1	
era c	e->1	
era d	a->2	e->86	i->1	
era e	f->3	g->2	l->1	n->27	r->5	t->19	u->1	x->2	
era f	e->1	i->1	l->2	o->3	r->10	u->1	ö->23	
era g	e->5	r->1	å->10	
era h	a->1	e->5	i->1	o->3	u->6	ö->1	
era i	 ->12	n->10	
era j	ä->1	
era k	l->1	o->21	v->2	
era l	a->2	e->2	i->2	ä->3	ö->1	
era m	a->2	e->10	i->10	o->3	y->1	ä->2	å->4	ö->1	
era n	a->2	e->1	y->1	ä->1	å->1	
era o	b->1	c->21	f->1	k->1	l->5	m->9	p->1	r->7	s->4	
era p	a->4	e->1	o->6	r->6	u->1	å->17	
era r	e->13	i->1	å->1	
era s	a->2	e->2	i->13	k->4	n->4	o->3	p->1	t->4	y->1	ä->4	å->6	
era t	i->9	j->1	o->1	r->2	v->5	
era u	n->4	p->1	t->7	
era v	a->6	e->1	i->8	ä->4	å->3	
era Ö	s->2	
era ä	g->1	n->4	r->2	
era å	r->4	t->1	
era ö	s->1	v->10	
era! 	D->1	
era".	.->1	
era, 	a->3	f->2	h->1	m->1	o->1	u->1	v->1	ä->2	
era. 	M->1	
era.B	a->1	
era.D	e->3	ä->2	
era.E	n->2	
era.F	ö->1	
era.H	e->1	ä->1	
era.I	 ->2	
era.J	a->6	
era.L	ä->1	å->1	
era.M	e->2	i->1	
era.P	å->1	
era.V	i->1	
erad 	a->7	b->3	d->1	e->4	f->5	g->1	i->9	k->4	m->6	o->1	p->4	r->1	s->6	t->4	u->1	v->3	y->1	ä->1	ö->3	
erad,	 ->2	
erad.	D->1	M->3	U->1	V->1	
erade	 ->137	,->4	.->5	s->16	
erahu	s->1	
eral 	I->2	p->1	s->1	å->1	
erala	 ->24	,->1	
erald	e->1	i->17	
erale	n->1	r->2	
erali	s->12	
erall	t->9	
erals	e->2	
eralt	 ->4	
eran-	 ->1	
eranb	i->8	
erand	e->55	
erans	 ->4	,->3	.->2	e->1	k->2	
erant	ö->3	
eranv	ä->18	
erar 	-->1	1->1	3->1	E->1	I->1	a->24	b->4	d->37	e->19	f->9	g->1	h->11	i->30	j->11	k->7	l->1	m->17	n->7	o->10	p->9	r->3	s->18	t->5	u->3	v->11	ä->3	ö->4	
erar!	T->1	
erar,	 ->9	
erar.	.->1	A->1	D->1	F->3	H->1	N->1	S->1	V->1	
erare	 ->1	,->2	s->1	
erark	i->4	
erart	r->1	
eras 	4->1	E->1	a->32	b->2	c->2	d->6	e->12	f->16	g->5	h->2	i->31	k->5	l->5	m->8	n->5	o->17	p->13	r->5	s->22	t->8	u->6	v->4	ä->3	å->2	ö->2	
eras,	 ->13	
eras.	 ->1	D->6	F->4	I->2	J->1	M->1	P->1	S->1	V->4	Y->1	
erat 	-->2	E->1	a->8	b->4	d->13	e->5	f->7	g->1	h->4	i->7	k->3	l->2	m->4	n->3	o->7	p->1	r->1	s->10	t->2	v->4	å->1	
erat,	 ->11	
erat.	 ->1	.->1	D->1	E->1	J->3	K->1	T->1	V->1	
erat;	 ->1	
erati	o->9	v->6	
erato	g->2	
erats	 ->21	,->3	.->1	?->1	
eratu	r->13	
eratö	r->2	
eray,	 ->1	
erb, 	e->1	
erbal	a->1	
erbar	 ->1	a->2	
erbay	e->1	
erbel	a->3	
erbem	a->1	
erber	 ->2	,->3	n->2	
erbet	a->1	ä->6	
erbil	d->1	
erbis	k->6	
erbju	d->19	
erbjö	d->1	
erbli	c->1	
erblå	s->2	
erbri	n->1	
erbry	g->3	
erböl	d->1	
erbör	a->1	l->10	
ercen	t->1	
erdam	 ->9	,->3	.->1	f->27	r->1	
erdel	a->2	n->2	
erdo 	R->1	
erdom	l->1	s->1	
erdri	f->1	v->13	
erdst	o->3	
erdör	r->1	
ere a	n->1	
ere k	r->1	
ere.M	e->1	
ereda	 ->7	,->1	n->2	
eredd	 ->20	a->13	e->2	
erede	l->5	r->7	
ereds	 ->1	k->1	
eregl	e->3	
erell	 ->3	a->6	t->7	
erend	 ->4	!->2	,->2	-->1	b->1	s->2	
ereng	u->2	
erens	 ->60	,->8	.->7	?->2	e->129	k->18	r->1	s->21	
erent	i->5	
erera	 ->4	d->2	r->6	s->6	t->1	
ererö	v->1	
eresu	r->1	
eret 	s->1	
eret,	 ->1	
erett	 ->4	.->1	s->1	
erext	r->6	
erfal	l->3	
erfar	e->23	i->2	n->1	t->1	
erfek	t->7	
erfin	n->3	
erfir	a->2	
erfis	k->1	
erfly	t->2	
erflö	d->1	
erfor	d->5	s->22	
erfrå	g->8	
erfun	n->2	
erföl	j->3	l->2	
erför	a->5	d->1	e->2	i->12	t->1	v->1	
erg f	ö->1	
erg g	j->1	
erg k	r->1	
erg o	m->1	
ergav	s->2	
erge 	e->1	v->2	
ergen	 ->1	s->4	
erger	 ->15	,->2	.->2	M->1	b->1	i->1	
erges	 ->2	,->1	
ergi 	b->1	g->2	h->1	l->1	m->1	o->4	s->3	
ergi,	 ->2	
ergi-	,->1	
ergi.	A->1	E->2	F->1	M->1	
ergia	g->1	n->6	
ergib	e->3	
ergic	e->1	
ergie	f->4	
ergif	o->1	t->2	ö->4	
ergii	m->1	
ergik	a->1	o->1	ä->37	
ergim	i->1	y->1	
ergin	 ->3	,->1	
ergio	r->2	
ergip	o->2	r->5	
ergis	e->4	k->1	n->1	ä->7	
ergiv	e->4	l->1	n->3	
ergiä	k->1	
ergiå	t->1	
ergne	 ->1	
ergri	p->14	
ergru	p->1	
ergrä	v->4	
ergäl	l->1	
ergå 	t->1	
ergån	g->11	
ergår	 ->3	
ergåt	t->1	
erhan	d->6	
erhea	d->1	
erhet	 ->133	,->12	.->24	?->3	J->1	e->46	s->62	
erheu	g->2	
erhus	 ->1	e->1	
erhäm	t->2	
erhän	g->1	
erhål	l->12	
erhög	h->2	
erhöl	l->3	
erhör	d->3	t->9	
eri -	 ->1	
eri a	v->1	
eri f	ö->2	
eri i	 ->1	
eri k	o->1	
eri m	e->1	o->1	
eri n	ä->1	
eri o	c->5	
eri ä	r->2	
eri ö	k->1	
eri, 	d->1	e->1	l->2	m->2	n->1	
eri- 	o->1	
eri.J	a->1	
eri.L	i->1	
eri.M	a->1	
erial	 ->12	,->2	.->5	e->4	
eribe	k->4	
eriel	l->4	
erien	 ->1	
erier	 ->23	,->3	.->2	n->11	
eries	m->1	
eriet	 ->5	.->3	s->1	
erife	r->6	
erifi	e->1	
erige	 ->5	.->2	n->19	
erika	 ->6	,->1	n->17	r->1	s->1	
eriko	m->1	n->1	
eril 	u->1	
erila	g->1	
erims	a->2	b->2	p->1	r->2	å->1	
erimå	l->1	
erin 	s->1	
erin.	J->1	
erinf	ö->4	
ering	 ->197	!->1	"->2	)->1	,->28	.->37	;->1	?->1	a->96	e->119	s->227	å->1	
erinr	a->13	e->1	ä->1	
erins	e->1	t->8	
erint	a->1	
erinä	r->3	
eriod	 ->23	,->5	.->2	?->1	e->41	i->14	
eripo	l->1	
erise	k->2	r->2	
erisk	a->1	
erite	r->1	
eriut	s->1	
eriös	 ->1	a->3	t->4	
erk -	 ->1	
erk a	t->1	
erk b	y->1	
erk f	i->1	å->1	ö->1	
erk g	e->1	
erk i	 ->5	n->3	
erk k	a->1	
erk m	e->2	
erk o	c->1	
erk p	å->1	
erk s	e->1	o->3	
erk u	t->1	
erk ä	r->2	
erk, 	g->1	m->1	s->1	
erk.B	e->1	
erk.D	e->1	
erk.S	y->1	
erk.V	a->1	
erk?R	e->1	
erka 	a->1	b->1	d->3	e->1	f->10	h->1	i->5	k->1	m->1	n->1	o->1	p->1	r->1	s->4	t->4	u->1	v->1	ä->1	å->1	
erka,	 ->1	
erkad	e->2	
erkan	 ->18	,->1	.->1	d->1	
erkar	 ->57	a->5	e->25	n->34	
erkas	 ->8	,->1	t->2	
erkat	 ->3	,->1	e->2	s->5	
erken	 ->5	,->1	
erket	 ->33	,->5	s->2	
erkla	g->6	
erkli	g->205	
erkni	n->15	
erkom	m->6	s->1	
erkra	n->1	
erkrä	v->1	
erksa	m->51	n->1	
erkst	ä->19	
erkty	g->8	
erkur	s->1	
erkän	d->5	n->35	t->2	
erlag	 ->4	,->1	.->2	t->1	
erlev	a->2	e->3	n->4	s->1	
erlig	 ->5	,->1	a->60	e->38	g->1	h->2	t->7	
erlin	 ->4	,->2	.->1	
erlys	e->1	t->1	
erläg	g->5	s->2	
erläm	n->18	
erlän	d->18	
erlät	t->18	
erlåt	a->6	e->2	i->2	s->1	
ermaj	o->1	
erman	.->1	e->8	s->1	
ermat	e->1	
ermen	i->1	
ermer	 ->2	,->1	
ermid	d->9	
ermin	e->1	
ermis	.->1	
ermo,	 ->1	
ermod	i->1	
ermor	g->1	
ermål	i->1	
ermöt	e->2	
ern (	f->1	
ern -	 ->1	
ern E	r->2	
ern b	i->1	
ern d	e->1	
ern e	n->1	
ern f	r->1	ö->5	
ern g	r->1	
ern h	a->3	
ern i	 ->2	n->1	
ern k	o->3	
ern l	i->2	
ern m	e->1	
ern n	y->1	
ern o	c->7	m->2	
ern p	å->1	
ern r	e->1	
ern s	a->1	k->2	o->2	å->1	
ern t	a->1	o->1	
ern u	n->1	
ern v	a->1	i->1	
ern ä	r->1	
ern, 	B->1	R->1	h->1	i->2	j->1	m->1	s->1	v->1	
ern.)	 ->1	
ern..	 ->1	
ern.D	e->3	ä->1	
ern.H	e->1	
ern.J	a->1	u->1	
ern.O	m->1	
ern.V	i->1	
ern.Ö	g->1	
ern/N	o->2	
erna 	(->1	-->14	1->4	A->1	I->1	P->1	T->1	a->65	b->26	d->14	e->17	f->135	g->20	h->41	i->132	j->3	k->31	l->7	m->55	n->8	o->125	p->21	r->11	s->84	t->39	u->30	v->17	ä->36	å->3	ö->5	
erna!	D->1	H->1	
erna"	.->1	
erna,	 ->168	
erna.	 ->4	)->1	-->1	.->1	A->8	B->2	D->38	E->9	F->6	G->2	H->7	I->11	J->19	K->7	L->3	M->14	N->6	O->4	P->5	R->1	S->8	T->3	U->2	V->27	Ä->2	Å->1	
erna/	s->1	
erna:	 ->3	
erna;	 ->4	
erna?	H->1	I->1	J->1	M->1	V->3	Ä->1	
ernaH	e->1	
ernar	d->1	e->1	
ernas	 ->144	,->1	.->1	
ernat	i->94	
ernd 	L->3	
ernea	r->1	
erner	 ->1	i->1	n->1	
ernet	 ->4	,->4	.->2	
ernfr	e->1	
ernis	e->24	
ernit	i->1	
erniv	å->1	
ernié	 ->1	
erns 	d->1	f->2	h->1	n->1	o->2	p->2	s->2	u->1	v->1	
ernt 	s->3	u->1	
ernt.	S->1	
erntu	n->1	
ernör	,->1	
erodd	e->5	
eroen	d->69	
eroga	t->1	
erois	k->1	
eromr	å->1	
eroni	.->1	
eropa	r->1	
eror 	a->1	i->4	j->1	m->1	o->1	p->8	t->2	
eror,	 ->1	
erord	n->5	
erott	 ->1	
erpar	l->1	t->1	
erpol	i->1	
erpop	u->1	
erpos	t->2	
erpre	s->1	
erpri	s->1	
err A	l->1	
err B	a->2	e->5	o->3	
err C	o->3	
err E	v->2	
err F	r->1	
err G	o->1	r->1	
err H	ä->2	
err J	o->1	
err K	i->4	o->2	
err L	a->1	
err M	o->1	
err N	o->1	
err P	a->3	o->5	
err R	a->1	
err S	c->2	e->2	p->1	
err W	y->1	
err f	ö->5	
err g	e->1	
err k	o->82	
err l	e->15	
err m	i->2	
err o	r->5	
err p	a->3	
err r	å->12	
err t	a->319	j->1	
err v	a->3	
erran	d->2	
errar	 ->8	!->20	,->16	n->1	
erras	k->1	
erreg	e->3	l->2	
errep	r->2	
erres	 ->1	
errez	,->1	
errik	a->7	e->74	i->49	
errit	o->17	
erron	g->1	
error	.->1	i->10	
errät	t->1	
erråd	 ->1	,->1	e->12	
errón	 ->3	
errös	t->1	
ers a	l->1	n->7	r->2	
ers b	e->9	i->1	
ers e	k->2	r->1	
ers f	r->2	u->2	ö->1	
ers i	n->3	
ers j	u->1	
ers k	a->1	
ers l	e->1	i->2	ö->1	
ers n	a->1	
ers o	k->1	l->1	
ers p	a->5	o->1	
ers r	a->1	e->1	ä->2	
ers s	a->1	o->1	t->3	
ers t	y->1	
ers u	p->1	t->4	
ers v	a->2	
ers å	s->1	
ers ö	p->1	
ers, 	L->1	
ers-b	i->1	
ersai	l->1	
ersal	m->1	
ersam	l->1	m->1	t->1	
ersat	t->5	
erse 	k->1	o->1	
ersel	l->3	
ersen	 ->2	
erser	 ->1	
ershi	p->1	
ersie	l->9	
ersif	i->2	
ersik	t->18	
ersio	n->13	
erska	l->2	p->22	
ersko	t->1	
erskr	i->19	o->1	
erskå	d->6	
erslu	n->1	
ersmå	l->1	
ersom	 ->189	,->1	
erson	 ->6	,->1	a->23	e->43	l->34	s->1	
erspe	g->3	k->17	r->2	
erst 	a->1	d->1	f->1	i->1	k->1	m->1	n->1	p->1	s->2	v->8	
ersta	 ->17	t->5	
ersti	g->5	
erstr	e->1	y->27	ä->12	ö->2	
erstä	l->40	
erstå	e->1	r->13	
erstö	d->6	
ersun	d->3	
ersvä	m->7	
ersyn	 ->1	
ersät	t->35	
ersåt	e->1	
ersök	a->19	e->2	n->23	t->4	
ert C	a->1	
ert G	o->1	
ert a	t->1	
ert b	e->6	i->1	r->1	
ert d	j->1	
ert e	g->1	
ert f	a->1	ö->4	
ert g	e->1	o->1	
ert h	u->1	
ert i	 ->1	n->5	
ert k	a->1	o->2	ä->1	
ert l	ö->1	
ert m	e->1	
ert o	c->4	m->1	r->1	
ert p	a->4	
ert s	a->1	o->3	t->2	v->3	ä->1	
ert t	o->1	
ert u	t->5	
ert v	e->1	i->1	
ert y	t->1	
ert ä	m->1	n->2	
ert ö	g->1	
ert!J	a->1	
ert, 	e->2	m->2	
ert.J	a->1	
erta 	a->1	d->1	u->1	
ertag	,->1	a->8	n->1	
ertal	 ->2	a->1	e->4	
ertan	k->3	
ertar	 ->1	,->1	
ertas	 ->1	
ertec	k->17	
erter	 ->7	.->2	n->11	
ertgr	u->3	
erthe	t->1	
erthu	 ->1	
ertid	 ->64	,->3	
ertif	i->6	
ertik	a->3	
ertil	l->1	
ertin	o->1	
ertis	 ->1	,->1	.->1	
ertko	m->17	
ertog	 ->1	
erton	e->1	
ertra	k->1	m->1	p->1	
ertre	g->1	
erträ	d->6	f->1	
ertut	s->1	
ertyg	a->34	e->4	
ertän	k->2	
erupp	b->12	l->1	r->7	s->3	t->11	
erusa	l->2	
erutb	i->2	
erutv	e->1	
ervak	a->14	n->11	
ervat	i->9	s->1	ö->1	
ervec	k->1	
erven	e->2	t->5	
erver	 ->2	a->2	k->1	
ervic	e->7	
ervin	n->74	
ervis	a->1	
ervju	 ->2	a->1	
ervri	d->1	
ervtr	u->1	
ervun	n->3	
erväg	a->25	d->1	e->7	t->2	
erväl	d->3	
ervän	d->3	
ervär	d->5	l->1	t->1	
ery, 	H->1	
erykt	a->1	
eräga	r->1	
eräkn	a->2	i->2	
erän 	n->1	s->1	
eräna	 ->3	
eräni	t->12	
erätt	 ->2	a->9	e->4	i->20	
eråri	g->12	
eråt 	k->1	
erömt	 ->1	
erömv	ä->1	
erör 	P->1	a->1	d->1	f->1	k->1	o->3	s->1	
erörd	 ->2	a->18	e->1	
erörs	 ->8	
erört	 ->2	s->2	
erös 	o->1	p->1	
erösa	 ->1	
eröst	 ->2	
eröva	r->1	
erövr	a->2	
es - 	i->1	t->1	
es 19	5->1	6->1	9->1	
es 2 	4->1	
es 3,	8->1	
es Ad	o->1	
es De	l->3	
es Gi	l->1	
es Sp	a->1	
es Vi	c->1	
es Wi	e->1	
es al	l->1	
es an	g->1	s->6	
es ar	b->2	
es at	t->9	
es au	k->1	
es av	 ->24	g->2	s->1	
es ba	r->1	
es be	f->1	l->1	t->2	v->1	
es bl	i->1	
es bo	r->1	
es br	å->1	
es by	r->1	
es bä	t->1	
es de	 ->2	l->1	m->1	n->4	t->6	
es di	t->1	
es dä	r->3	
es då	 ->1	
es dö	d->1	
es eg	e->1	
es ek	o->1	
es el	l->6	
es em	e->1	o->1	
es en	 ->4	v->1	
es et	 ->1	t->4	
es fa	s->1	
es fi	n->1	s->1	
es fl	e->1	
es fo	l->2	r->1	
es fr	a->2	å->9	
es fö	r->24	
es ge	n->2	
es gö	r->1	
es ha	 ->2	d->1	r->2	
es he	l->1	
es hi	s->1	
es hä	n->1	
es hå	r->1	
es hö	g->1	j->1	
es i 	A->2	B->1	E->1	G->2	J->1	M->1	S->4	T->2	a->1	d->4	e->1	f->1	g->2	h->2	j->1	k->2	m->3	p->2	r->2	s->2	
es ig	e->1	
es ih	o->1	
es in	 ->1	,->1	g->2	n->1	r->2	s->1	t->7	
es ju	s->2	
es kl	.->2	a->2	
es ko	l->1	m->5	n->1	
es kr	i->1	
es ku	n->1	s->1	
es kv	o->1	
es le	d->3	t->1	
es lo	b->1	
es ma	k->1	n->2	
es me	d->5	
es mo	t->2	
es my	c->1	
es mö	j->4	
es na	c->1	
es no	g->1	
es ny	a->2	l->3	s->1	
es nå	g->2	
es nö	d->2	
es ob	l->1	
es oc	h->10	k->4	
es of	ö->1	
es om	 ->3	r->1	
es or	o->1	
es ph	a->1	
es po	r->1	s->1	
es pr	e->1	o->1	
es på	 ->5	
es re	d->2	g->2	s->1	
es ri	k->2	
es ro	t->1	
es ry	k->1	
es rä	k->1	t->4	
es rö	r->1	s->1	
es sa	m->1	
es se	 ->1	
es si	t->1	
es sj	ä->1	
es sk	u->1	
es sl	o->2	
es so	m->9	
es sp	e->2	
es st	a->1	o->1	r->1	å->1	
es sv	a->1	
es sä	r->1	
es ti	d->3	l->11	
es tj	ä->1	
es tv	i->1	ä->1	
es ty	d->3	
es un	d->3	
es up	p->6	
es ur	 ->1	
es ut	 ->1	a->1	g->1	m->1	r->1	
es va	n->1	r->2	
es vi	 ->1	d->1	l->2	s->1	
es vo	t->1	
es vä	c->1	g->2	
es yt	t->1	
es än	d->2	
es är	 ->2	
es åt	g->1	
es ög	o->1	
es ök	a->1	
es öv	e->5	
es".K	a->1	
es, W	u->1	
es, a	t->1	
es, e	f->1	n->1	
es, g	ö->1	
es, j	a->2	o->1	
es, o	c->5	m->1	
es, s	o->1	
es, t	.->1	
es, v	a->1	
es- o	c->6	
es-Ca	r->1	
es.)Å	t->1	
es.An	t->1	
es.De	t->1	
es.Dä	r->1	
es.Fl	o->1	
es.Hu	v->1	
es.I 	d->1	
es.Ja	g->1	
es.Ko	m->1	
es.Me	l->1	
es.Mä	n->1	
es.Om	 ->1	
es.Re	d->1	
es.Rå	d->1	
es.Un	d->1	
es.Va	d->1	
es.Vi	 ->1	
es; o	c->1	
esa b	e->1	
esa d	r->1	
esa e	r->1	
esa f	a->1	
esa i	 ->2	n->1	
esa m	i->1	
esa o	c->3	
esa p	å->1	
esa t	i->1	
esa ö	v->1	
esa, 	f->1	g->1	
esa.J	a->1	
esamm	a->7	
esan 	o->1	
esarb	e->1	
esare	 ->1	
esats	,->1	e->6	
esaur	o->1	
esbed	ö->1	
esbes	t->1	
esdig	r->2	
ese i	 ->1	
esegr	a->2	
esekt	o->3	
esen 	i->1	
esent	 ->1	.->1	a->23	e->23	
eser 	f->1	i->1	t->1	
eser,	 ->1	
esern	a->1	
eserv	a->2	e->3	t->1	
eseti	k->1	
esfor	m->1	
esfrå	g->4	
esför	s->1	
esgem	e->1	
esgil	l->1	
esgå 	K->1	d->1	
esgås	:->1	
eshan	d->4	
eside	n->9	
esidi	g->5	
esidu	e->1	
esikt	n->2	
esisk	 ->2	a->10	
esitt	e->2	
eskad	e->1	
eskap	 ->18	,->1	.->3	e->89	s->2	
eskar	r->1	
eskat	t->5	
esked	 ->3	
eskif	t->3	
eskre	v->3	
eskri	f->13	v->35	
eskva	l->1	
eskyd	d->3	
eskyl	d->1	l->2	
eskål	e->1	
eslag	e->1	i->14	n->10	r->1	
esliv	e->2	
eslog	 ->9	s->2	
eslut	 ->79	,->10	.->9	;->1	a->62	e->46	n->2	s->32	
esläk	t->1	
eslå 	a->5	e->3	k->3	p->1	r->1	s->1	v->1	
eslår	 ->35	"->1	.->1	?->1	
eslås	 ->16	
eslöt	 ->3	
esman	n->2	
esmin	i->9	
esmit	t->1	
esmän	 ->1	
esmär	k->1	
esmäs	s->1	
esnål	a->4	
esolu	t->100	
esona	n->1	
esone	m->3	
esor 	m->1	
esp. 	s->1	t->1	
espar	a->2	i->3	
espeg	l->1	
espek	t->80	
esper	i->7	
espo,	 ->1	
espol	i->3	
espon	d->1	s->1	
espos	 ->1	
esprå	k->9	
esque	,->1	
esrap	p->2	
esrör	e->1	
ess a	l->1	n->2	r->1	t->1	v->4	
ess b	e->4	i->1	r->1	u->1	
ess d	a->2	e->1	o->2	
ess e	g->3	k->1	n->1	x->1	
ess f	o->4	r->1	u->3	ö->3	
ess g	e->2	r->2	
ess h	a->1	i->1	
ess i	 ->3	n->8	
ess k	l->1	o->5	v->1	
ess l	a->1	i->2	
ess m	a->1	e->4	o->2	y->1	å->1	
ess n	a->2	y->1	ä->1	
ess o	c->1	m->1	r->4	
ess p	e->1	r->1	å->3	
ess r	e->4	y->1	ä->2	ö->1	
ess s	a->1	j->1	k->3	o->11	t->3	v->1	y->1	
ess t	i->2	o->1	
ess u	t->3	
ess v	i->1	ä->2	
ess ä	n->1	r->1	
ess å	s->2	t->1	
ess ö	d->1	r->1	
ess".	D->1	
ess, 	d->1	å->1	
ess.A	l->1	
ess.D	e->3	i->1	
ess.H	e->1	
ess.M	a->1	å->1	
ess.N	ä->1	
ess.V	i->3	å->1	
ess?J	o->1	
essa 	1->1	2->3	3->1	a->16	b->18	c->1	d->5	e->4	f->49	g->9	h->9	i->15	k->20	l->12	m->25	n->4	o->15	p->34	r->21	s->34	t->16	u->9	v->12	ä->24	å->8	ö->1	
essa!	L->1	
essa,	 ->4	
essa.	B->1	D->2	I->1	J->1	M->2	
essad	e->1	
essan	d->1	t->21	
essar	 ->1	
essbe	l->5	
esse 	(->1	a->6	d->3	f->5	l->1	o->1	p->1	s->2	t->1	
esse,	 ->5	
esse.	F->1	M->2	
esse?	E->1	
essen	 ->54	,->20	.->31	?->1	N->1	a->5	s->3	t->1	
esser	 ->4	,->2	a->13	n->6	
esset	 ->4	,->1	
esshä	n->1	
essim	i->2	
essio	n->9	
essiv	 ->2	a->3	t->3	
esska	t->1	
essko	n->2	
essme	d->1	
essni	n->1	
essor	 ->6	
essre	g->1	
essrä	t->2	
esstr	u->1	
essue	l->1	
essut	o->61	
essvä	r->4	
est M	i->1	
est a	c->1	n->3	v->3	
est b	e->3	
est d	e->1	r->2	y->1	
est e	f->1	
est f	r->2	ö->2	
est g	e->1	r->1	
est h	a->1	
est k	o->1	r->1	
est l	a->1	å->2	ö->1	
est m	o->2	
est n	ä->1	
est o	c->1	m->1	
est p	o->1	
est r	e->2	
est s	k->1	t->1	v->1	
est t	i->1	r->2	
est u	t->2	
est v	ä->1	
est ä	r->1	
est, 	s->1	
est?N	e->1	
esta 	a->7	d->2	f->2	h->2	i->2	k->1	m->2	s->4	t->2	v->1	ä->2	
esta,	 ->2	
estad	e->2	
estan	d->1	t->2	
estar	k->1	
estas	 ->1	
estat	e->1	i->4	
estau	r->1	
estei	n->1	
estel	s->3	
esten	 ->2	"->1	,->3	a->1	s->1	
ester	 ->4	"->1	.->1	a->8	f->2	i->12	n->4	
estie	r->1	
estin	a->10	i->4	s->8	
estni	n->1	
esto 	h->1	v->1	
estod	 ->1	
estor	e->3	
estra	f->2	t->1	
estri	d->2	k->4	
estru	k->1	
estrå	l->1	
ests.	D->1	
estun	d->7	
estyr	k->1	
estäl	l->16	
estäm	d->15	m->127	s->1	t->16	
estän	d->2	g->4	
estå 	a->4	
eståe	l->1	n->10	
estån	d->28	
estår	 ->18	
estör	t->1	
esult	a->109	e->7	
esurs	b->1	e->46	f->1	s->1	t->1	
esutb	i->7	
esval	,->1	
esvar	a->17	
esvik	e->7	n->1	
esvis	 ->2	
esvär	e->1	l->6	
esynn	e->1	
esyst	e->1	
esätt	:->1	e->2	n->3	
esök 	i->5	o->1	
esöka	 ->1	
esöke	t->1	
esökt	e->1	
esörj	a->2	
et "E	U->1	
et "K	u->2	v->1	
et "O	l->1	
et "e	g->1	n->1	u->1	
et "k	u->1	
et "r	e->2	
et (B	5->2	
et (C	E->1	
et (E	U->2	
et (F	P->1	
et (I	C->1	F->1	
et (S	P->1	
et (a	r->1	
et (d	e->1	
et (f	i->2	
et (h	ä->1	
et (i	 ->1	n->1	
et (k	o->1	
et (t	y->1	
et (Ö	V->1	
et , 	d->1	
et - 	a->4	d->3	e->2	f->1	g->1	h->1	i->2	k->2	m->1	o->5	p->1	s->5	u->1	v->3	ä->1	
et 19	4->1	9->13	
et 21	:->1	
et 22	 ->1	
et AB	B->1	
et Ak	k->1	
et Al	e->1	t->2	
et BN	P->1	
et Be	r->1	
et Br	e->1	
et Ca	s->1	
et Da	l->1	
et De	 ->1	
et EU	-->1	
et El	l->1	
et Eq	u->8	
et Er	i->1	
et Eu	r->4	
et Fö	r->1	
et Gr	e->1	ö->1	
et I 	T->1	
et It	a->1	
et Ko	s->1	
et Ku	l->3	
et Le	a->2	
et Mi	n->1	
et Mo	r->3	
et Po	r->4	
et RI	N->1	
et Ra	n->1	
et SE	M->1	
et Sa	v->1	
et Sj	u->1	
et St	o->1	
et Sv	e->1	
et TV	-->1	
et Tu	r->1	
et Va	t->1	
et Ve	r->1	
et Vo	d->1	
et ab	s->4	
et ac	c->4	
et ak	t->6	u->1	
et al	d->1	l->31	
et am	b->2	
et an	d->56	g->6	l->3	n->6	s->15	t->14	v->4	
et ar	a->1	b->22	t->1	
et at	t->258	
et av	 ->306	b->2	d->1	g->3	h->1	s->20	t->4	
et ba	d->1	k->1	r->13	
et be	a->2	d->2	f->6	g->5	h->18	k->6	l->4	r->18	s->13	t->37	v->1	
et bi	d->1	l->2	s->1	t->1	
et bl	.->1	a->2	e->1	i->22	y->1	
et bo	r->6	
et br	a->9	i->5	å->2	
et bu	d->3	
et by	g->1	r->2	
et bä	s->7	t->4	
et bå	t->1	
et bö	r->25	
et ce	m->2	n->1	
et ch	a->1	
et ci	r->1	v->4	
et da	g->3	n->7	t->5	
et de	 ->14	l->4	m->4	n->14	s->3	t->9	
et di	r->3	s->4	
et dj	ä->1	
et do	c->4	k->2	m->1	
et dr	a->4	ö->2	
et dy	r->2	
et dä	r->14	
et då	 ->11	l->3	
et dö	l->1	r->1	
et ef	f->1	t->11	
et eg	e->9	n->3	
et ek	o->8	
et el	e->2	l->19	
et em	e->3	
et en	 ->26	a->9	b->1	d->20	e->1	g->3	h->3	k->9	l->5	o->1	s->1	t->2	v->1	
et er	b->2	f->1	h->1	k->2	s->1	
et et	t->13	
et eu	r->31	
et ev	e->2	
et ex	 ->1	a->4	e->5	t->3	
et f.	d->1	
et fa	i->1	k->58	l->13	n->9	r->5	s->3	t->5	
et fe	l->1	m->11	
et fi	c->3	n->188	
et fj	ä->4	
et fl	e->3	y->1	
et fo	r->16	
et fr	a->18	i->7	u->1	ä->9	å->48	
et fu	l->4	n->5	
et fä	s->1	
et få	 ->4	r->21	t->1	
et fö	d->1	l->2	r->503	
et ga	m->3	n->1	r->1	v->3	
et ge	 ->1	m->9	n->14	o->2	r->10	s->1	
et gi	c->1	l->1	v->3	
et gj	o->4	
et gl	a->5	o->1	ä->8	
et go	d->18	t->3	
et gr	a->7	u->6	
et gy	n->1	
et gä	l->208	r->1	
et gå	r->14	t->3	
et gö	r->24	
et ha	 ->3	d->6	f->2	n->57	r->139	
et he	l->15	m->2	s->1	
et hi	n->3	s->1	t->4	
et hj	ä->2	
et ho	p->2	r->1	s->8	t->2	
et hu	r->1	s->1	
et hy	c->1	
et hä	n->12	r->56	
et hå	r->2	
et hö	g->8	j->1	l->2	r->4	
et i 	A->2	B->5	E->6	F->4	G->1	H->9	I->2	K->2	M->2	N->1	P->2	S->2	T->7	a->8	b->3	d->44	e->7	f->19	g->5	h->11	j->1	k->3	l->1	m->10	n->4	o->3	p->5	r->8	s->31	t->1	u->1	v->13	Ö->2	å->2	
et ib	l->3	
et id	e->1	
et ig	e->2	
et il	l->1	s->1	
et im	p->1	
et in	f->8	g->9	i->6	k->1	l->1	n->35	o->21	r->4	s->5	t->163	v->1	
et ir	l->1	r->2	
et it	a->3	
et ja	g->16	
et jo	r->1	
et ju	 ->6	r->2	s->7	
et jä	m->3	
et ka	l->1	n->59	p->2	
et ke	m->1	
et kl	a->12	
et kn	a->1	
et ko	l->1	m->109	n->13	r->7	s->4	
et kr	a->5	i->8	ä->32	
et ku	l->4	n->7	
et kv	a->6	
et ky	l->1	
et kä	m->1	n->8	
et kö	t->1	
et la	d->1	g->5	n->10	
et le	d->5	
et li	b->1	d->1	g->9	k->4	l->3	t->9	
et lo	g->2	
et lu	t->1	
et ly	c->1	d->1	s->1	
et lä	g->13	m->4	n->11	t->5	
et lå	g->2	n->5	
et lö	f->1	p->4	s->1	
et ma	k->2	n->9	t->2	
et me	d->157	l->32	n->7	r->12	s->7	
et mi	g->3	n->7	s->1	t->1	
et mo	d->4	n->1	t->20	
et mu	l->1	n->2	
et my	c->16	t->1	
et mä	r->1	
et må	h->1	l->4	n->3	s->77	
et mö	d->1	j->29	t->1	
et na	t->10	
et ne	g->2	
et ni	 ->8	
et no	g->8	r->2	t->1	
et nu	 ->24	,->2	v->9	
et ny	a->18	l->2	t->2	v->1	
et nä	m->2	r->19	s->2	
et nå	g->11	
et nö	d->12	j->1	
et oa	c->4	v->1	
et ob	e->3	
et oc	h->327	k->34	
et oe	r->1	
et of	f->5	t->3	ö->1	
et og	r->1	
et ok	l->1	
et ol	a->1	j->2	
et om	 ->90	f->3	r->8	s->2	v->1	ö->4	
et on	d->2	t->1	ö->1	
et op	r->1	t->1	
et or	d->1	g->2	o->8	s->1	w->1	
et os	a->1	ä->1	
et ot	i->1	y->1	ä->1	
et oö	v->1	
et pa	r->7	s->1	
et pe	k->1	n->2	r->5	
et pl	a->7	
et po	l->12	r->60	s->13	
et pr	a->5	e->1	i->1	o->9	
et på	 ->66	,->1	:->1	b->1	g->4	p->1	s->1	t->2	v->2	
et ra	k->3	t->1	
et re	a->1	d->11	e->1	f->2	g->7	k->2	n->1	s->6	t->3	
et ri	k->8	m->3	n->1	s->2	
et ry	k->1	
et rä	c->12	t->11	
et rå	d->21	k->1	
et rö	r->16	s->3	
et sa	d->2	k->12	m->19	n->6	t->1	
et se	 ->1	d->4	g->4	k->1	n->13	r->5	s->1	t->1	
et si	g->2	n->2	s->5	t->1	
et sj	u->2	ä->6	
et sk	a->68	e->15	i->2	r->4	u->69	ä->9	ö->1	
et sl	a->2	u->7	ä->2	å->1	
et sm	ä->1	å->1	
et sn	a->8	
et so	c->9	l->1	m->212	r->1	
et sp	a->4	e->12	
et st	a->21	e->1	i->1	o->31	r->8	ä->14	å->25	ö->23	
et su	b->2	n->1	
et sv	a->4	e->1	å->8	
et sy	f->6	m->1	n->3	s->8	
et sä	g->8	k->9	m->2	r->7	t->34	
et så	 ->23	,->1	.->2	d->2	g->1	l->3	s->2	v->2	
et sö	d->1	k->1	
et ta	 ->2	g->1	r->6	
et te	r->1	
et ti	b->1	d->9	l->109	o->1	
et tj	u->1	ä->1	
et to	g->1	t->2	
et tr	a->6	e->19	o->4	ä->4	
et tu	f->1	n->2	
et tv	e->2	i->5	å->1	
et ty	c->3	d->12	s->4	v->2	
et tä	n->6	
et tå	l->1	
et un	d->21	
et up	p->41	
et ur	s->3	v->1	
et ut	 ->1	a->11	e->2	f->1	g->10	h->1	l->1	m->4	s->5	t->7	v->2	ö->1	
et va	c->1	d->10	l->4	n->2	r->77	
et ve	r->20	t->7	
et vi	 ->37	d->18	k->70	l->55	s->16	t->2	
et vo	l->1	r->12	
et vä	l->26	n->2	r->5	s->3	x->2	
et vå	g->1	r->3	
et yt	t->7	
et Ös	t->1	
et äc	k->1	
et äg	e->1	n->2	
et äm	b->1	
et än	 ->4	,->1	d->15	n->5	t->2	
et är	 ->785	:->1	e->1	
et äv	e->13	
et ål	i->4	
et år	 ->3	e->1	h->1	l->1	
et åt	 ->7	a->2	e->10	m->1	
et öd	e->2	
et ög	o->1	
et ök	a->3	
et ön	s->2	
et öp	p->3	
et ös	t->14	
et öv	e->13	
et!(P	a->1	
et!. 	(->1	
et!.(	N->1	
et!He	r->1	
et!Ku	l->1	
et!Pr	e->1	
et" (	s->1	
et" g	ö->1	
et" m	e->1	
et" o	c->1	
et" ä	r->1	
et", 	b->1	s->1	
et".E	n->1	
et".J	a->1	
et) (	C->1	
et) C	5->1	
et) h	a->2	
et) p	å->1	
et) s	o->1	
et), 	d->1	s->1	t->1	
et).D	e->1	
et).H	e->2	
et).L	i->1	
et)Nä	s->1	
et, C	o->1	
et, D	a->1	
et, E	f->1	
et, G	i->1	
et, H	a->1	
et, I	I->2	n->1	
et, J	o->1	
et, W	e->1	
et, a	n->4	r->1	t->11	v->5	
et, b	e->2	l->2	ö->2	
et, d	e->27	v->4	ä->4	å->1	
et, e	f->8	l->1	n->8	t->2	x->1	
et, f	a->1	i->2	r->11	å->1	ö->19	
et, g	e->3	å->3	ö->1	
et, h	a->10	e->14	j->1	
et, i	 ->11	n->11	
et, j	a->3	ä->2	
et, k	a->4	o->9	u->1	ä->3	
et, l	a->1	e->1	i->1	ä->1	
et, m	e->33	i->1	o->1	y->3	ä->1	å->2	
et, n	a->3	ä->9	
et, o	a->2	c->51	l->1	m->12	
et, p	a->1	l->1	o->1	r->2	å->4	
et, r	a->1	e->1	ä->1	å->2	
et, s	a->1	e->3	k->5	o->35	p->2	t->2	ä->32	å->13	
et, t	a->1	i->2	v->1	y->3	
et, u	n->2	p->1	t->18	
et, v	a->9	e->2	i->20	o->1	ä->3	å->1	
et, ä	r->8	v->4	
et, å	 ->1	
et, ö	k->1	p->1	
et- o	c->1	
et-fr	å->1	
et. (	P->1	
et. D	e->7	ä->1	
et. E	t->1	
et. J	a->1	
et. K	o->1	
et. M	e->1	
et. S	o->1	
et. V	i->1	å->1	
et. a	i->1	
et.(A	r->1	
et.(F	R->1	
et.(P	T->1	
et.)A	n->1	
et.)B	e->2	
et.)R	e->1	
et.- 	H->1	
et.. 	(->2	
et...	F->1	
et.19	9->1	
et.Al	d->1	
et.An	s->1	v->1	
et.At	t->1	
et.Av	 ->3	s->5	
et.Be	t->2	
et.Bl	a->1	
et.Br	i->1	
et.De	 ->14	l->1	n->15	s->3	t->83	
et.Dä	r->9	
et.Då	 ->1	
et.EG	-->1	
et.Ef	f->1	t->3	
et.Ek	o->1	
et.En	 ->3	d->2	l->3	
et.Et	t->5	
et.Eu	r->9	
et.Fl	e->1	o->1	
et.Fr	a->4	u->4	å->4	
et.Fö	l->1	r->13	
et.Ha	n->4	
et.He	l->1	r->22	
et.Hi	t->1	
et.Hu	r->1	v->1	
et.Hä	r->4	
et.I 	F->1	N->1	a->2	b->1	d->8	e->2	f->1	k->1	l->1	o->1	r->2	s->1	ä->1	
et.Ib	l->1	
et.In	g->1	n->1	s->1	
et.Ja	 ->1	g->78	
et.Ju	 ->1	
et.Ko	m->4	n->1	
et.Ku	l->1	
et.Kä	r->1	
et.La	 ->1	
et.Li	k->1	t->1	
et.Lå	t->3	
et.Ma	n->8	
et.Me	d->5	n->23	
et.Mi	n->6	
et.Na	t->1	
et.Ni	 ->4	
et.Nu	 ->4	m->1	v->1	
et.Nä	r->4	s->1	
et.Nö	d->1	
et.Oc	h->7	
et.Om	 ->5	
et.Or	d->1	k->1	
et.Pa	r->3	
et.Po	r->1	
et.Pr	o->2	
et.Pu	n->1	
et.På	 ->5	
et.Ra	p->1	
et.Re	d->1	s->1	
et.Rä	t->1	
et.Sk	o->1	u->1	
et.Sl	u->1	
et.So	c->1	m->3	
et.St	a->2	o->1	
et.Så	 ->7	v->1	
et.Ta	c->3	n->1	
et.Th	e->1	
et.Ti	l->2	
et.Tr	e->1	o->1	
et.Tu	s->1	
et.Ty	 ->1	v->1	
et.Un	i->1	
et.Ur	 ->1	
et.Ut	s->1	
et.Va	d->2	r->2	
et.Vi	 ->47	d->1	s->1	
et.Vä	s->1	
et.Vå	r->2	
et.Än	d->1	
et.Äv	e->1	
et.Å 	e->1	
et.År	 ->1	
et.Åt	e->1	
et.Ös	t->1	
et: "	M->1	
et: F	r->1	
et: J	a->1	
et: U	t->1	
et: d	e->2	
et: e	n->1	
et: f	ö->1	
et: k	a->1	
et: o	m->1	
et: t	a->1	
et: v	å->1	
et: ö	n->1	
et; D	a->1	
et; a	r->1	
et; d	e->1	
et; f	o->1	r->1	
et; u	n->1	
et? R	å->1	
et?. 	(->1	
et?.(	E->1	
et?At	t->1	
et?De	 ->1	t->2	
et?He	r->1	
et?Hu	r->2	
et?I 	v->1	
et?Ja	g->2	
et?Ko	m->1	
et?Kä	r->1	
et?Ni	 ->2	
et?Nä	r->1	
et?Oc	h->1	
et?RI	N->1	
et?Sk	u->1	
et?Va	d->1	
et?Vi	l->1	s->1	
et?Är	 ->1	
etJag	 ->1	
eta -	 ->1	
eta a	l->1	t->9	v->1	
eta b	e->1	i->1	
eta d	e->2	i->1	
eta e	f->2	n->6	t->2	
eta f	a->1	r->3	ö->21	
eta h	i->1	u->1	
eta i	 ->7	n->2	
eta k	l->1	o->1	r->1	
eta m	e->17	
eta n	ä->1	
eta o	c->1	m->6	r->1	
eta p	r->6	å->5	
eta r	e->3	i->1	
eta s	a->1	n->1	
eta t	e->1	i->3	
eta u	p->1	
eta v	a->4	e->1	i->2	
eta å	t->6	
eta ö	v->1	
eta, 	e->1	i->1	r->1	s->1	
eta. 	D->1	
eta.D	e->1	
eta.T	r->1	
eta?V	i->1	
etabl	e->13	
etade	 ->2	
etag 	a->1	b->1	e->2	f->3	h->5	i->6	k->4	l->2	n->1	o->6	p->2	s->18	u->1	v->1	ä->2	
etag,	 ->14	
etag.	A->1	D->4	E->2	F->1	J->1	K->2	M->1	R->1	T->1	V->1	
etaga	n->1	r->22	
etage	n->61	t->5	
etagn	e->8	i->1	
etags	 ->3	a->4	e->5	g->2	i->1	j->2	k->1	l->1	n->1	r->2	s->3	
etakt	.->1	
etala	 ->19	"->1	,->3	.->6	?->2	d->3	r->29	s->3	t->7	
etalj	 ->2	,->2	.->1	a->1	e->26	f->1	k->2	
etall	,->1	d->1	e->8	i->1	
etaln	i->15	
etalt	.->1	s->1	
etand	e->16	
etane	r->5	
etank	e->3	f->2	r->4	
etans	k->5	l->1	
etapp	 ->1	e->4	
etar 	a->1	b->1	e->3	f->4	g->1	i->2	m->4	o->3	p->2	u->1	
etar,	 ->1	
etar.	D->1	
etare	 ->5	,->2	.->2	
etari	a->2	s->1	
etark	l->1	
etarn	a->5	
etas 	ä->1	
etas.	F->1	
etat 	b->2	d->1	e->1	f->2	h->1	i->1	m->2	s->1	u->1	
etats	 ->2	
etbeh	o->1	
etc. 	o->1	Ä->2	
etc.D	e->1	
etc.E	n->1	
etc?A	t->1	
etder	a->1	
ete (	K->2	
ete -	 ->2	,->1	
ete a	n->1	t->1	
ete b	e->1	l->1	ö->1	
ete d	e->1	ä->1	
ete f	ö->9	
ete h	a->5	o->1	
ete i	 ->5	n->4	
ete k	a->2	o->1	r->1	u->1	v->1	
ete l	a->1	e->2	
ete m	e->22	
ete o	c->11	m->3	
ete p	å->6	
ete r	e->1	
ete s	e->1	k->2	o->19	
ete t	i->1	
ete u	p->1	
ete v	i->2	
ete ä	r->1	
ete å	t->1	
ete, 	a->1	d->1	f->1	g->1	l->1	o->2	p->1	s->1	v->2	
ete. 	D->1	
ete..	 ->1	
ete.A	k->1	
ete.D	e->5	
ete.F	r->1	
ete.H	e->1	
ete.I	 ->1	
ete.J	a->3	
ete.K	o->1	
ete.L	i->1	ä->1	å->1	
ete.M	e->2	
ete.N	i->1	
ete.P	å->1	
ete.R	e->1	å->1	
ete.S	o->1	
ete.U	p->1	
ete.V	i->1	å->1	
ete.Å	t->1	
ete?H	u->1	
ete?I	 ->1	
ete?S	o->1	
eteck	e->2	n->10	
eteen	d->3	
eten 	(->1	-->2	1->1	a->47	b->2	d->1	e->4	f->38	g->4	h->11	i->40	j->1	k->8	l->1	m->17	o->40	p->17	r->2	s->22	t->7	u->4	v->10	ä->13	å->2	ö->1	
eten)	 ->1	
eten,	 ->31	
eten.	A->2	D->12	E->2	F->3	H->2	I->1	J->6	K->4	L->1	M->4	N->3	O->3	S->2	V->7	Å->1	
eten:	 ->1	
etena	 ->3	
etenh	e->1	
etens	 ->35	,->3	.->2	k->71	
etent	 ->2	a->2	
eter 	-->3	E->1	O->1	a->20	b->2	d->3	e->3	f->21	g->3	h->6	i->22	k->5	l->3	m->9	o->54	p->8	r->3	s->37	t->12	u->5	v->2	ä->10	å->1	ö->2	
eter,	 ->31	
eter.	 ->2	A->1	D->14	E->5	F->1	J->4	K->2	M->2	O->1	S->1	T->2	V->3	Ä->1	
eter?	D->1	
etera	n->9	r->2	
eteri	n->4	
eterl	i->1	
etern	 ->1	a->120	
eters	 ->3	e->1	
etess	 ->4	b->5	e->2	h->1	
etet 	a->3	f->5	h->3	i->5	k->2	m->11	o->9	p->4	s->2	t->1	u->1	v->1	ä->2	
etet"	.->1	
etet,	 ->3	
etet.	D->2	H->1	I->1	J->1	K->1	R->1	T->1	
etete	n->1	
etets	 ->1	
etfrå	g->2	
etför	f->2	o->6	s->1	
eth S	c->1	
etik 	o->2	
eting	e->2	
etise	r->2	
etisk	.->1	a->3	t->3	
etiti	o->1	
etjän	t->1	
etkon	t->16	
etkra	v->1	
etlig	 ->15	.->2	?->1	a->7	h->3	t->8	
etmat	c->1	
etmäs	s->1	
etna 	b->1	o->16	
etnis	k->14	
etod 	a->1	b->1	f->2	m->2	s->5	ä->1	å->1	
etode	n->4	r->12	
etona	 ->26	d->6	r->7	s->1	t->5	
etoni	n->1	
etori	k->3	
etpla	n->3	
etpol	i->1	
etpos	t->10	
etrak	t->23	
etran	s->1	
etrar	n->1	
etroa	k->12	
etrol	e->1	
etrus	t->1	
etryc	k->3	
etryg	g->1	
eträd	a->59	d->3	e->9	s->2	
eträf	f->79	
eträt	t->1	
ets "	g->1	
ets -	 ->1	
ets B	a->1	
ets L	e->1	
ets a	b->1	l->1	m->2	n->4	r->6	u->1	
ets b	e->25	i->2	u->1	
ets c	e->1	
ets d	e->8	i->11	o->2	
ets e	f->2	g->2	
ets f	a->2	e->1	i->1	j->1	o->1	r->4	u->2	ö->28	
ets g	e->13	i->3	r->14	å->1	
ets h	a->1	i->2	j->1	u->1	ä->2	å->1	
ets i	k->1	n->2	
ets k	l->1	o->2	r->2	u->1	ä->1	
ets l	a->2	e->6	i->1	o->2	ö->1	
ets m	a->1	e->4	i->2	o->2	y->1	å->1	ö->5	
ets n	e->1	u->1	y->2	
ets o	c->21	h->1	i->1	r->17	t->1	
ets p	a->1	e->2	l->1	o->4	r->4	u->1	
ets r	e->13	i->2	ä->5	
ets s	a->1	e->2	i->5	k->3	l->5	o->1	p->1	t->13	u->1	y->4	ä->1	
ets t	a->3	e->1	i->4	j->1	r->3	
ets u	p->3	t->6	
ets v	e->2	ä->2	
ets y	t->3	
ets ä	n->2	
ets å	l->1	s->1	
ets ö	n->1	v->1	
ets, 	S->1	f->1	
ets- 	o->5	
ets.E	n->1	
etsak	t->1	
etsam	m->6	
etsan	d->5	
etsar	 ->2	.->1	b->1	g->1	
etsas	p->3	
etsav	b->1	t->1	
etsba	s->1	
etsbe	s->5	
etsbu	d->1	
etsbö	r->5	
etsce	r->1	
etsch	e->3	
etsdo	k->4	
etsen	 ->3	h->3	
etsfi	e->1	
etsfl	a->15	
etsfo	r->1	
etsfr	å->9	
etsfå	n->1	
etsfö	r->4	
etsga	r->3	
etsgi	v->8	
etsgr	e->2	u->5	ä->1	
etsha	n->2	
etsin	s->2	
etsit	u->1	
etska	m->1	p->1	
etskl	a->1	i->1	
etsko	e->1	n->2	
etskr	a->5	i->3	
etsla	g->3	
etsli	v->2	
etslo	p->2	
etslä	n->1	
etslö	s->43	
etsma	n->1	r->12	
etsme	t->2	
etsmy	n->8	
etsmä	n->2	
etsni	v->2	
etsno	r->6	
etsnä	t->1	
etsom	r->5	
etsor	d->10	g->1	
etspa	k->4	
etspe	r->2	
etspl	a->9	
etspo	l->6	
etspr	i->70	o->6	
etsra	m->1	p->2	
etsre	g->3	
etsri	s->1	
etsru	m->1	t->1	
etsrä	t->3	
etsrå	d->18	
etssa	n->1	
etssi	f->2	
etssk	ä->2	
etssp	r->1	
etsst	a->1	y->2	
etssy	n->1	s->2	
etsta	g->40	
etsti	d->10	l->38	
etstä	n->2	
etstö	d->2	
etsut	b->5	
etsva	n->1	
etsve	n->1	
etsvi	l->5	
etsyn	p->1	
etsåt	g->2	
ett "	o->1	
ett 5	0->1	
ett A	m->1	
ett E	G->1	u->14	
ett a	b->1	d->3	k->3	l->15	m->2	n->52	r->4	t->17	v->31	
ett b	a->1	e->37	i->3	l->1	r->31	u->1	y->1	ä->11	ö->1	
ett c	e->3	i->1	
ett d	a->2	e->12	i->19	j->3	o->9	r->1	u->1	
ett e	-->1	f->14	g->2	k->3	l->2	m->1	n->26	r->2	t->3	u->9	v->2	x->15	
ett f	a->11	e->1	i->1	l->13	o->8	r->16	u->7	å->1	ö->67	
ett g	a->2	e->21	i->1	o->14	r->2	
ett h	a->5	e->3	i->4	j->1	o->4	u->5	y->1	å->7	ö->5	
ett i	 ->4	c->1	f->1	m->1	n->43	r->3	t->1	
ett j	a->2	u->3	ä->3	
ett k	a->3	l->8	o->23	r->6	u->2	v->4	ä->2	
ett l	a->20	e->3	i->5	j->1	o->1	u->1	y->1	ä->4	å->2	ö->2	
ett m	a->4	e->27	i->18	o->5	u->2	y->40	ä->1	å->13	ö->3	
ett n	a->3	e->3	u->1	y->20	ä->3	å->1	ö->3	
ett o	a->1	b->2	c->4	d->1	e->2	f->4	g->1	l->2	m->36	n->1	p->3	r->13	s->3	ä->1	ö->1	
ett p	a->27	e->6	i->1	o->20	r->29	å->6	
ett r	a->1	e->24	i->6	u->1	y->1	ä->6	å->1	ö->1	
ett s	.->1	a->15	e->6	i->5	j->6	k->6	l->11	n->1	o->5	p->3	t->54	u->1	v->7	y->18	ä->22	å->45	
ett t	a->7	e->2	i->25	o->3	r->9	y->8	å->1	
ett u	l->1	n->5	p->5	r->5	t->33	
ett v	a->3	e->7	i->27	r->1	ä->9	
ett w	o->1	
ett y	p->1	t->4	
ett ä	n->12	r->8	
ett å	l->1	r->16	t->6	
ett ö	k->2	m->1	p->4	v->9	
ett, 	f->1	i->1	k->1	o->1	t->2	u->1	
ett. 	I->1	
ett..	(->1	
ett.D	e->2	
ett.F	ö->1	
ett.H	e->1	
ett.J	a->1	
ett.M	e->1	o->1	
ett.Ä	v->1	
ett: 	H->1	s->1	
etta 	-->6	A->1	E->6	F->1	a->23	b->66	c->2	d->40	e->12	f->75	g->10	h->31	i->45	k->37	l->13	m->52	n->8	o->59	p->75	r->8	s->119	t->18	u->20	v->28	y->2	ä->159	å->6	ö->3	
etta!	F->1	
etta,	 ->39	
etta.	 ->1	(->1	.->1	A->1	B->1	C->1	D->19	E->5	F->1	G->1	H->2	I->6	J->7	K->1	M->6	N->1	O->3	P->1	S->4	T->1	V->9	Ä->1	
etta:	 ->1	
etta?	J->1	
ette 	d->1	
ette-	L->1	
etter	a->13	i->5	
ettet	,->1	
ettic	h->1	
ettid	e->1	
ettig	 ->1	a->1	t->1	
ettio	f->1	t->1	
etton	 ->3	s->1	
etts 	a->2	f->1	g->1	i->2	m->1	o->1	u->2	ö->1	
etts,	 ->1	
etts.	D->1	E->1	I->1	
ettvi	l->1	
etung	a->1	
etuts	k->10	
etvis	 ->25	,->1	.->1	
etviv	l->3	
ety ä	r->1	
ety-p	r->1	
etyda	 ->1	n->16	
etydd	e->1	
etyde	l->73	r->18	
etydi	g->7	
etydl	i->13	
etänk	a->287	e->1	l->5	
etära	 ->6	
etåre	t->10	
etête	 ->2	
etöve	r->1	
eugen	 ->1	.->1	
eum v	ä->1	
eundr	a->3	
euro 	1->1	b->1	f->6	h->1	i->1	o->1	p->3	t->1	u->1	
euro!	A->1	
euro,	 ->6	
euro.	D->3	H->1	K->1	N->1	S->1	V->1	
eurof	e->1	
euron	 ->3	,->1	s->2	
euroo	m->1	
europ	a->9	e->355	r->1	é->10	
euros	k->2	
eussa	g->1	
eutbi	l->1	
eutiq	u->1	
eutra	l->2	
eutro	t->1	
eutsc	h->1	
eutsl	ä->2	
eutve	c->4	
ev an	s->1	
ev av	 ->1	s->1	
ev di	r->1	
ev dj	u->1	
ev dä	r->2	
ev fa	l->1	
ev fr	å->1	
ev fö	r->1	
ev in	 ->1	t->1	v->1	
ev kv	a->1	
ev ny	l->1	
ev ob	e->1	l->1	
ev oc	k->1	
ev om	 ->1	
ev so	m->1	
ev ti	l->2	
ev tv	u->1	
ev un	d->1	i->1	
ev.Fr	u->1	
eva d	ä->1	
eva e	n->1	t->1	
eva f	l->1	
eva h	u->1	
eva i	 ->4	
eva l	i->1	
eva m	e->2	
eva n	å->1	
eva p	å->1	
eva s	j->1	
eva u	p->1	
eva v	å->1	
eva, 	u->1	
eva?N	e->1	
evaka	 ->2	r->1	
evakn	i->3	
evald	 ->4	a->2	
evand	e->3	
evant	 ->3	a->6	
evara	 ->13	n->8	t->1	
evatt	n->2	
evde 	d->1	g->1	
evebr	ö->1	
eveka	 ->1	
evel 	s->1	
evels	e->1	
evene	m->1	
event	u->20	
ever 	a->3	e->1	f->1	i->1	j->1	l->1	m->1	u->3	
ever.	K->1	
evera	n->3	
evere	r->4	
evide	r->18	
evig 	v->1	
evigt	 ->1	.->1	
evilj	a->48	
evis 	-->1	a->1	e->1	f->3	i->2	l->1	m->1	o->2	p->7	s->4	t->1	ä->2	
evis,	 ->1	
evis.	D->1	H->1	
evisa	 ->3	d->2	s->1	
evisb	ö->7	
evise	n->2	t->3	
evisi	o->22	
evisn	i->1	
evitt	n->1	
evlig	 ->2	t->1	
evlåd	e->1	
evnad	 ->2	,->2	.->1	?->1	s->6	
evolu	t->1	
evs a	v->1	
evs o	c->1	
evs s	o->3	
evs u	t->1	
evt d	e->1	
evt e	n->1	t->1	
evt i	 ->1	
eväck	a->3	
evärd	 ->4	a->4	
evärt	 ->3	,->1	.->2	
evåna	r->2	
ew Yo	r->1	
ewies	 ->1	
ewood	 ->1	s->1	
ex al	l->1	
ex an	t->4	
ex av	 ->1	
ex eu	r->1	
ex fl	e->1	
ex mi	n->1	
ex må	n->10	
ex pl	a->1	
ex po	s->1	
ex ti	l->1	
ex tu	n->1	
ex öv	e->1	
ex, s	j->1	
ex. E	u->1	
ex. F	r->1	
ex. N	e->1	
ex. U	S->1	
ex. a	t->1	v->1	
ex. d	e->2	
ex. e	t->1	
ex. i	n->1	
ex. k	u->1	ä->1	
ex. m	i->2	
ex. n	ä->2	
ex. o	l->1	
ex. p	å->1	
ex. u	t->1	
ex. v	a->1	
ex.Ja	g->1	
exa, 	t->1	
exakt	 ->10	,->1	a->6	h->1	
exame	n->6	
exami	n->10	
exand	e->2	
exas 	g->1	i->1	
excep	t->5	
exemp	e->109	l->8	
exibe	l->11	
exibi	l->10	
exibl	a->6	
exiko	,->1	
exilr	e->1	
exilt	i->1	
exism	e->1	
exist	e->19	
exklu	s->3	
exmån	a->1	
expan	d->5	s->1	
exped	i->1	
exper	t->44	
expli	c->1	
explo	s->2	
expon	e->2	
expor	t->4	
ext a	v->1	
ext f	å->1	
ext i	 ->1	
ext k	o->1	
ext l	i->1	
ext o	c->2	m->1	
ext s	k->1	o->4	
ext, 	o->1	s->3	ä->1	
ext.M	e->1	
exten	 ->11	"->2	,->2	.->2	
exter	 ->2	,->2	.->2	n->11	
exton	.->1	
extra	 ->5	o->1	
extre	m->30	
exuel	l->3	
exvär	t->1	
ey Ca	n->3	
eyer 	h->1	n->1	
eyer.	O->1	
eyhun	 ->1	
ez Go	n->1	
ez an	g->1	
ez oc	h->1	
ez to	g->1	
ez, i	n->1	
ez, u	t->1	
ez-ka	t->2	
ezuel	a->1	
eägar	e->2	
eåter	f->1	
f - a	t->1	
f Hit	l->2	
f av 	d->1	
f ell	e->1	
f ext	r->1	
f för	 ->4	e->1	
f had	e->1	
f har	 ->2	
f i f	ä->1	
f inn	a->1	
f int	r->1	
f kun	n->1	
f lik	s->1	
f nol	l->1	
f och	 ->3	
f ock	s->1	
f om 	f->1	
f som	 ->4	
f the	 ->1	
f uta	n->1	
f ägt	 ->1	
f, ha	d->1	
f, me	n->1	
f, oc	h->1	
f, på	 ->1	
f, so	m->1	
f- oc	h->2	
f-Mat	h->2	
f.Det	 ->1	
f.Där	f->1	
f.End	a->1	
f.Jag	 ->1	
f.d. 	Ö->1	ö->1	
fa al	l->2	
fa ar	b->1	
fa bu	d->1	
fa de	n->2	
fa ek	o->2	
fa en	 ->3	
fa fo	t->1	
fa fr	a->1	
fa fö	r->1	
fa in	o->1	
fa ko	m->1	n->2	
fa mi	s->1	
fa oc	h->1	
fa re	a->1	
fa si	g->2	
fa un	i->1	
fa ut	a->1	
fa, o	c->1	
fa, å	t->1	
fa.Me	n->1	
fabet	e->1	
fabri	k->1	
fackf	ö->4	
fadde	r->1	
fade 	2->1	i->1	j->1	k->1	n->1	s->1	t->1	
fader	,->1	
fades	 ->1	.->1	
fael 	-->1	l->1	
fael.	N->1	
failu	r->1	
fakta	 ->6	.->1	i->2	
fakti	s->49	
fakto	r->14	
faktu	m->64	
fala 	f->1	
fald 	i->2	ä->1	
fald,	 ->5	
falde	n->5	
faldi	g->2	
fall 	K->1	a->6	b->5	d->4	e->5	f->10	g->3	h->4	i->4	j->2	k->8	l->1	m->4	o->4	p->1	r->1	s->16	t->2	u->3	v->1	ä->5	ö->1	
fall,	 ->11	
fall.	 ->2	B->1	D->4	E->1	H->1	J->3	M->1	S->1	V->2	
falla	s->1	
falle	n->8	r->36	t->56	
falli	t->4	
falls	f->1	h->1	m->1	s->3	t->1	ä->1	
falsk	a->2	n->1	t->1	
famil	j->15	
fande	 ->41	t->1	
fann 	d->1	t->1	
fanns	 ->14	
fant 	i->1	
fanta	s->11	
fantl	i->2	
far E	v->1	
far L	y->1	
far S	w->1	
far a	r->1	s->1	
far b	a->1	ö->1	
far d	e->9	
far e	n->2	
far h	a->1	u->1	
far i	 ->1	a->1	g->1	
far k	a->1	o->1	
far l	i->1	
far m	y->1	
far o	c->1	
far p	u->1	
far s	a->1	t->1	ä->1	å->1	
far u	n->1	
far ä	r->1	
far ö	v->1	
far, 	a->1	m->1	o->1	u->1	
far. 	E->1	
far.D	e->3	å->1	
far.I	 ->1	
far.J	a->2	
far.V	i->1	
far: 	v->1	
far?K	a->1	
fara 	e->1	f->4	r->1	t->2	y->1	
fara,	 ->2	
fara.	A->1	
faran	 ->2	d->165	
farar	 ->3	
fare 	n->1	
faren	 ->1	h->24	
farhå	g->2	
farit	 ->2	
farli	g->59	
farma	k->1	
farna	 ->1	
faror	 ->3	.->1	
farso	t->1	
fart 	p->1	
fart,	 ->1	
fart.	V->1	
farte	n->2	
farts	i->1	m->1	o->2	s->3	
farty	g->69	
farva	t->9	
fas h	å->1	
fas o	l->1	
fas t	y->1	
fas v	i->1	
fas, 	a->1	d->1	
fas.D	å->1	
fasci	s->11	
fasen	 ->2	,->1	.->1	
fasni	n->3	
fasor	,->1	
fast 	a->4	d->1	f->1	i->4	m->1	n->2	t->1	v->9	ö->1	
fast.	K->1	N->1	
fasta	 ->5	
fasti	g->1	
fastk	u->1	
fastl	a->3	ä->2	
fastn	a->1	
fasts	l->21	t->51	
fastä	n->1	
fat e	n->1	
fat g	e->1	
fat i	 ->1	
fat p	å->1	
fat s	j->1	
fat.D	e->2	ä->1	
fat.V	a->1	
fats 	e->1	h->1	
fatta	 ->37	.->1	d->7	n->40	r->40	s->29	t->18	
fatti	g->30	
fattn	i->55	
fauna	 ->1	
favor	i->1	
faxa 	e->1	
fbest	ä->1	
fdrab	b->1	
febru	a->16	
feder	a->12	
fekt 	i->1	k->1	m->2	p->1	s->1	u->1	
fekt.	I->1	M->1	
fekta	 ->1	
fekte	n->12	r->25	
fekti	o->1	v->114	
fel a	t->2	v->2	
fel o	c->3	
fel s	i->1	o->1	ä->1	
fel u	p->1	
fel! 	I->1	
fel, 	m->1	o->2	s->1	
fel.D	e->2	
fel.G	e->1	
fel.J	a->1	
felak	t->12	
felan	d->1	
felba	r->1	
felbe	r->1	
felen	,->1	
felkv	o->1	
felrä	k->1	
felsy	n->1	
fem a	l->1	n->1	v->1	
fem d	a->1	
fem g	å->1	
fem k	o->2	
fem m	å->1	
fem p	u->2	
fem v	e->1	i->1	
fem å	r->14	t->1	
fem, 	s->1	
fem: 	p->1	
fempu	n->1	
femte	 ->14	d->2	
femti	e->1	o->2	
femto	n->5	
femår	i->1	s->2	
fen D	u->1	
fen S	S->1	
fen d	å->1	
fen g	e->1	
fen i	 ->1	
fen l	o->1	
fen m	e->3	å->1	
fen o	c->2	
fen u	t->2	
fen v	a->1	
fen ä	r->2	
fen, 	d->1	e->1	n->1	o->1	s->1	
fen-S	S->1	
fen.D	e->1	
fen.F	o->1	
fen.I	 ->1	
fen.Ä	r->1	
fenom	e->3	
fens 	o->1	
fensi	v->3	
fentl	i->80	
fer a	v->1	
fer e	l->1	
fer f	ö->7	
fer h	a->1	ä->1	
fer i	 ->3	n->3	
fer m	e->1	å->1	
fer o	c->3	
fer p	å->2	
fer s	k->1	o->3	
fer u	t->1	
fer ä	r->1	
fer" 	m->1	
fer, 	d->1	h->1	k->1	o->5	s->2	
fer.D	e->2	
fer.N	a->1	
fer.O	m->1	
fer.V	i->2	
fera 	l->2	r->1	
fera.	J->1	
feren	s->174	t->5	
ferer	a->3	
ferie	n->1	
ferin	.->1	
ferna	 ->8	,->2	s->2	
fert.	J->1	
ferta	r->1	
fessi	o->2	
fesso	r->6	
festa	t->1	
fety-	p->1	
ff no	l->1	
ff oc	h->2	
ff, p	å->1	
ff- o	c->2	
ffa a	l->2	r->1	
ffa b	u->1	
ffa d	e->2	
ffa e	k->2	n->3	
ffa f	o->1	r->1	ö->1	
ffa i	n->1	
ffa k	o->3	
ffa m	i->1	
ffa o	c->1	
ffa r	e->1	
ffa s	i->2	
ffa u	n->1	t->1	
ffa, 	o->1	å->1	
ffa.M	e->1	
ffade	 ->7	s->2	
ffand	e->42	
ffar 	E->1	L->1	S->1	a->1	b->2	d->9	e->2	h->2	i->3	k->2	l->1	m->1	o->1	p->1	s->4	u->1	ä->1	ö->1	
ffar,	 ->4	
ffar.	 ->1	D->4	I->1	J->2	V->1	
ffar:	 ->1	
ffar?	K->1	
ffare	 ->1	
ffas 	h->1	o->1	t->1	v->1	
ffas.	D->1	
ffat 	e->1	g->1	i->1	p->1	s->1	
ffat.	D->3	V->1	
ffats	 ->1	
ffbes	t->1	
ffekt	 ->2	.->1	e->36	i->114	
ffen 	S->1	
ffen-	S->1	
ffens	 ->1	i->3	
ffent	l->80	
ffer 	f->7	i->1	s->1	
ffer,	 ->3	
ffere	n->5	
ffert	a->1	
ffice	 ->1	
ffici	e->6	
fflag	s->1	
fflig	a->1	h->1	
ffpro	c->2	
ffra 	e->1	f->1	s->1	ä->1	
ffra,	 ->3	
ffrad	e->1	
ffrar	 ->1	
ffren	 ->11	,->1	s->2	
ffror	 ->6	.->2	?->1	n->6	
ffrät	t->28	
ffäre	n->3	r->8	
ffärs	m->1	
fhjäl	p->1	
fi oc	h->1	
fi på	 ->1	
fi so	m->1	
fi, m	e->1	
fi.De	t->1	
fi.Vi	 ->1	
fice 	n->1	
ficer	a->29	i->9	
ficie	l->7	n->1	
fick 	K->1	d->1	e->3	h->2	i->4	j->3	m->2	n->2	o->2	s->2	u->1	v->3	
ficko	r->1	
fiden	t->2	
fiend	e->1	
fient	l->33	
fiera	 ->7	d->7	s->3	t->5	
fierb	a->2	
fieri	n->3	
fik o	c->1	
fik s	t->1	å->1	
fik ä	r->1	
fik å	t->1	
fik- 	o->1	
fik.B	y->1	
fik.D	e->1	
fika 	b->1	f->5	k->2	l->1	p->2	r->3	t->1	u->1	å->1	
fikat	 ->4	i->1	
fiken	 ->2	.->1	
fikle	d->1	
fikt 	d->1	f->1	g->1	h->1	k->1	v->1	ä->1	
fil u	t->1	
fil.D	e->1	
fil.L	y->1	
filme	n->1	r->1	
filos	o->5	
filsk	a->1	
filtr	e->1	
fin i	 ->1	
fin s	å->1	
fin-r	å->3	
fin.V	i->1	
fina 	b->1	s->1	
finan	s->81	
fing-	P->1	
finge	r->1	
finie	r->13	
finin	g->1	
finit	i->23	u->1	
finlä	n->5	
finna	 ->21	s->39	
finne	r->39	
finns	 ->309	,->3	.->5	
finsk	 ->1	a->5	
fintl	i->10	
fique	s->1	
fira 	m->1	
firar	e->1	n->1	
fisk 	o->2	u->1	
fiska	 ->7	d->1	r->4	s->1	
fiskb	e->4	
fiske	 ->4	)->2	,->4	.->2	k->1	m->4	o->2	r->9	s->1	t->8	v->2	
fiskt	 ->2	
fit-a	n->5	
fjol 	o->2	
fjol,	 ->1	
fjol.	K->1	
fjort	o->9	
fjärd	e->11	
fkrig	e->1	
flagg	 ->6	,->7	.->5	;->1	a->5	e->2	n->1	o->1	
flagr	a->1	
flags	t->1	
flams	k->4	
flekt	e->3	i->4	
fler 	a->2	b->2	d->1	f->1	i->1	k->3	l->2	m->3	n->1	p->3	s->2	t->2	ä->1	
fler,	 ->1	
flera	 ->56	
flers	t->1	
flert	a->5	
flerå	r->12	
flest	a->25	
flexi	b->27	
flick	o->1	
fliga	 ->1	
fligh	e->1	
flikt	 ->4	e->11	f->1	
flirt	a->1	
flit 	p->1	
flite	n->1	
flod 	t->2	
flode	n->2	
flora	 ->1	
flott	a->3	o->1	
flute	t->1	
flutn	a->13	
flyg,	 ->1	
flyga	 ->1	n->1	
flygb	l->1	
flyge	r->1	t->1	
flygk	r->1	
flygn	i->1	
flygp	l->4	
flygt	r->2	
flykt	e->3	i->13	
flyr 	f->1	
flyta	n->12	
flyte	l->1	
flytt	 ->1	.->1	a->11	n->4	
fläck	a->1	
fläkt	a->1	
flöde	n->1	t->2	
flödi	g->1	
fmann	 ->1	
fobin	,->1	
foder	 ->2	,->2	.->4	m->1	t->1	
fog f	ö->1	
foga 	a->4	f->1	ö->1	
fogad	.->1	e->2	
fogan	d->11	
fogar	 ->7	
fogat	 ->3	
fogen	h->27	
fokus	 ->1	.->1	e->3	
folk 	a->1	b->2	h->1	i->2	o->2	s->2	u->1	
folk,	 ->1	
folk.	A->1	D->1	M->1	O->1	V->4	
folka	d->1	
folke	n->6	t->14	
folkg	r->2	
folkh	ä->9	
folkl	i->1	
folkn	i->43	
folko	m->6	
folkp	a->10	
folkr	e->2	ä->1	
folks	 ->3	t->1	ä->1	
folkv	a->2	
fon, 	5->1	
fond 	f->4	k->1	s->2	
fonde	n->43	r->69	
fondm	e->3	
fonds	p->3	
fondu	p->1	
fone-	M->1	
for o	c->1	
for s	o->1	
fora 	p->1	
force	 ->1	
ford-	f->1	
forde	r->5	
fordo	n->65	
fordr	a->17	i->1	
form 	a->26	b->1	d->1	e->1	f->1	i->3	j->1	k->2	l->1	o->2	p->1	s->6	v->2	ä->1	
form,	 ->8	
form.	D->1	E->1	M->1	N->1	S->1	V->1	Ä->1	
form:	 ->1	
forma	 ->7	d->1	n->4	r->3	s->3	t->75	
forme	l->16	n->15	r->98	
formf	ö->2	
formi	s->1	
formn	i->26	
formp	a->1	r->14	
forms	t->1	
formu	l->18	
formå	t->1	
fors 	b->2	e->1	f->3	g->1	h->3	i->4	k->2	o->3	s->2	t->2	u->1	
fors,	 ->7	
fors.	D->5	J->1	M->1	T->1	U->1	V->1	
forsb	e->1	
forsk	a->5	n->34	
fort 	h->1	s->2	
fortb	i->1	
fortf	a->89	
fortg	å->5	
fortl	e->1	
forts	a->12	k->1	ä->82	
forum	 ->4	e->1	
forêt	s->1	
fossi	l->3	
foste	r->1	
fotbo	l->1	
fotfä	s->1	
fotsp	å->2	
fproc	e->2	
fra e	n->1	
fra f	ö->1	
fra s	o->1	
fra ä	r->1	
fra, 	1->1	h->1	m->1	
frade	s->1	
frakt	a->10	f->1	
fram 	8->1	a->6	b->2	d->19	e->55	f->15	g->1	h->3	i->8	k->3	l->2	m->3	n->3	o->7	p->3	r->5	s->12	t->45	u->2	v->4	ä->4	å->1	ö->1	
fram,	 ->8	
fram.	.->1	D->1	F->2	H->1	K->1	R->1	
framf	a->1	ö->142	
framg	i->1	å->52	
framh	ä->5	å->17	ö->2	
framk	a->1	o->10	
framl	a->13	ä->7	
framm	e->1	
frams	k->2	t->46	
framt	 ->1	a->4	i->106	r->2	v->2	
framå	t->21	
framö	v->2	
franc	,->1	a->1	
frans	k->33	m->3	
frar 	y->1	
frase	r->1	
frast	r->15	
fred 	i->6	m->1	o->7	v->1	
fred,	 ->1	
fred.	D->1	H->2	I->1	
frede	n->2	
fredl	i->8	
freds	 ->1	,->1	.->1	a->4	b->2	f->3	p->22	s->28	u->1	
free-	f->1	l->1	
free.	D->1	
frekv	e->1	
fren 	f->9	o->1	v->1	
fren,	 ->1	
frens	 ->2	
frest	a->1	e->3	n->1	
fri f	r->1	ö->1	
fri i	n->2	
fri k	o->2	
fri r	ö->8	
fri ö	p->1	
fri, 	o->1	
fri- 	o->8	
fria 	P->1	a->2	d->1	f->1	i->1	m->1	o->1	r->10	s->1	t->1	v->4	å->1	
fria,	 ->2	
frias	 ->3	
friat	 ->1	
friel	s->6	
frigj	o->1	
frigö	r->5	
friha	n->2	
frihe	t->113	
frika	 ->3	.->3	
frikt	i->1	
frisl	ä->2	
frist	 ->4	e->7	i->1	ä->1	å->1	
fritt	 ->3	,->1	.->1	
frivi	l->12	
froda	s->4	
front	a->1	e->3	
fror 	f->1	p->2	s->1	u->1	ö->1	
fror.	J->1	V->1	
fror?	H->1	
frorn	a->6	
fru A	h->1	n->1	
fru F	r->1	
fru P	e->1	
fru R	e->3	
fru S	c->2	u->1	
fru T	h->1	
fru W	a->1	
fru k	o->42	
fru t	a->13	
fru, 	s->1	
frukt	 ->1	.->1	a->11	b->2	e->1	
frust	r->2	
fruta	l->1	
frysa	 ->2	
frysn	i->1	
frytt	e->2	
fräck	h->1	
främj	a->61	
främl	i->34	
främm	a->2	
främs	t->47	
frätt	 ->6	,->2	?->1	e->4	s->15	
fråga	 ->211	!->1	,->24	.->40	:->7	?->1	d->8	n->187	r->20	s->20	t->5	v->1	
fråge	k->1	s->8	t->2	
frågn	i->8	
frågo	r->272	
från 	(->21	-->1	1->7	2->1	3->1	5->3	8->1	9->1	A->10	B->5	C->3	D->2	E->29	F->6	G->4	H->2	I->5	J->1	K->5	L->3	M->1	N->3	O->1	P->7	R->1	S->6	T->6	U->2	V->1	W->2	a->35	b->13	d->94	e->43	f->30	g->4	h->6	i->1	j->4	k->36	l->8	m->21	n->6	o->21	p->18	r->17	s->25	t->25	u->22	v->19	Ö->1	ä->1	å->1	ö->4	
från,	 ->3	
från.	D->1	Ä->1	
frång	å->1	
frånk	o->3	
frånt	a->2	o->1	
frånv	a->8	ä->1	
fsitu	a->1	
fstra	t->1	
fströ	m->3	
fstöd	 ->1	.->1	
ft 20	0->1	
ft al	l->1	
ft at	t->4	
ft av	 ->4	
ft be	h->1	t->1	
ft de	n->3	t->1	
ft dä	r->1	
ft en	 ->1	
ft er	s->1	
ft et	t->2	
ft ex	 ->1	
ft fa	l->1	
ft fl	e->1	
ft fr	a->2	å->2	
ft fö	r->8	
ft ge	r->1	
ft ha	r->1	
ft i 	I->1	a->1	l->1	m->1	å->1	
ft in	o->1	
ft ka	n->1	
ft ko	m->1	
ft la	w->1	
ft me	d->2	n->1	
ft my	c->1	
ft må	n->1	
ft mö	j->1	
ft nä	r->2	
ft nå	g->2	
ft oc	h->4	
ft om	 ->2	
ft pr	o->2	
ft på	 ->3	
ft re	d->1	
ft sa	m->1	
ft se	x->1	
ft si	n->1	
ft sk	a->2	u->1	
ft so	m->6	
ft st	o->1	ä->1	ö->1	
ft sv	å->1	
ft så	 ->1	d->1	
ft ta	r->1	
ft ti	l->4	
ft un	d->1	
ft ut	g->1	
ft vi	 ->2	
ft vä	g->1	
ft vå	r->1	
ft är	 ->3	a->1	
ft!He	r->1	
ft, S	c->1	
ft, f	ö->1	
ft, i	n->1	
ft, m	e->2	å->1	
ft, o	c->2	
ft, s	k->1	o->1	
ft, u	t->1	
ft, v	a->1	i->1	
ft. D	e->1	
ft.At	t->1	
ft.De	 ->1	t->1	
ft.Dä	r->1	
ft.Ef	t->1	
ft.He	r->1	
ft.Ja	g->1	
ft.Me	r->1	
ft.Om	 ->1	
ft.Vi	 ->3	d->1	
ft: d	e->1	
ft? M	e->1	
ft?Ne	j->1	
fta a	n->2	t->6	
fta b	e->1	i->1	l->1	o->1	r->1	
fta d	e->3	
fta e	n->1	
fta f	r->4	u->1	ö->3	
fta g	ö->2	
fta h	a->6	u->1	
fta i	 ->1	n->2	
fta k	a->1	
fta l	a->1	i->1	
fta m	o->1	
fta n	o->1	ä->1	
fta o	c->2	g->1	r->2	
fta p	å->2	
fta s	a->2	e->1	k->1	t->1	y->1	ä->1	å->1	
fta t	i->1	v->1	
fta u	n->1	t->2	
fta v	a->1	å->1	
fta ä	r->5	
fta, 	l->1	
fta.O	c->1	
ftade	 ->5	s->1	
ftan 	i->1	m->1	
ftand	e->5	
ftar 	a->2	b->1	d->2	f->1	i->1	j->1	m->1	n->1	o->2	s->1	t->24	
ftare	 ->3	
ftarl	ø->2	
ftarn	a->2	
ftas 	a->2	i->5	
ftas.	J->1	
ftast	 ->1	
ftat 	a->3	m->1	o->1	p->1	
ftats	 ->2	
ftbur	e->1	
fte a	t->9	
fte d	e->1	
fte g	å->1	
fte i	n->1	
fte m	e->1	
fte o	c->1	
fte s	k->1	o->1	
fte u	t->1	
fte v	a->1	
fte ä	n->1	r->1	
fte, 	o->1	
fte.D	e->1	
fte.V	a->1	
ftels	e->1	
ften 	a->5	b->1	f->3	i->4	m->3	o->5	p->1	s->4	v->2	ä->2	å->2	
ften,	 ->2	
ften.	D->4	E->1	V->2	
ftena	 ->1	
fter 	-->2	1->1	A->2	E->3	H->1	L->1	M->2	O->1	S->1	T->1	a->38	b->5	d->33	e->15	f->8	g->2	h->8	i->6	j->4	k->4	l->1	m->4	n->2	o->13	p->5	r->3	s->15	t->3	u->2	v->8	ä->3	å->5	ö->1	
fter,	 ->9	
fter.	D->2	F->1	H->1	I->1	J->2	L->1	V->1	
fter:	 ->1	
fter;	 ->1	
fterb	i->1	
fterf	r->8	ö->3	
fterg	i->8	
fterh	a->5	
fterl	e->3	y->2	ä->1	
fterm	i->9	
ftern	a->21	
fters	a->3	o->190	t->12	
ftert	a->3	r->2	ä->1	
fterå	t->1	
ftet 	a->5	b->2	f->1	h->1	m->13	o->1	ä->2	
ftet.	F->1	
ftful	l->12	
ftig 	e->1	g->1	l->1	m->1	o->3	p->1	r->1	u->1	å->1	ö->1	
ftig,	 ->1	
ftiga	 ->15	.->1	r->4	
ftigt	 ->11	,->2	.->3	
ftlig	 ->1	a->1	e->3	t->3	
ftnin	g->113	
ftomr	å->1	
ftone	n->1	
ftor,	 ->1	
ftorn	a->2	
fts- 	o->1	
ftsan	l->4	
ftsfö	r->2	
ftslä	m->2	
ftsmå	l->1	
ftsol	y->1	
ftspl	a->1	
ftspo	l->1	
ftspr	i->1	o->1	
ftsre	a->1	
ftsse	k->1	
ftssä	k->1	
ftsta	k->1	
ftsve	r->1	
ftsäk	e->1	
fttag	.->1	
ftträ	d->4	
ftver	k->8	
full 	a->2	e->1	g->3	h->2	n->1	o->1	p->1	r->2	s->1	ö->1	
full.	D->2	O->1	
fulla	 ->19	,->1	.->2	r->1	s->1	
fullb	o->3	
fullf	ö->3	
fullg	j->1	ö->1	
fullh	e->1	
fullk	o->5	
fullo	 ->5	
fulls	t->41	
fullt	 ->40	,->1	.->2	
fullv	ä->2	
fullä	n->2	
fult 	d->1	
funda	m->1	
funde	r->12	t->5	
funge	r->54	
funkt	i->32	
funna	 ->1	.->1	
funne	n->1	
funni	t->9	
fuse"	,->1	
fusio	n->8	
fusk.	H->1	
futti	g->1	
fylla	 ->23	.->1	n->2	s->9	
fylld	e->1	
fylle	r->19	
fylls	 ->2	.->1	
fyllt	 ->1	,->2	s->1	
fyra 	f->2	k->1	l->1	m->3	n->1	o->2	p->6	r->1	s->2	ä->2	å->2	
fyra,	 ->1	
fyra:	 ->1	
fyrti	o->3	
fysis	k->9	
fäder	n->1	
fäkta	r->1	
fälha	v->1	
fälld	a->1	e->1	
fälle	 ->24	.->1	n->54	r->1	t->12	
fälli	g->18	
fällt	s->2	
fält 	i->1	
fälte	t->5	
fängd	a->1	
fänge	l->1	
fär 1	,->1	/->1	0->1	
fär 7	 ->1	
fär l	i->1	
fär s	a->1	o->1	
fär t	v->2	
färan	d->1	
färd 	m->1	o->1	
färd,	 ->2	
färd;	 ->1	
färda	 ->4	n->5	s->1	t->2	
färdi	g->13	
färds	b->1	m->1	s->3	v->1	
fären	 ->1	,->2	?->1	
färer	 ->2	,->3	.->1	n->2	
färg,	 ->2	
färga	d->1	
färli	g->2	
färre	 ->2	
färsk	t->1	
färsm	ä->1	
fäst 	d->1	f->1	s->1	
fästa	 ->7	n->1	
fäste	 ->2	l->1	r->8	s->1	
fästn	i->1	
fästs	 ->1	
få 10	0->1	
få Eu	r->1	
få Go	l->1	
få al	l->1	
få an	d->1	
få ar	b->1	
få av	g->2	
få be	s->1	t->2	
få bo	r->2	
få bä	r->2	
få bö	r->1	
få de	l->1	m->1	n->5	r->1	s->3	t->3	
få di	s->1	
få do	m->1	
få ef	f->2	
få en	 ->26	o->1	
få er	s->1	
få et	t->11	
få fa	r->1	
få fi	n->1	
få fl	e->1	
få fo	l->1	
få fr	a->4	
få fu	l->1	
få fö	l->1	r->3	
få ga	r->1	
få ge	m->1	
få hi	n->1	
få hj	ä->1	
få i 	d->1	g->1	l->1	
få ig	å->1	
få in	f->1	r->1	s->1	
få ko	m->2	n->2	
få kv	i->2	
få la	n->1	
få li	k->1	
få lo	s->1	v->1	
få lä	g->2	s->1	
få ma	j->1	s->1	
få me	d->2	
få my	c->1	
få må	l->1	n->2	
få mö	j->1	
få nå	g->3	
få ob	l->1	
få om	f->1	
få or	d->2	
få os	s->2	
få pa	r->1	
få pe	r->2	
få po	s->1	ä->1	
få pr	e->1	o->1	
få pu	n->1	
få på	m->1	
få re	d->1	g->1	s->1	
få ry	g->1	
få rä	t->1	
få sa	k->1	m->1	
få se	 ->6	
få si	n->2	
få sl	u->1	
få st	a->1	o->2	r->2	ö->4	
få sä	g->2	
få så	 ->2	v->1	
få ta	 ->3	c->1	l->2	
få ti	l->16	
få up	p->1	
få ut	 ->1	f->1	
få va	r->1	
få ve	t->6	
få vi	s->3	
få vå	r->1	
få är	 ->1	
få åt	m->1	
få ök	a->1	
få, o	c->1	f->1	
få, r	ä->1	
få.Eu	r->1	
få.Gr	a->1	
få.Vi	 ->1	
fågel	l->1	s->1	v->1	
fågla	r->6	
fång 	f->1	
fånga	r->3	s->1	
fånge	t->1	
fångs	r->1	t->7	
får M	a->1	
får O	L->1	
får a	k->1	l->4	n->1	r->1	
får b	e->2	o->1	
får d	e->11	o->1	r->1	u->1	
får e	l->1	m->1	n->13	t->4	
får f	a->2	i->2	å->1	ö->1	
får g	e->2	l->1	ö->2	
får h	a->1	ä->1	å->1	
får i	 ->2	b->1	n->36	
får j	a->2	
får k	l->1	o->4	
får l	i->1	å->1	
får m	a->1	e->3	i->4	ö->2	
får n	i->1	å->2	ö->1	
får o	c->1	f->2	m->1	r->1	
får p	r->1	å->1	
får r	e->1	
får s	e->3	i->3	j->1	n->1	t->7	
får t	a->4	i->6	r->1	
får u	n->1	t->1	
får v	e->1	i->19	ä->1	
får y	t->1	
får ä	n->2	
får å	 ->1	
får, 	e->1	o->1	
får?N	ä->1	
fårkö	t->1	
fås f	ö->1	
fåtal	 ->1	
fått 	8->1	9->1	a->1	b->3	d->3	e->12	f->2	h->4	i->3	k->1	l->1	m->4	n->3	o->1	s->2	t->6	u->1	v->5	y->2	
fått.	P->1	
féren	d->1	
född.	M->1	
födde	s->1	
födel	s->2	
föder	 ->2	
födni	n->1	
födoä	m->1	
föds 	b->1	
föga 	m->1	r->1	
följa	 ->26	,->1	k->9	n->37	r->1	s->6	
följd	 ->18	.->1	e->20	r->1	s->2	å->1	
följe	l->3	r->14	
följn	i->10	
följs	 ->3	,->1	
följt	 ->2	s->2	
föll 	d->2	i->1	o->2	t->1	
föll.	H->1	
fönst	r->1	
för "	a->2	f->1	n->1	
för -	 ->3	,->1	
för 1	9->15	
för 2	0->5	7->1	9->1	
för 3	3->1	
för 5	 ->1	,->1	
för 7	5->1	6->1	
för A	g->1	l->3	
för B	e->1	i->1	o->1	r->3	
för C	S->1	e->1	
för D	a->2	e->1	
för E	C->1	G->4	U->9	r->1	u->55	
för F	P->1	o->2	ö->2	
för G	e->1	o->1	
för H	a->1	
för I	M->1	N->1	n->1	s->1	
för K	a->3	o->1	u->2	y->1	
för L	a->1	e->1	
för O	L->1	
för P	P->1	a->1	o->1	
för S	a->2	ã->1	
för T	a->1	i->6	u->1	
för V	o->1	
för W	T->1	a->1	
för a	c->1	i->1	l->130	m->2	n->40	r->12	s->2	t->724	v->23	
för b	a->1	e->39	i->9	j->1	l->3	o->2	r->4	u->14	ä->1	å->3	ö->6	
för c	e->2	h->1	i->4	
för d	a->4	e->513	i->10	j->1	o->2	u->1	ä->2	å->4	ö->1	
för e	f->1	g->3	k->16	l->4	n->130	r->30	t->50	u->1	v->2	x->3	
för f	a->10	e->3	i->10	j->1	l->3	o->8	r->29	u->1	y->1	å->5	ö->52	
för g	a->1	e->18	i->3	l->1	o->4	r->12	u->2	ä->1	
för h	a->34	e->17	i->1	j->3	o->6	u->11	ä->6	å->2	ö->4	
för i	 ->11	c->1	k->1	l->1	n->46	
för j	a->13	o->11	u->3	ä->3	
för k	a->19	l->1	n->1	o->96	r->9	u->22	v->9	ä->4	
för l	a->9	e->2	i->26	o->3	ä->11	å->7	ö->1	
för m	a->7	e->49	i->48	o->6	y->15	ä->12	å->27	ö->3	
för n	a->11	e->1	i->1	o->6	u->2	y->7	ä->34	å->11	ö->3	
för o	c->10	f->13	l->5	m->11	p->1	r->6	s->50	t->1	v->2	
för p	a->22	e->25	l->1	o->4	r->17	u->1	å->3	
för r	a->2	e->60	i->3	o->1	ä->28	å->9	ö->6	
för s	a->10	e->7	i->38	j->3	k->31	l->1	m->5	n->3	o->3	p->3	t->54	v->3	y->19	ä->14	å->12	
för t	a->3	e->2	i->41	j->7	o->1	r->25	u->3	v->4	y->3	å->1	
för u	n->33	p->7	r->1	t->60	
för v	a->22	e->9	i->49	o->1	u->1	ä->4	å->39	
för y	n->1	r->1	t->1	
för Ö	s->2	
för ä	n->7	r->23	v->1	
för å	k->1	r->12	t->21	
för ö	a->1	g->6	k->3	p->5	s->1	v->30	
för".	O->1	
för, 	1->1	a->5	e->1	f->3	h->1	i->2	k->3	o->3	s->3	t->1	u->1	v->1	ä->2	
för. 	D->1	
för.(	L->1	
för..	.->1	
för.D	e->3	i->1	
för.H	e->1	
för.J	a->1	
för.M	a->1	e->2	
för.V	i->4	å->1	
för: 	D->1	F->1	a->1	
för; 	d->1	
för?D	ä->1	
för?F	r->2	
för?I	 ->1	
för?Ä	r->1	
föra 	a->9	b->4	d->29	e->36	f->2	g->4	h->1	i->3	k->4	l->3	m->11	n->2	o->1	p->4	r->4	s->11	t->4	u->11	v->3	y->1	ä->1	å->1	ö->2	
föra,	 ->1	
föra.	D->1	J->1	O->1	
förak	t->1	
föral	l->1	
föran	d->304	k->4	l->2	s->1	
förar	b->1	n->1	
föras	 ->28	!->1	,->3	.->9	;->1	
förba	n->2	r->12	
förbe	h->6	r->27	
förbi	 ->1	f->2	g->6	n->22	s->1	
förbj	u->14	
förbl	e->1	i->14	
förbr	u->1	y->2	ä->2	
förbu	d->24	n->9	
förbä	t->78	
förd 	f->1	
förd,	 ->1	
förda	 ->5	
förde	 ->14	,->1	.->2	l->41	s->8	
fördj	u->11	
fördo	m->2	
fördr	a->162	ö->1	
fördu	b->2	n->1	
fördä	r->4	
fördö	m->20	
före 	2->1	A->1	K->1	d->5	e->1	m->2	n->2	o->3	s->2	u->4	v->2	å->1	ö->1	
föreb	i->1	r->2	y->22	
föred	r->158	ö->2	
föref	a->20	ö->1	
föreg	i->1	r->1	å->17	
föreh	a->1	
förek	o->22	
förel	e->1	i->26	s->2	
förem	å->13	
fören	a->10	i->12	k->8	l->8	
föres	a->6	k->28	l->104	p->10	t->15	ä->1	
föret	a->199	r->72	
förfa	l->1	r->75	t->7	
förfi	n->1	
förfj	o->1	
förfl	u->14	y->4	
förfo	g->18	
förfr	y->1	å->4	
förfä	k->1	r->2	
förfå	n->1	
förfö	l->5	
förgl	ö->2	
förgr	u->3	
förgä	v->1	
förha	n->92	s->3	
förhi	n->30	
förho	p->9	
förhå	l->56	
förhö	l->1	
förin	g->12	t->3	
förir	r->1	
förka	s->9	
förkl	a->76	
förkn	i->3	
förko	r->2	
förkr	o->1	
förku	n->2	
förla	g->3	
förle	g->2	
förli	g->3	k->45	s->2	t->10	v->19	
förlo	r->20	
förlu	s->9	
förlä	g->2	n->4	
förlå	t->4	
förme	d->3	n->2	
förmi	d->3	
förmo	d->11	
förmy	n->1	
förmå	 ->2	g->31	n->14	r->1	
förmö	g->1	
förna	m->1	
förne	d->2	k->8	
förnu	f->14	
förny	a->4	b->39	e->6	
förol	ä->2	
föror	d->44	e->27	s->6	
förpa	c->4	s->1	
förpl	i->21	
förr 	d->1	e->2	
förr,	 ->1	
förra	 ->42	
förre	 ->2	s->2	
förrg	å->3	
förri	n->1	
förrä	d->1	n->4	
förrå	d->1	
förs 	a->2	b->1	d->1	e->4	f->4	i->3	p->3	t->1	u->1	ä->1	ö->1	
förs,	 ->2	
förs.	 ->1	.->1	D->1	H->1	J->1	O->1	
försa	m->12	
förse	 ->2	n->27	r->1	s->1	
försi	k->66	
försk	i->2	j->1	o->2	r->4	ä->1	
försl	a->484	
förso	n->5	
först	 ->48	.->1	a->210	e->1	k->1	o->3	ä->30	å->82	ö->21	
försu	m->9	
försv	a->62	i->15	u->4	å->2	
försä	k->44	l->5	m->9	n->1	
förså	g->1	
försö	k->60	r->4	
fört 	-->1	a->1	d->1	e->2	f->3	k->1	l->1	m->9	n->2	o->1	p->1	s->3	u->1	v->1	
fört,	 ->2	
fört.	K->1	
förte	c->3	
förti	d->6	
förtj	u->1	ä->19	
förtr	o->59	y->2	ä->3	ö->1	
förts	 ->22	,->3	.->4	
förtv	i->1	
förty	d->3	
förtä	c->1	
förun	d->1	
förut	 ->2	.->1	b->1	o->9	s->62	v->2	
förva	l->48	n->6	r->1	
förve	r->22	
förvi	r->12	s->7	
förvr	ä->1	
förvä	g->14	n->28	r->11	
förvå	n->6	
förän	d->73	
förål	d->3	
föröd	a->3	e->2	
föröv	a->3	
fötte	r->3	
g (19	9->1	
g (EG	,->1	
g (ar	t->2	
g (re	c->1	
g (åt	e->1	
g - S	a->1	
g - a	t->1	
g - d	e->5	
g - g	e->1	
g - i	n->1	
g - j	a->1	
g - m	e->1	o->1	
g - o	c->6	f->1	
g - s	o->2	
g - t	r->1	
g - ä	r->1	
g -, 	i->1	ä->1	
g 1 m	e->1	
g 1 o	c->1	
g 1, 	o->1	
g 1,2	 ->1	
g 10 	k->1	r->1	s->1	ä->1	
g 10.	K->1	
g 11,	 ->1	
g 12 	i->1	
g 13 	ä->1	
g 15 	o->1	
g 17 	s->1	
g 17,	 ->1	
g 18 	h->1	i->1	
g 19 	s->1	ä->1	
g 199	4->1	9->2	
g 2, 	s->2	
g 20 	p->1	
g 200	 ->1	
g 22 	a->1	
g 22,	 ->2	
g 23 	i->1	
g 26 	m->1	
g 3 o	c->1	
g 34 	t->1	
g 37/	6->1	
g 38 	f->1	o->1	
g 38:	 ->1	
g 4 o	c->1	
g 4.I	 ->2	
g 43 	h->1	
g 44 	o->1	
g 45.	 ->1	"->1	H->1	
g 5, 	d->1	u->1	
g 6 o	c->2	
g 600	 ->1	
g 685	/->1	
g 80 	p->2	
g Det	 ->1	
g Ece	m->1	
g Eur	o->2	
g Fäs	t->1	
g Gaz	a->1	
g Hai	d->14	
g INT	E->1	
g IV 	i->2	
g Irl	a->1	
g OLA	F->1	
g Tad	z->1	
g VI 	i->1	
g [KO	M->1	
g abs	o->1	
g acc	e->3	
g ajo	u->1	
g akt	i->1	
g ald	r->2	
g all	a->2	e->1	t->6	v->1	
g an 	d->1	å->1	
g and	r->1	
g ang	å->1	
g anl	e->2	
g anm	ä->1	
g ann	a->5	
g ans	e->86	l->3	v->2	
g ant	a->5	i->1	y->1	
g anv	ä->3	
g ara	b->1	
g arb	e->5	
g art	i->1	
g ass	i->2	
g att	 ->203	
g av 	B->4	D->1	E->7	H->1	J->1	M->1	O->1	S->1	T->2	a->21	b->19	c->1	d->69	e->19	f->29	g->7	h->7	i->7	j->3	k->27	l->7	m->15	n->6	o->5	p->7	r->9	s->34	t->12	u->8	v->17	ä->1	å->4	ö->2	
g ave	u->1	
g avg	e->1	
g avl	ä->1	
g avr	u->1	ä->1	
g avs	e->2	l->4	t->1	
g avt	a->1	
g avv	i->3	
g bad	 ->2	
g bak	o->4	
g bar	a->14	
g bas	e->2	
g be 	f->1	k->1	o->1	
g bea	k->2	
g bef	a->1	i->3	o->1	r->1	
g beg	r->1	ä->5	
g beh	a->3	ö->1	
g bek	l->14	r->1	
g ber	 ->20	,->1	o->1	ä->1	ö->2	
g bes	k->2	t->5	v->1	
g bet	a->1	o->4	r->4	v->1	ä->1	
g beu	n->1	
g bev	a->1	i->1	
g bid	r->1	
g bil	d->2	
g bla	n->2	
g ble	v->5	
g bli	r->5	v->1	
g bor	 ->1	t->4	
g bra	 ->1	n->1	
g bro	t->2	
g byr	å->3	
g bär	 ->2	
g bör	 ->8	j->2	
g cit	e->2	
g dag	o->1	
g de 	f->2	m->1	s->3	t->1	v->1	
g deb	a->8	
g del	 ->9	a->9	
g dem	 ->1	o->2	
g den	 ->12	n->2	
g des	s->3	
g det	 ->14	a->1	t->4	
g dia	l->2	
g dir	e->1	
g dis	k->3	
g dju	p->1	
g doc	k->5	
g dra	 ->1	r->1	
g dro	g->1	
g dyl	i->1	
g där	 ->8	.->1	f->7	t->1	
g då 	k->1	
g död	 ->1	
g dör	 ->2	
g e.d	.->1	
g eff	e->2	
g eft	e->6	
g eko	l->1	
g ell	e->22	
g eme	l->4	
g emo	t->6	
g en 	a->1	b->1	d->2	e->1	f->1	g->1	k->2	l->2	m->4	o->1	p->1	s->6	u->1	v->2	ö->2	
g enb	a->1	
g end	a->3	
g enh	ä->1	
g ens	a->1	
g er 	a->3	g->1	k->3	o->1	
g er,	 ->2	
g erh	å->1	
g eri	n->2	
g erk	ä->2	
g ett	 ->20	
g eur	o->1	
g eve	n->1	
g ex 	a->1	
g exa	m->1	
g exi	s->1	
g exp	a->1	
g fak	t->1	
g far	t->1	
g fas	t->2	
g fel	k->1	
g fic	k->3	
g fie	n->1	
g fin	n->8	
g for	t->7	
g fra	m->27	n->1	
g fre	d->4	
g fri	t->1	
g frä	m->1	
g frå	g->28	n->56	
g ful	l->2	
g fun	d->1	g->1	k->3	
g fäl	l->1	
g får	 ->13	
g fåt	t->3	
g föl	j->1	
g för	 ->173	,->3	a->1	b->6	d->3	e->23	h->3	k->22	l->1	m->1	o->1	p->3	s->36	t->2	u->3	v->14	ä->1	
g gan	s->1	
g gar	a->3	
g gav	 ->1	
g ge 	e->1	h->1	p->1	u->1	
g gen	d->1	e->1	o->9	t->2	
g ger	 ->5	
g gic	k->1	
g giv	e->2	
g gjo	r->5	
g gla	d->2	
g glo	b->1	
g glä	d->9	
g god	t->1	
g gra	d->6	n->3	t->8	
g gro	u->1	
g gru	n->8	p->1	
g gäl	l->4	
g gär	n->8	
g går	 ->2	
g gör	a->4	
g ha 	f->1	n->1	p->1	v->1	
g had	e->5	
g han	 ->4	d->3	t->1	
g har	 ->137	m->1	
g hed	r->1	
g hel	h->3	l->1	t->7	
g hem	 ->1	
g hen	n->1	
g hie	r->1	
g hin	d->1	
g his	t->1	
g hit	 ->1	
g hjä	l->3	
g hop	p->54	
g hos	 ->3	
g hot	a->1	
g hur	 ->3	
g huv	u->1	
g häl	s->2	
g hän	d->3	s->3	v->2	
g här	 ->9	,->1	
g häv	d->5	
g hål	l->15	
g höj	d->1	
g höl	l->1	
g hör	 ->3	d->3	
g i "	g->1	
g i B	e->2	
g i D	a->1	
g i E	U->1	t->1	u->13	
g i F	r->1	
g i I	r->1	
g i K	o->3	
g i M	e->1	
g i S	h->1	t->1	y->1	
g i T	h->1	y->1	
g i Y	a->1	
g i a	k->1	l->1	n->1	r->1	v->1	
g i b	e->1	i->1	u->1	ö->1	
g i d	a->9	e->35	i->1	
g i e	g->4	n->16	t->3	
g i f	e->3	o->1	r->9	ö->11	
g i g	å->1	
g i h	a->1	e->1	ä->2	
g i j	ä->2	
g i k	a->1	l->1	o->4	r->1	
g i m	e->4	i->4	o->1	y->1	å->1	
g i o	l->1	ö->1	
g i p	r->2	u->1	
g i r	e->3	ä->4	å->1	
g i s	a->3	e->2	i->2	j->1	l->2	t->7	y->3	ä->1	å->1	
g i t	r->1	v->1	
g i u	n->1	t->4	
g i v	a->3	i->1	ä->2	å->3	
g i Ö	s->2	
g i, 	s->1	
g i.S	å->1	
g iak	t->1	
g iho	p->1	
g in 	e->1	i->6	p->2	
g ind	u->1	
g inf	i->1	o->8	ö->7	
g ing	a->2	e->2	i->1	å->2	
g ink	l->1	o->1	
g inn	a->2	e->7	
g ino	m->18	
g inr	e->1	i->2	
g ins	e->7	i->1	k->1	t->9	
g int	a->1	e->76	o->1	r->1	
g inv	ä->1	
g irr	i->1	
g ivä	g->1	
g jag	 ->2	
g jon	i->1	
g ju 	b->1	t->1	
g jur	i->1	
g jus	t->2	
g jäm	f->2	s->1	
g kam	m->1	
g kan	 ->72	s->2	
g kap	i->1	
g kar	a->2	
g kat	a->2	
g kl.	 ->2	
g kla	r->3	
g kna	p->2	
g kol	l->1	
g kom	m->57	p->7	
g kon	c->1	k->3	s->4	t->6	v->1	
g kop	p->1	
g kor	t->1	
g kos	t->3	
g kra	v->1	
g kri	t->2	
g krä	n->1	v->1	
g kul	t->2	
g kun	d->3	n->2	s->1	
g kva	l->1	r->1	
g kän	n->10	
g kär	n->1	
g köp	t->1	
g lad	e->1	
g lag	,->1	a->1	s->6	t->1	
g lan	s->1	
g lar	m->1	
g led	a->3	e->2	
g leg	a->1	i->1	
g lid	e->1	
g lig	g->1	
g lik	a->1	s->1	
g lis	t->1	
g lit	a->1	e->3	
g lyf	t->2	
g lys	s->5	
g läg	g->4	
g läm	n->2	
g län	g->3	
g lär	d->1	
g läs	a->1	t->2	
g läx	a->1	
g lån	g->1	
g låt	 ->1	e->1	
g lös	n->5	t->1	
g maj	o->1	
g mak	t->3	
g man	 ->9	.->1	d->1	
g mar	k->2	
g max	i->1	
g med	 ->62	.->1	b->1	d->3	f->1	g->1	l->3	v->4	
g mel	l->15	
g men	 ->4	,->1	a->7	i->2	
g mer	 ->9	!->1	a->1	
g mes	t->1	
g mig	 ->16	
g mil	j->2	
g min	 ->3	d->1	n->3	s->1	
g mis	s->2	
g mot	 ->21	p->1	s->5	
g myc	k->13	
g myn	d->1	
g mär	k->3	
g måh	ä->1	
g mål	e->1	
g mån	g->5	
g mås	t->34	
g möj	l->2	
g nai	v->1	
g nat	u->6	
g ned	 ->1	e->1	s->1	
g neg	a->1	
g ni 	a->1	h->2	j->1	k->1	s->1	u->1	
g niv	å->7	
g nog	 ->2	a->1	
g nol	l->1	
g not	e->4	
g nr 	1->2	
g nu 	a->1	f->2	h->1	k->2	u->1	
g num	e->1	
g nyn	a->1	
g nys	s->1	
g nyt	t->1	
g näm	n->7	
g när	 ->13	a->1	i->1	v->1	
g näs	t->3	
g någ	r->2	
g nöd	v->3	
g obe	r->3	
g och	 ->234	,->1	
g ock	s->29	
g oer	h->1	
g of 	t->1	
g off	e->2	
g oft	a->2	
g olj	a->1	
g om 	"->1	4->1	F->1	H->1	L->1	T->1	a->17	b->1	d->16	e->13	f->2	g->2	h->3	i->1	j->2	k->3	l->1	m->5	n->6	o->1	p->3	r->7	s->5	t->4	u->2	v->4	ä->1	
g om.	D->1	
g omb	a->1	u->1	
g ome	d->1	
g omf	a->1	
g omp	r->1	
g oms	ä->1	
g omö	j->1	
g ond	s->1	
g onö	d->1	
g ord	e->2	
g ori	e->1	
g oro	.->1	
g osv	.->1	
g par	l->2	
g pek	a->1	
g per	 ->1	s->9	
g pla	n->1	
g plä	d->1	
g pol	i->8	
g pos	i->3	
g poä	n->2	
g pra	x->1	
g pre	s->2	
g pri	v->1	
g pro	c->2	f->1	g->2	p->1	t->2	
g pun	k->7	
g på 	1->2	2->1	5->2	C->1	E->2	G->1	I->1	M->1	a->5	b->1	c->1	d->17	e->6	f->12	g->6	i->2	j->1	k->2	l->2	m->7	n->6	p->2	r->1	s->5	t->2	v->8	å->1	ö->1	
g på,	 ->2	
g på.	D->1	O->1	
g påb	ö->1	
g påg	å->1	
g påm	i->5	
g påp	e->2	
g pås	t->1	
g påv	e->3	
g rad	 ->1	
g ram	 ->1	.->1	
g rap	p->1	
g rat	i->1	
g rea	g->1	k->1	l->1	
g red	a->14	o->1	
g ref	e->1	o->4	
g reg	e->3	i->1	l->1	
g rek	o->4	
g rel	a->1	
g res	a->1	o->2	p->3	u->1	
g rev	i->1	
g rik	t->4	
g ris	k->3	
g rol	l->8	
g rum	.->1	
g ryk	t->1	
g räd	d->1	
g räk	n->7	
g rät	t->3	
g råd	e->3	g->2	
g rör	 ->2	a->2	
g rös	t->11	
g sad	e->11	
g sag	t->1	
g sak	 ->1	n->1	
g sam	l->2	m->4	t->3	
g sat	t->1	
g se 	a->1	
g sed	a->3	
g seg	e->1	
g sei	s->1	
g sek	t->3	
g sem	e->1	
g sen	a->1	
g ser	 ->12	v->1	
g set	t->1	
g sig	 ->1	.->1	n->3	
g sik	t->9	
g sim	m->1	
g sin	a->2	s->1	
g sit	t->3	u->2	
g sjä	l->25	
g ska	l->50	p->4	
g ske	r->1	
g ski	c->1	l->1	
g skr	i->1	
g sku	l->124	
g sky	d->1	l->1	n->1	
g skä	n->1	
g slu	k->1	t->1	
g soc	i->2	
g sol	i->2	
g som	 ->226	,->3	
g spe	c->1	
g spr	i->1	
g sta	d->1	g->1	n->2	r->1	
g sto	d->1	p->1	
g str	a->4	i->1	u->1	ä->1	
g stä	l->8	n->1	
g stå	 ->1	r->4	
g stö	d->12	r->1	
g sub	s->1	
g sva	r->3	
g syf	t->4	
g sym	p->2	
g syn	 ->1	
g sys	s->3	
g säg	a->18	e->20	
g säk	e->5	
g sän	d->1	
g sär	s->5	
g sät	t->1	
g så 	a->1	l->2	v->1	
g såd	a->1	
g såg	 ->2	
g sål	e->2	
g såv	ä->2	
g t.e	x->1	
g ta 	e->1	u->3	ö->1	
g tac	k->29	
g tag	i->4	
g tal	a->15	
g tan	k->1	
g tar	 ->6	
g tas	 ->1	
g tek	n->2	
g ter	r->1	
g tid	 ->15	e->1	i->4	s->2	
g til	l->200	
g tog	 ->1	s->1	
g tol	k->1	
g tra	n->1	
g tro	 ->1	d->1	r->114	t->1	
g trä	d->1	f->1	
g tve	k->1	
g tvi	n->1	v->2	
g tvu	n->1	
g två	 ->1	
g tyc	k->42	
g tyd	e->1	l->4	
g tyv	ä->2	
g tän	k->16	
g täv	l->1	
g und	a->1	e->20	r->5	v->1	
g upp	 ->8	.->1	e->1	f->2	g->3	m->20	r->14	s->8	
g urv	a->1	
g ut 	f->2	i->1	p->3	
g uta	n->15	
g utb	i->4	
g ute	l->1	s->1	
g utf	o->1	r->2	
g utg	å->5	ö->2	
g utk	o->1	
g utm	a->1	ä->1	
g uto	m->1	
g uts	k->1	t->6	
g utt	a->5	r->6	
g utv	e->1	ä->1	
g utö	k->1	
g vad	 ->11	
g vak	s->1	
g val	d->1	
g var	 ->7	a->9	e->1	f->1	i->3	j->1	k->1	m->2	n->1	
g ver	k->11	
g vet	 ->21	,->2	a->1	
g vi 	a->1	e->1	g->1	h->4	m->1	t->3	
g vid	 ->9	h->1	
g vil	j->28	k->3	l->236	s->1	
g vis	a->3	s->3	
g vor	e->1	
g väd	j->2	
g väg	.->3	e->1	
g väl	 ->2	d->1	k->15	
g vän	d->3	t->4	
g vär	d->1	
g väx	e->1	
g våg	a->2	
g yrk	e->1	
g ytt	e->1	
g Öst	e->2	
g ägn	a->2	
g äls	k->1	
g än 	a->1	d->1	s->1	
g änd	a->1	r->4	å->5	
g änn	u->1	
g är 	a->12	b->3	d->22	e->9	f->13	g->12	h->4	i->7	k->3	l->7	m->10	n->4	o->8	p->1	r->2	s->17	t->3	u->2	v->8	ä->1	ö->12	
g är,	 ->2	
g ärl	i->1	
g äro	 ->1	
g äve	n->6	
g å P	P->1	
g å e	n->1	
g å u	t->1	
g åkl	a->1	
g åsi	k->3	
g åst	a->1	
g åt 	E->1	a->1	b->1	d->6	e->3	f->1	i->1	k->3	m->1	u->1	Ö->1	å->1	
g åt,	 ->1	
g åte	r->3	
g åtg	ä->5	
g åts	t->1	
g öka	 ->1	r->1	
g ökn	i->1	
g öns	k->6	
g öpp	n->1	
g öve	r->17	
g övn	i->1	
g!".D	e->1	
g!Han	 ->1	
g!Jag	 ->1	
g" av	 ->1	
g" oc	h->1	
g" so	m->1	
g", m	e->1	
g", o	c->1	
g".Eu	r->1	
g".Ja	g->1	
g".Nä	r->1	
g) i 	h->1	
g) in	n->1	
g) oc	h->2	
g), t	v->1	
g).Vi	l->1	
g)Näs	t->1	
g, Br	y->1	
g, Il	e->1	
g, OL	A->1	
g, ac	c->1	
g, an	s->1	
g, at	t->9	
g, av	 ->3	
g, be	v->1	
g, bl	.->3	a->1	
g, bå	d->2	
g, bö	r->1	
g, de	 ->3	l->1	n->5	t->6	
g, dr	i->1	
g, dv	s->5	
g, dä	r->3	
g, ef	t->15	
g, el	l->3	
g, en	 ->10	
g, et	c->1	n->1	t->3	
g, fa	s->3	
g, fi	n->1	
g, fo	r->2	
g, fr	a->1	u->2	ä->1	å->4	
g, fö	r->26	
g, ge	n->2	r->1	
g, gr	u->1	ä->1	
g, gu	l->1	
g, gö	r->1	
g, ha	n->1	r->4	
g, he	r->8	
g, hå	l->1	
g, i 	b->1	d->1	e->1	l->1	m->1	p->1	s->4	u->1	
g, in	f->3	g->1	k->1	s->1	t->4	
g, ir	o->1	
g, ju	s->1	
g, jä	r->6	
g, ka	o->1	
g, kl	a->1	
g, ko	m->2	n->1	
g, kr	a->1	
g, ku	r->1	
g, le	d->1	g->2	
g, li	d->1	k->2	
g, lå	n->2	
g, ma	r->1	
g, me	d->9	n->15	r->1	
g, mi	k->1	l->3	n->1	
g, mo	d->1	t->1	
g, må	s->1	
g, nu	 ->2	
g, ny	a->1	
g, nä	m->4	r->7	
g, nå	g->1	
g, oa	k->1	
g, oc	h->35	k->1	
g, om	 ->2	
g, ot	y->1	
g, pe	n->1	
g, pr	e->1	i->1	
g, på	 ->6	
g, rä	d->1	
g, rå	d->1	
g, sa	m->2	t->1	
g, sj	u->1	
g, sk	u->4	
g, sn	a->1	
g, so	m->28	
g, sp	a->1	e->2	
g, st	r->1	ö->1	
g, sä	g->1	r->3	
g, så	 ->8	s->3	v->2	
g, ta	c->2	r->1	
g, ti	l->2	
g, tj	ä->1	
g, to	l->1	
g, tr	o->2	
g, tv	i->1	
g, tä	c->1	
g, up	p->1	
g, ut	a->12	t->2	v->2	
g, va	d->1	r->4	
g, vi	 ->2	a->1	c->1	d->1	l->16	s->1	
g, vo	r->1	
g, är	 ->6	
g, äv	e->4	
g, åt	e->2	m->1	
g, öv	e->1	
g-PM 	s->1	
g. De	n->1	t->2	
g. En	 ->1	
g. Fö	r->1	
g. Hä	r->1	
g. Me	n->1	
g. På	 ->1	
g. Sk	o->1	
g. Så	 ->1	
g.(Ap	p->2	
g.)Fö	r->2	
g.)He	a->1	
g.. (	E->2	
g.. F	ö->1	
g..(D	A->1	
g.All	a->4	
g.And	r->1	
g.Ans	v->1	
g.Arb	e->1	
g.Av 	a->2	b->1	d->1	s->1	
g.Avs	l->1	
g.Bek	v->1	
g.Bet	ä->1	
g.Bil	i->1	
g.Bri	s->1	
g.Dal	a->1	
g.Dan	m->1	
g.De 	1->1	a->1	f->1	g->1	m->2	n->1	u->1	
g.Den	 ->19	n->4	
g.Des	s->2	
g.Det	 ->56	t->11	
g.Dis	k->1	
g.Dok	u->1	
g.Dom	s->1	
g.Där	 ->1	e->1	f->6	i->1	m->1	
g.Eff	e->1	
g.Eft	e->3	
g.Eme	l->1	
g.En 	k->1	v->1	
g.End	a->1	
g.Enl	i->4	
g.Eri	k->2	
g.Ett	 ->1	
g.Eur	o->3	
g.Fle	r->1	
g.Fra	m->1	
g.Fru	 ->4	
g.Frå	g->4	
g.För	 ->10	e->2	s->4	t->1	u->1	v->1	
g.Gen	o->4	
g.Gru	n->1	
g.Han	 ->2	
g.Her	r->20	
g.Hur	 ->2	
g.Hyc	k->1	
g.Här	 ->1	
g.Hög	e->1	
g.I d	a->4	e->9	
g.I e	t->1	
g.I f	ö->1	
g.I n	o->1	
g.I s	j->2	
g.I v	i->1	o->1	
g.Ing	e->2	
g.Int	e->1	
g.Jag	 ->62	
g.Jus	t->1	
g.Kan	s->1	
g.Kat	a->1	
g.Kom	m->9	
g.Kon	k->2	
g.Kor	t->1	
g.Kos	t->1	
g.Led	n->1	
g.Lik	a->1	
g.Liv	s->1	
g.Låt	 ->3	
g.Mal	t->1	
g.Man	 ->7	
g.Mar	g->1	
g.Med	 ->2	
g.Men	 ->6	,->1	
g.Min	a->1	
g.Myn	d->1	
g.Måh	ä->1	
g.Mål	e->1	
g.Mån	g->2	
g.Möj	l->1	
g.Nat	i->1	u->1	
g.Ni 	k->2	m->1	
g.Nu 	v->1	ä->1	å->1	
g.När	 ->3	
g.Nåj	a->1	
g.Oav	s->1	
g.Och	 ->11	
g.Oft	a->1	
g.Om 	5->1	E->1	d->2	e->1	k->1	m->1	v->3	
g.PPE	-->1	
g.Par	l->2	
g.Pro	b->1	c->1	
g.På 	d->1	p->1	
g.Rap	p->1	
g.Ref	o->1	
g.Ret	r->1	
g.Sam	m->1	t->2	
g.Sed	a->1	
g.Ska	d->1	
g.Sku	l->1	
g.Slu	t->4	
g.Syf	t->1	
g.Så 	ä->1	
g.Tac	k->2	
g.Til	l->3	
g.Tit	t->1	
g.Tro	t->1	
g.Und	e->1	
g.Ung	e->1	
g.Vad	 ->4	
g.Var	 ->1	f->1	
g.Vi 	b->1	f->1	h->3	i->3	k->3	m->2	p->1	s->3	t->1	v->5	ä->3	
g.Vil	k->1	
g.Vis	s->2	
g.Vår	 ->1	a->1	
g.a. 	k->1	
g.Är 	I->1	d->1	r->1	
g.Ära	d->1	
g: De	 ->1	
g: de	t->2	
g: di	r->1	
g: et	t->1	
g: fö	r->1	
g: ha	n->1	
g: in	s->1	
g: ja	,->1	
g:Den	 ->1	
g:Det	 ->1	
g; de	n->1	t->1	
g; en	 ->1	
g; fö	r->3	
g; mi	n->1	
g; sl	u->1	
g?Den	 ->2	
g?Det	 ->2	
g?Där	f->1	
g?Fin	n->1	
g?Fru	 ->1	
g?För	 ->1	
g?Hur	 ->1	
g?Här	 ->1	
g?Jag	 ->1	
g?Jo,	 ->1	
g?Oli	k->1	
g?Tyc	k->1	
g?Vad	 ->1	
g?Är 	v->1	
gNäst	a->1	
ga "A	m->1	
ga "i	r->1	
ga - 	a->1	d->1	h->1	m->2	o->1	r->1	v->1	
ga 2 	p->1	
ga 37	0->1	
ga Be	r->2	
ga Bo	w->1	
ga EU	-->1	:->1	
ga El	i->1	
ga Eu	r->4	
ga Ev	a->1	
ga Fi	s->1	
ga Fl	a->1	o->2	
ga Fr	a->3	
ga Ha	i->2	
ga Hu	l->1	
ga Iz	q->1	
ga Ja	n->1	
ga Je	a->1	
ga Jo	n->1	
ga Ko	c->1	
ga Li	i->1	
ga Mu	l->1	
ga Na	n->1	
ga Ni	e->1	
ga Ra	c->1	
ga Ro	b->1	
ga Sa	l->1	v->1	
ga Sv	e->1	
ga ad	m->2	
ga ag	e->2	
ga ak	t->1	
ga al	l->3	
ga an	d->12	g->3	l->1	m->1	n->1	s->1	
ga ap	p->2	
ga ar	b->7	g->2	
ga at	t->121	
ga av	 ->21	f->1	s->6	t->2	
ga ba	k->2	
ga be	f->2	g->1	h->2	k->4	m->1	r->2	s->19	t->2	v->9	
ga bi	d->6	l->6	
ga bl	a->1	i->1	
ga bo	r->1	s->1	
ga br	i->3	o->4	u->1	
ga bu	d->5	
ga bä	t->1	
ga bå	t->1	
ga ce	n->1	
ga ch	a->1	
ga da	g->2	n->1	
ga de	 ->4	b->2	l->5	m->5	n->12	s->1	t->17	
ga di	r->3	s->4	
ga do	g->1	k->3	
ga dä	r->1	
ga då	 ->2	l->1	
ga ef	f->3	t->3	
ga eg	n->1	
ga ek	o->1	
ga el	e->1	l->4	
ga en	 ->8	e->1	g->1	h->1	
ga er	 ->1	,->1	f->2	
ga et	t->7	
ga eu	r->2	
ga ex	e->1	p->1	
ga fa	l->3	m->1	r->5	s->1	
ga fe	l->1	m->1	
ga fi	n->4	
ga fl	e->3	i->1	
ga fo	r->6	s->1	
ga fr	a->53	e->1	i->5	å->49	
ga få	 ->1	g->1	
ga fö	l->7	r->84	
ga ga	l->1	r->2	
ga ge	m->4	n->6	
ga gi	v->3	
ga gn	ä->1	
ga go	d->2	
ga gr	a->3	u->11	ä->2	
ga gä	l->3	
ga gå	n->3	
ga ha	d->1	n->6	r->5	
ga he	l->3	
ga hi	n->2	
ga ho	t->1	
ga hu	r->6	
ga hy	l->1	
ga hä	l->2	n->4	
ga hö	l->1	r->1	
ga i 	E->3	P->1	W->1	a->1	b->1	d->9	e->3	f->2	k->1	l->1	r->1	s->2	t->1	v->1	
ga i.	D->1	
ga ia	k->1	
ga ic	k->1	
ga id	e->1	é->1	
ga if	r->1	
ga ig	e->1	
ga im	a->1	
ga in	 ->3	d->1	f->6	g->1	l->1	o->1	r->1	s->9	t->7	v->1	
ga ir	r->1	
ga ja	,->1	g->1	
ga ju	r->1	
ga ka	n->3	t->2	
ga ke	d->1	
ga kl	a->2	
ga ko	l->2	m->18	n->20	r->1	s->8	
ga kr	a->6	i->1	
ga kv	a->2	i->2	
ga kä	r->1	
ga la	g->2	n->1	
ga le	d->2	
ga li	g->1	k->1	n->1	s->1	v->8	
ga lo	k->1	
ga lä	g->1	m->1	n->7	
ga lö	f->2	s->2	
ga ma	k->1	r->3	
ga me	d->32	g->1	k->3	n->6	r->1	t->2	
ga mi	l->4	n->4	s->2	
ga mo	n->5	t->1	
ga mu	s->1	
ga my	c->1	n->1	
ga mä	n->5	
ga må	l->6	n->2	s->1	
ga mö	j->2	
ga na	t->3	
ga ne	d->3	j->1	
ga ni	 ->1	v->2	
ga no	g->1	
ga nr	 ->24	
ga ny	a->4	h->1	å->1	
ga nä	r->6	t->2	
ga nå	g->10	
ga ob	e->1	
ga oc	h->73	k->3	
ga oe	g->1	
ga of	f->1	r->1	
ga ok	l->1	
ga ol	i->2	y->2	ö->1	
ga om	 ->82	f->2	r->8	s->2	
ga or	d->3	g->11	s->1	
ga os	s->5	ä->1	
ga pa	r->5	
ga pe	r->2	
ga pl	a->2	
ga po	l->6	
ga pr	e->1	i->2	o->16	
ga pu	n->3	
ga på	 ->8	f->1	g->1	p->1	
ga ra	m->4	p->2	
ga re	a->3	d->1	f->7	g->12	k->1	l->1	n->1	p->1	s->10	v->1	
ga ri	k->3	
ga ro	l->1	
ga ru	m->18	
ga rä	d->1	k->1	t->38	
ga rå	d->9	
ga rö	r->1	
ga sa	d->1	k->2	m->7	
ga sc	e->1	
ga se	k->8	
ga si	g->10	n->3	t->3	
ga sk	a->3	i->3	j->1	o->1	r->2	u->3	y->1	ä->1	
ga sl	u->1	
ga sm	å->1	
ga so	c->1	m->51	
ga sp	e->4	
ga st	a->4	e->1	o->4	r->5	u->2	ä->2	ö->49	
ga su	b->2	
ga sv	a->4	å->4	
ga sy	d->1	m->1	n->1	s->3	
ga sä	k->2	t->3	
ga så	 ->2	n->1	
ga ta	g->1	l->4	n->1	r->1	s->1	
ga te	c->1	l->1	m->1	x->4	
ga ti	d->4	l->24	
ga tj	ä->5	
ga to	g->1	n->1	
ga tr	a->5	
ga tu	n->2	s->1	
ga ty	c->1	n->1	
ga un	d->2	g->1	i->2	
ga up	p->19	
ga ut	 ->5	a->3	f->3	k->1	m->1	s->4	v->3	
ga va	d->2	l->3	n->4	r->1	
ga ve	c->1	r->4	t->2	
ga vi	 ->1	c->1	d->6	k->4	l->3	n->1	s->1	
ga vr	a->2	
ga vä	g->1	l->2	n->1	r->6	
ga vå	l->1	r->2	
ga yt	t->2	
ga äm	b->1	n->12	
ga än	 ->1	d->11	t->1	
ga är	 ->12	:->2	e->1	
ga äv	e->1	
ga åk	l->1	
ga år	 ->5	,->3	.->1	
ga ås	k->1	
ga åt	a->1	e->3	f->1	g->10	
ga öa	r->1	
ga ön	s->1	
ga öp	p->2	
ga ös	t->1	
ga öv	e->9	
ga! V	i->1	
ga!De	t->1	
ga!Fr	u->1	
ga!Fö	r->1	
ga!Ja	g->1	
ga!Äv	e->1	
ga, E	v->1	
ga, a	t->7	
ga, b	l->1	
ga, d	e->3	v->1	
ga, e	f->5	n->2	
ga, f	r->2	ö->7	
ga, h	a->1	e->4	
ga, i	 ->2	n->3	
ga, k	a->1	o->5	
ga, l	i->2	
ga, m	e->2	i->1	
ga, n	a->1	y->1	ä->1	
ga, o	c->12	m->4	
ga, p	e->1	r->3	
ga, r	a->1	
ga, s	o->4	ä->1	
ga, u	t->2	
ga, v	a->1	e->1	i->6	
ga, ä	g->1	
ga, å	t->1	
ga. M	e->2	
ga.(T	a->1	
ga.- 	(->1	
ga.Al	l->1	
ga.An	s->1	
ga.Av	 ->2	
ga.De	n->2	t->10	
ga.Dä	r->1	
ga.En	 ->2	
ga.Et	t->1	
ga.Fr	å->1	
ga.Fö	r->5	
ga.He	r->5	
ga.I 	d->1	e->1	p->2	r->1	
ga.In	t->1	
ga.Ja	g->14	
ga.Ma	j->1	
ga.Me	d->2	n->3	
ga.Ni	 ->3	
ga.Oc	h->1	
ga.Om	 ->2	
ga.På	 ->2	
ga.So	m->1	
ga.Så	 ->1	
ga.Ti	l->1	
ga.Ut	f->1	
ga.Vi	 ->9	a->1	d->1	k->1	
ga.Äv	e->1	
ga/ha	l->1	
ga: "	D->1	
ga: D	e->1	
ga: F	ö->1	
ga: N	ä->1	
ga: d	e->1	
ga: h	u->2	
ga: o	m->1	
ga: v	e->2	i->1	
ga; v	i->1	
ga?. 	(->1	
ga?De	t->1	
ga?Fö	r->1	
gad d	a->1	
gad m	a->2	
gad o	m->15	
gad p	o->1	
gad r	o->1	
gad s	u->1	
gad, 	a->1	
gad.D	e->1	
gad.K	o->1	
gad.M	e->1	
gad.V	i->1	
gade 	H->1	a->3	b->1	d->1	e->2	f->1	h->1	i->2	j->1	k->1	m->1	o->7	r->1	s->4	t->2	u->1	v->1	
gade,	 ->1	
gade.	D->1	
gades	 ->7	
gado,	 ->1	
gagem	a->9	
gager	a->9	
gagn 	f->3	
gagna	d->4	r->2	t->2	
gagån	g->6	
gaktu	e->1	
gal K	a->1	
gal b	e->1	
gal i	n->1	
gal k	a->1	
gal o	c->9	
gal p	r->2	å->1	
gal s	t->1	
gal t	i->1	
gal ä	r->1	
gal, 	T->1	l->1	m->1	v->1	
gala 	f->1	i->2	p->1	s->3	
galen	s->1	
galis	e->1	
galit	e->1	
gallr	i->1	
galna	 ->1	
gals 	f->2	i->1	o->2	p->1	s->1	
galt 	i->4	s->2	u->2	ä->1	
galun	d->3	
gam g	ö->1	
gam, 	e->1	
gamla	 ->28	
gamma	l->4	
gan -	 ->2	
gan 1	9->1	
gan B	r->2	
gan D	e->1	
gan J	u->1	
gan K	o->2	
gan L	a->1	
gan N	i->1	
gan P	r->1	
gan S	c->1	
gan W	i->3	
gan a	n->2	p->1	t->2	v->1	
gan c	e->1	
gan d	e->1	i->2	
gan f	i->1	l->1	r->2	ö->7	
gan g	ä->5	ö->1	
gan h	a->1	ä->1	
gan i	 ->10	n->4	
gan j	a->1	
gan k	a->1	o->2	
gan m	e->1	å->1	
gan n	ä->3	
gan o	c->11	m->93	
gan p	å->2	
gan r	ö->1	
gan s	a->2	e->1	k->2	o->7	p->1	t->1	å->1	
gan t	i->2	
gan u	r->1	t->1	
gan v	a->4	o->1	
gan y	t->1	
gan ä	r->15	v->1	
gan å	t->1	
gan",	 ->1	
gan, 	a->1	d->1	e->1	f->2	h->2	m->1	o->5	s->2	u->3	v->1	ä->1	
gan.D	e->1	
gan.E	f->1	
gan.F	ö->3	
gan.H	e->1	u->1	
gan.I	n->1	
gan.J	a->4	
gan.K	o->2	
gan.S	e->1	å->1	
gan.U	n->1	
gan.V	a->1	
gan: 	K->1	V->2	n->1	v->1	
gan; 	s->1	
gan?J	a->1	
ganda	,->2	.->1	
gande	 ->203	!->2	,->14	.->12	:->3	?->1	f->3	n->107	r->1	t->39	
ganen	 ->3	.->1	s->1	
ganet	 ->2	,->1	.->1	
gani 	s->1	
gani,	 ->4	
ganis	a->43	e->17	m->1	
gans 	o->1	
gansk	a->26	
gansv	ä->3	
gant 	s->1	
ganti	s->5	
gapro	j->1	
gar (	C->2	F->1	
gar -	 ->3	
gar E	u->2	
gar R	å->1	
gar a	l->1	n->2	t->18	v->24	
gar b	a->1	e->1	l->1	ö->2	
gar d	e->6	i->1	o->1	ä->2	å->2	
gar e	f->2	l->2	n->6	
gar f	a->1	r->7	ö->26	
gar g	e->3	j->1	å->1	
gar h	a->6	e->1	i->1	o->1	ä->1	ö->1	
gar i	 ->23	f->1	g->1	n->9	
gar j	a->5	u->1	
gar k	a->2	l->1	o->2	r->1	
gar m	a->1	e->12	i->4	o->1	å->3	
gar n	ä->4	
gar o	c->52	f->1	m->17	r->1	s->3	
gar p	å->15	
gar r	ö->1	
gar s	a->1	e->2	i->3	k->6	l->1	o->46	p->1	ä->1	å->1	
gar t	i->18	y->1	
gar u	n->1	p->2	t->2	
gar v	a->1	e->2	i->12	
gar ä	g->1	m->1	n->3	r->11	
gar å	r->1	t->1	
gar ö	v->7	
gar!M	e->1	
gar" 	o->1	
gar).	)->1	
gar, 	a->2	b->2	d->3	e->4	f->4	i->3	j->2	k->1	l->1	m->6	n->3	o->11	p->1	r->1	s->8	t->1	u->3	v->4	ä->4	
gar- 	s->1	
gar. 	A->1	V->1	
gar.)	S->1	
gar.-	 ->1	
gar..	 ->1	
gar.B	e->1	o->1	
gar.D	e->17	ä->3	
gar.E	f->1	n->2	u->1	
gar.F	P->1	r->1	ö->6	
gar.H	e->3	u->1	
gar.I	 ->5	n->1	
gar.J	a->12	
gar.K	o->2	r->1	
gar.L	i->1	å->2	
gar.M	e->1	
gar.N	i->1	
gar.O	b->1	c->1	m->4	
gar.P	å->1	
gar.R	i->1	å->1	
gar.T	a->1	i->3	
gar.U	n->1	
gar.V	a->1	i->10	å->1	
gar.Ä	n->1	
gar: 	P->1	a->2	d->2	f->1	u->1	
gar; 	i->1	
gar?J	a->1	
garan	d->2	s->1	t->93	
garde	-->1	m->1	
gare 	-->3	1->2	3->1	D->1	a->12	b->7	d->3	e->14	f->37	g->8	h->12	i->28	k->17	l->1	m->11	n->8	o->9	p->7	r->5	s->25	t->7	u->6	v->3	ä->12	å->1	ö->1	
gare!	S->1	
gare"	 ->1	
gare,	 ->27	
gare.	A->1	D->9	E->2	F->1	J->2	M->3	R->1	S->1	T->2	Ä->1	
gare:	 ->1	
gare?	K->1	
garel	ä->1	
garen	 ->19	,->4	.->7	?->1	
gares	 ->10	
garie	n->1	
garik	e->15	
garin	 ->1	
garla	n->2	
garlä	n->1	
garmy	n->14	
garna	 ->191	"->1	,->25	.->34	?->1	s->34	
gars 	E->1	o->1	s->1	u->1	v->1	
garsk	a->7	
garvä	r->1	
garäm	b->1	
gas a	t->5	
gas b	ä->1	
gas d	e->1	ä->1	
gas e	l->2	n->1	t->1	
gas f	r->4	ö->1	
gas i	 ->2	n->1	
gas k	o->2	
gas m	y->1	
gas p	a->1	o->1	å->2	
gas r	ä->1	
gas s	a->1	
gas t	a->1	i->1	y->1	
gas u	n->1	p->2	t->1	
gas v	a->2	i->1	
gas ä	r->1	
gas ö	r->1	
gas, 	a->1	e->1	f->1	i->2	n->1	o->1	p->1	
gas.D	e->1	
gas.E	t->2	
gas.J	a->1	
gas.N	ä->1	
gas.P	r->1	
gas.R	e->1	
gas.V	a->1	i->2	
gasat	t->1	
gaser	 ->2	.->1	n->2	
gaska	m->1	r->1	
gast 	g->1	
gast,	 ->1	
gaste	 ->49	,->1	.->3	:->1	
gasät	t->19	
gat E	u->2	
gat a	t->4	
gat e	n->3	
gat f	i->1	l->1	ö->2	
gat l	å->1	
gat m	i->1	o->1	
gat n	å->1	
gat o	r->1	
gat r	e->1	
gat s	i->2	o->1	t->1	
gat t	a->1	
gat, 	e->1	k->1	o->1	
gat.D	e->1	
gat.V	i->1	
gata 	m->1	
gatel	l->2	
gatio	n->16	
gativ	 ->6	.->1	a->12	i->1	t->7	
gator	i->14	n->1	
gats 	E->1	a->1	f->1	m->1	p->1	v->1	
gats.	D->1	
gau f	ö->3	
gau o	c->1	
gau s	a->3	
gau, 	L->1	e->1	h->1	s->2	
gau.E	t->1	
gauMe	d->1	
gaube	t->1	
gaus 	b->3	
gav K	i->1	
gav e	f->1	
gav h	a->1	o->1	ä->1	
gav i	 ->1	
gav m	a->1	i->1	
gav n	å->1	
gav o	r->1	
gav p	r->1	
gav s	i->1	
gav u	p->1	
gav v	ä->1	
gav, 	d->1	
gavar	a->1	
gavs 	a->1	i->2	o->1	u->1	
gbar 	m->1	n->1	
gbar.	H->1	
gbara	 ->1	.->1	
gbart	 ->4	!->1	.->5	
gbero	e->1	
gblad	 ->1	
gboxn	i->1	
gbro 	o->1	
gbygg	n->1	
gd at	t->1	
gd av	f->1	
gd ba	k->1	
gd br	a->1	
gd fo	r->1	
gd fr	a->1	å->1	
gd fö	r->2	
gd ge	m->1	
gd i 	p->2	
gd in	f->1	v->1	
gd lö	s->1	
gd ni	 ->1	
gd oc	h->3	
gd ol	i->1	
gd om	 ->1	
gd ot	i->1	
gd på	 ->2	
gd sa	k->1	
gd so	m->1	
gd yt	t->1	
gd än	d->1	
gd åt	g->1	
gd, m	e->1	
gd.De	n->1	t->1	
gda a	g->1	
gda f	ö->1	
gda h	a->2	
gda o	c->1	
gda r	ö->1	
gda t	a->1	
gda ä	n->1	
gda.V	i->1	
gde "	d->1	
gde p	å->1	
gde s	i->1	
gde v	i->1	
gden 	a->1	b->1	f->3	h->1	k->1	m->1	o->4	p->3	s->1	u->1	å->1	
gden,	 ->3	
gden.	D->3	F->1	I->1	J->1	V->1	
gdens	 ->8	
gder 	f->2	g->1	s->1	t->1	
gdes 	a->1	
gdom 	b->1	g->1	i->1	o->1	
gdom,	 ->2	
gdom.	D->1	
gdom/	r->1	
gdoma	r->7	
gdome	n->4	
gdoms	-->3	b->1	f->3	g->1	
gdpun	k->4	
gdrag	e->2	
gdsbe	f->1	
gdsko	m->1	
gdsom	r->4	
gdsre	g->2	
gdstu	r->1	
gdsut	v->1	
gdyrk	a->1	
ge Eu	r->1	
ge Fr	a->1	
ge Fu	n->1	
ge ak	t->2	
ge al	l->3	
ge an	l->2	s->1	t->1	
ge ar	b->1	t->1	
ge at	t->4	
ge be	t->1	
ge bi	d->1	s->2	
ge bu	r->1	
ge bä	s->1	
ge bå	d->1	
ge de	 ->4	m->6	n->3	s->1	t->3	
ge dä	r->1	
ge då	 ->1	
ge en	 ->13	
ge er	 ->5	a->1	f->1	
ge et	t->12	
ge fe	m->1	
ge fö	r->3	
ge ga	r->1	
ge ge	n->1	
ge gr	ö->1	
ge ha	n->1	r->2	
ge hj	ä->2	
ge hö	g->1	
ge i 	p->1	s->1	
ge in	d->1	f->1	n->1	t->1	
ge jo	u->1	
ge kl	a->2	
ge ko	l->1	m->2	n->1	
ge ku	n->1	
ge ma	n->1	t->1	
ge me	d->3	
ge mi	g->1	n->1	
ge nu	 ->1	
ge nä	r->1	
ge nå	g->2	
ge oc	h->8	
ge of	f->1	
ge om	 ->1	
ge or	d->1	
ge os	s->8	
ge pa	r->3	
ge pe	k->1	n->1	
ge pi	l->1	
ge po	l->1	
ge pr	o->2	
ge på	 ->2	,->1	
ge ra	p->1	
ge re	a->1	g->1	p->1	
ge ri	k->1	
ge ro	s->1	
ge rä	t->1	
ge rå	d->3	
ge se	d->5	
ge si	g->4	
ge sn	a->1	
ge so	m->10	
ge st	o->1	ö->1	
ge sä	g->1	
ge så	 ->2	
ge ti	l->2	
ge tr	o->1	
ge ty	d->1	
ge un	d->2	
ge up	p->2	
ge ut	 ->3	l->1	r->1	t->4	
ge va	d->1	r->2	
ge ve	l->1	
ge vi	 ->2	k->1	
ge vä	g->1	r->1	
ge vå	r->1	
ge än	 ->1	
ge är	 ->1	
ge åt	e->1	
ge, b	l->1	
ge, d	e->1	
ge, m	e->1	
ge, s	o->1	
ge. D	ä->1	
ge.He	r->1	
ge.Ja	g->2	
ge.Om	 ->1	
ge.Vå	r->1	
ge?He	r->1	
gedi 	-->1	
gedi.	D->1	
gedie	r->2	
gedig	e->1	n->1	
gefär	 ->9	l->1	
gekom	p->1	
gel r	ö->1	
gel s	o->1	
gel ä	r->2	
gel, 	å->1	
gelbr	o->1	
gelbu	n->15	
gelil	l->1	
gelli	v->1	
gellö	s->1	
gelme	d->1	
gelmä	s->2	
geln 	f->2	i->1	k->1	o->1	ä->1	
gelns	 ->2	
gelrä	t->2	
gelse	 ->4	,->4	.->1	f->2	n->2	r->6	
gelsk	-->1	a->7	t->1	y->1	
gelsm	ä->1	
gelsy	s->2	
gelve	r->19	
gelvä	n->1	
geläg	e->20	n->2	
gelän	d->1	
geman	g->13	
gemen	s->385	t->1	
gen -	 ->7	
gen 1	 ->2	,->1	2->1	3->1	4->1	7->1	8->1	9->1	
gen 2	 ->1	,->1	9->1	
gen 3	,->1	1->1	8->1	9->1	
gen 4	,->2	
gen 7	 ->1	
gen A	B->1	D->1	
gen B	a->2	
gen E	n->1	u->1	
gen F	N->1	
gen J	a->1	
gen K	i->1	
gen W	o->1	
gen a	c->1	g->1	k->1	l->1	n->17	r->1	t->56	v->214	
gen b	a->1	e->28	l->11	o->4	r->1	ä->3	ö->4	
gen d	a->3	e->14	i->2	r->2	ä->2	å->1	ö->1	
gen e	f->6	j->1	l->3	n->17	r->1	t->9	u->1	x->1	
gen f	a->5	i->4	o->1	r->19	u->4	å->8	ö->66	
gen g	a->3	e->12	j->1	l->1	o->2	r->4	ä->3	å->3	ö->6	
gen h	a->51	e->3	j->1	o->3	u->1	ä->7	å->1	ö->2	
gen i	 ->76	l->1	n->47	
gen j	a->2	u->1	
gen k	a->20	l->3	o->32	r->3	u->5	ä->4	
gen l	a->1	e->2	i->3	y->2	ä->2	
gen m	a->2	e->36	i->2	o->6	y->2	å->22	ö->3	
gen n	a->1	e->1	y->1	ä->4	å->4	ö->1	
gen o	a->1	b->2	c->69	f->2	k->1	m->19	n->1	r->2	ö->2	
gen p	a->1	e->1	l->1	o->2	r->6	u->1	å->32	
gen r	a->1	e->11	i->4	ä->6	ö->1	
gen s	a->8	e->6	i->2	k->38	l->2	o->28	t->14	u->1	ä->4	å->3	ö->1	
gen t	a->9	i->51	o->2	r->2	v->8	y->2	ä->1	
gen u	n->11	p->8	r->2	t->3	
gen v	a->21	e->6	i->19	ä->4	
gen ä	n->3	r->44	v->1	
gen å	b->1	l->1	t->3	
gen ö	v->7	
gen!R	ö->1	
gen" 	a->1	
gen",	 ->2	
gen, 	1->1	E->1	R->1	a->3	b->3	d->9	e->3	f->10	g->1	h->13	i->10	j->1	k->4	l->2	m->9	n->7	o->16	p->1	s->15	t->5	u->2	v->8	ä->5	
gen. 	H->1	J->1	N->1	O->1	V->1	
gen.(	I->1	
gen..	(->1	
gen.A	l->2	v->1	
gen.B	r->1	
gen.C	u->1	
gen.D	e->31	ä->4	
gen.E	f->1	n->3	
gen.F	a->1	r->1	ö->4	
gen.G	o->1	
gen.H	a->3	e->6	o->1	ä->2	
gen.I	 ->4	
gen.J	a->16	
gen.K	a->2	o->2	
gen.L	å->2	
gen.M	e->7	o->2	
gen.N	a->1	
gen.O	m->1	
gen.P	å->2	
gen.R	o->1	
gen.S	l->2	n->1	o->1	u->1	
gen.T	a->2	i->1	r->1	
gen.U	n->2	
gen.V	e->1	i->11	
gen.Ä	v->1	
gen: 	E->1	T->1	d->1	f->2	m->1	v->3	
gen; 	d->2	p->1	
gen?D	e->4	
gen?F	ö->1	
gen?H	e->1	
gen?V	i->1	
genI 	d->1	
gena 	e->1	
gena,	 ->1	
genan	s->1	t->1	
genar	e->2	n->1	
genas	t->10	
genav	t->3	
genbe	t->1	
genda	 ->1	
gende	r->7	
gendo	m->5	
gener	a->16	e->18	ö->4	
genet	i->1	
genfö	r->5	
gengä	l->1	
genhe	t->39	
genjö	r->2	
genko	n->1	
genkä	n->1	
genom	 ->206	,->1	.->2	a->2	b->7	d->6	f->158	g->16	l->2	r->1	s->17	t->1	
genre	g->1	
gens 	E->1	a->4	b->5	d->6	e->1	f->7	i->1	j->2	k->5	l->4	m->7	o->5	p->2	r->5	s->17	t->4	u->1	v->3	ä->3	å->2	ö->3	
gens,	 ->2	
gense	n->3	
gensk	a->23	r->1	
genst	a->1	
gensv	a->1	
gent 	s->3	å->1	
gent.	O->1	
genta	,->1	
gente	m->27	
genti	n->22	
gentl	i->43	
gentu	r->1	
genus	d->1	
genäm	t->1	
geogr	a->8	
geost	r->2	
ger -	 ->1	
ger 1	 ->1	
ger 2	0->1	
ger 5	0->1	
ger E	r->1	u->2	
ger S	c->1	
ger a	l->3	n->6	t->33	v->2	
ger b	a->6	e->3	i->1	ä->1	
ger d	e->21	i->1	o->1	
ger e	f->1	l->1	m->1	n->13	r->1	t->7	
ger f	a->2	e->1	o->2	r->17	å->1	ö->11	
ger g	a->1	e->2	r->1	
ger h	a->6	e->1	i->1	o->2	
ger i	 ->24	g->1	h->1	n->16	
ger j	a->10	u->2	
ger k	o->6	r->2	ä->1	
ger l	a->2	i->1	ä->1	å->1	
ger m	a->7	e->5	i->8	
ger n	e->2	i->4	o->1	u->2	ä->1	å->2	
ger o	c->8	l->1	m->4	s->7	
ger p	a->1	r->1	å->13	
ger r	e->3	u->2	ä->1	å->1	
ger s	a->7	e->1	i->9	o->6	t->5	å->3	ö->1	
ger t	a->2	i->15	o->2	v->1	y->2	
ger u	n->4	p->4	t->9	
ger v	a->4	i->7	o->1	ä->1	å->4	
ger ä	n->1	r->2	
ger ö	p->1	
ger! 	D->12	E->5	F->3	G->2	I->7	J->15	K->1	L->1	M->1	N->1	T->2	V->5	Ä->2	Å->1	
ger!D	e->3	
ger!E	f->1	
ger!J	a->2	
ger!V	i->1	
ger, 	"->1	a->3	b->4	d->1	e->1	f->2	g->1	h->1	i->2	k->1	m->3	n->1	o->3	r->1	s->2	t->2	v->1	
ger. 	(->1	
ger.A	t->1	
ger.D	e->2	
ger.E	u->1	
ger.F	r->1	
ger.H	e->1	ä->1	
ger.J	a->2	
ger.N	ä->1	
ger.O	c->2	
ger.P	r->1	
ger.T	a->1	i->1	
ger: 	"->1	D->1	V->2	d->1	v->1	
ger; 	d->1	
gerMe	d->1	
gera 	b->2	d->1	e->4	f->6	i->3	k->3	m->3	n->2	o->3	p->10	s->10	t->1	u->2	v->2	ö->1	
gera!	 ->1	
gera,	 ->5	
gera.	D->2	E->2	J->1	M->1	P->1	
gerad	 ->1	e->4	
geran	d->18	
gerar	 ->21	,->4	.->4	t->1	
geras	 ->1	
gerat	 ->8	,->1	.->1	
gerbe	t->1	
gerex	t->6	
geri 	k->1	m->1	o->3	
geri,	 ->5	
geri-	 ->1	
geri.	J->1	L->1	
gerib	e->4	
gerie	r->15	t->3	
gerik	o->1	
geril	a->1	
gerim	å->1	
gerin	g->289	
gerkr	a->1	
gerli	g->3	
germa	j->1	
gern 	b->1	f->1	h->1	i->2	o->2	s->2	
gern,	 ->2	
gern.	.->1	O->1	V->1	
gerna	 ->8	
gerns	 ->7	
gerpo	l->1	p->1	
gers 	a->1	
gervr	i->1	
ges a	n->3	
ges b	e->1	
ges d	e->1	i->1	ä->1	
ges e	l->1	n->1	
ges f	ö->1	
ges i	 ->6	n->1	
ges k	o->1	
ges n	y->1	å->1	
ges o	c->1	
ges p	å->1	
ges s	p->1	
ges t	i->2	
ges u	t->1	
ges y	t->1	
ges ä	n->1	
ges ö	k->1	
ges, 	j->1	o->2	
ges- 	o->1	
ges.R	å->1	
gesbe	d->1	
gesfo	r->1	
gesra	p->2	
gest 	h->1	
gest?	N->1	
gestu	n->7	
gestä	l->3	
get (	a->1	d->1	
get -	 ->2	
get 1	9->1	
get A	B->1	
get R	I->1	
get a	c->1	l->1	n->4	t->10	v->5	
get b	e->3	l->1	ö->1	
get e	f->3	m->1	n->2	
get f	a->2	i->1	r->3	å->1	ö->13	
get g	e->5	i->1	l->1	o->2	r->1	
get h	a->4	e->2	j->1	u->1	
get i	 ->8	n->13	
get k	a->4	o->3	r->2	u->1	
get l	a->2	ä->1	ö->3	
get m	a->1	e->5	o->2	å->1	ö->1	
get n	y->1	ä->1	
get o	b->1	c->14	m->9	ö->1	
get p	a->1	o->2	r->2	å->3	
get r	a->1	e->2	
get s	a->4	e->6	k->9	o->9	p->2	t->2	v->1	y->3	ä->2	å->3	
get t	a->1	e->1	i->16	r->2	v->4	
get u	n->1	p->1	t->3	
get v	a->3	i->3	ä->1	
get y	t->1	
get ä	r->10	
get ö	d->2	
get) 	s->1	
get),	 ->1	
get).	H->1	L->1	
get, 	a->2	d->3	e->4	f->1	h->3	i->2	o->5	s->4	t->1	u->1	v->1	ä->1	
get. 	V->1	
get.A	v->1	
get.D	e->9	
get.E	n->1	u->1	
get.F	r->2	ö->2	
get.H	e->2	
get.I	 ->2	
get.J	a->8	
get.K	o->2	
get.L	å->1	
get.M	e->5	
get.N	ö->1	
get.O	c->1	m->1	
get.P	a->1	å->1	
get.S	t->1	å->1	
get.T	y->1	
get.V	i->1	
get: 	t->1	
get; 	f->1	
get?V	a->1	
getan	s->1	
getar	,->1	n->1	
getbe	h->1	
getde	r->1	
getec	k->2	
geten	 ->13	.->2	
geter	i->1	
getfr	å->2	
getfö	r->9	
getko	n->16	
getkr	a->1	
getmä	s->1	
getpl	a->3	
getpo	l->1	s->10	
gets 	a->4	b->3	c->1	f->2	g->1	h->1	l->2	m->2	n->1	o->1	p->2	s->2	u->2	å->1	
getsi	t->1	
getst	ö->2	
getsy	n->1	
gett 	a->1	d->2	e->2	h->1	k->1	m->2	n->1	o->1	p->2	r->2	s->2	t->1	u->5	v->1	
gett,	 ->1	
getut	s->10	
getår	e->10	
getöv	e->1	
gfald	 ->3	,->5	e->5	i->2	
gflöd	e->1	
gfond	e->1	
gfors	 ->12	,->2	.->6	
gfris	t->1	
gfrut	a->1	
gfunk	t->1	
gfärd	s->1	
gfärg	a->1	
gförs	l->5	
gg de	 ->1	
gg dä	r->1	
gg fa	r->1	
gg fr	å->1	
gg ge	 ->1	
gg ha	r->2	
gg i 	d->3	
gg in	o->1	s->1	
gg ku	n->1	
gg lå	n->1	
gg ma	n->1	
gg mä	r->1	
gg oc	h->1	
gg på	 ->3	
gg so	m->2	
gg ti	l->4	
gg un	d->2	
gg up	p->1	
gg ut	g->1	
gg vi	 ->1	
gg" s	o->1	
gg, e	n->1	t->2	
gg, i	n->1	
gg, k	r->1	
gg, m	e->1	
gg, t	i->1	
gg, v	i->1	
gg.Dä	r->1	
gg.Fö	r->2	
gg.Ko	r->1	
gg.Ma	l->1	
gg.Nu	 ->1	
gg; f	ö->1	
gga I	z->1	
gga a	l->1	t->7	v->1	
gga b	r->1	ä->1	
gga d	e->3	o->1	
gga e	n->3	t->4	
gga f	a->2	r->45	ö->1	
gga g	r->1	
gga h	e->1	i->1	
gga i	 ->2	d->1	n->2	
gga k	e->1	o->1	v->1	
gga m	y->1	
gga n	e->2	å->2	
gga o	c->2	l->2	m->2	
gga p	å->2	
gga r	e->1	ä->1	
gga s	i->3	k->3	o->1	t->1	
gga t	i->9	o->1	y->1	
gga u	n->1	p->12	t->7	
gga v	i->5	å->2	
gga ö	v->1	
gga, 	f->1	
ggade	 ->2	s->1	
ggan 	a->1	i->1	
ggand	e->109	
ggas 	e->1	f->3	p->2	t->1	u->4	
ggas,	 ->2	
ggas.	V->1	
ggbox	n->1	
ggd i	 ->1	
ggd p	å->1	
ggde 	p->1	
ggdes	 ->1	
gge s	o->1	
ggels	e->1	
ggen 	a->1	f->2	p->1	ä->1	å->1	
ggen"	 ->1	
ggens	 ->1	
gger 	E->1	a->3	b->7	d->10	e->11	f->18	g->2	h->4	i->19	j->1	k->1	l->1	m->5	n->4	o->7	p->11	r->1	s->3	t->7	u->4	v->6	ä->1	
gger,	 ->3	
gger.	O->1	P->1	
gger;	 ->1	
gget 	a->1	s->1	v->1	
gget,	 ->1	
ggets	 ->2	
gghet	 ->4	,->1	s->1	
ggigt	 ->1	,->1	.->1	
ggjor	d->5	t->8	
gglin	g->1	
ggnad	 ->6	.->1	e->9	s->3	
ggnin	g->28	
ggor 	m->1	
ggorn	a->1	
ggrad	 ->1	
ggran	n->3	t->9	
ggres	s->1	
ggs f	a->1	r->6	
ggs i	 ->2	n->1	
ggs n	u->1	
ggs p	å->5	
ggs u	p->1	t->1	
ggs v	i->1	
ggs, 	m->1	
ggsbu	d->1	
ggsfr	å->1	
ggskr	a->1	
ggste	n->1	
ggt i	n->1	
ggt p	å->1	
ggt s	n->1	
ggt u	p->1	
ggts 	u->1	
ggå l	a->1	
ggås,	 ->1	
ggör 	a->1	e->1	i->1	s->1	v->1	
ggöra	 ->10	s->2	
ggörs	 ->3	.->1	
gh le	v->1	
gh me	d->1	
gh.Vi	 ->1	
ghet 	-->1	D->1	a->44	b->2	d->3	e->6	f->18	g->1	h->4	i->28	k->2	l->1	m->36	n->1	o->29	p->3	r->2	s->23	t->6	u->1	v->4	ä->8	å->1	
ghet!	K->1	
ghet"	 ->1	
ghet,	 ->35	
ghet.	 ->1	D->9	E->2	F->3	H->3	J->6	L->1	M->3	N->3	P->1	R->1	S->1	T->2	V->3	Å->1	
ghet?	A->1	
ghete	n->148	r->317	t->1	
ghets	c->1	f->16	k->1	o->1	p->55	s->2	t->4	å->2	
ght k	a->1	
ght t	i->1	
ghts.	A->1	
ghåll	a->2	
gi - 	a->1	v->1	
gi be	r->1	
gi fö	r->5	
gi ge	n->1	
gi gö	r->1	
gi ha	 ->1	n->1	
gi i 	k->1	
gi ka	n->1	
gi le	d->1	
gi me	l->1	
gi må	s->1	
gi oc	h->8	
gi so	m->7	
gi ti	l->2	
gi, d	e->1	
gi, e	n->1	
gi, i	n->1	
gi, k	u->1	
gi, m	e->1	
gi, o	c->1	
gi-, 	t->1	
gi.. 	(->1	
gi.Al	l->1	
gi.De	t->1	
gi.Et	t->1	
gi.Eu	r->1	
gi.Fo	r->1	
gi.Fr	u->1	
gi.Ja	g->1	
gi.Ma	n->1	
gi.Vå	r->1	
giage	n->1	
gianv	ä->6	
gibes	p->3	
gicen	t->1	
gick 	-->1	b->2	d->1	e->1	f->1	i->1	j->2	k->1	m->2	n->1	s->1	t->3	v->1	
gick,	 ->2	
gick.	A->1	Ä->1	
gieff	e->4	
gien 	d->1	j->1	o->2	ä->1	
gien,	 ->3	
gien.	D->1	
gien?	V->1	
giens	 ->1	
gier 	-->1	f->2	m->1	o->2	p->1	r->1	s->3	
gier,	 ->4	
gier.	D->1	
giera	d->1	
giern	a->1	
giet,	 ->1	
giet.	V->1	
gifor	m->1	
gift 	a->2	d->1	e->1	f->2	i->2	k->1	m->1	p->1	r->1	s->5	t->1	v->1	ä->3	
gift!	H->1	
gift,	 ->2	
gift.	A->1	D->1	E->1	J->1	O->1	V->1	
gift:	 ->1	
gifte	n->7	r->52	
gifti	g->2	
gifts	f->1	l->2	m->1	p->2	s->1	t->1	
giför	b->1	r->1	s->2	
gigan	t->5	
giggj	o->1	
gigt 	a->1	e->1	
gigt,	 ->1	
gigt.	F->1	
giimp	o->1	
gik o	c->1	
gik, 	n->1	s->1	
gik.F	r->1	
gik.H	a->1	
gik.V	i->1	
gikap	a->1	
giken	 ->2	
gikon	t->1	
gikäl	l->37	
gilla	 ->1	r->1	
gilti	g->26	
gimen	 ->1	.->1	s->1	
gimix	e->1	
gimyn	d->1	
gin f	r->1	ö->1	
gin k	o->1	
gin m	o->1	
gin o	c->2	
gin s	o->1	
gin u	t->1	
gin, 	o->2	
gin.D	e->1	
gin.S	c->1	
ginal	 ->1	e->3	i->2	v->1	
ginel	l->1	
gins 	f->1	
ginär	a->1	
gion 	a->1	d->1	e->1	f->1	g->1	i->2	r->1	s->2	t->1	u->1	
gion,	 ->3	
gion.	 ->1	D->2	G->1	J->1	U->1	V->1	
giona	l->89	
gione	n->12	r->129	
giorg	a->2	
gipla	n->1	
gipol	i->1	
gipot	e->1	
gipro	d->3	g->2	
gisek	t->4	
gisis	k->70	
gisk 	a->1	b->2	i->2	k->1	p->2	r->2	
giska	 ->36	,->1	.->2	
giskt	 ->14	,->1	.->2	
gisnå	l->1	
gissl	a->1	
giste	r->10	
gistr	e->10	
gisäk	e->7	
git -	 ->1	
git a	k->1	l->1	n->1	t->2	
git b	e->2	o->1	
git d	e->6	i->1	
git e	l->1	n->4	t->5	
git f	e->1	l->1	r->1	ö->2	
git h	u->1	ä->7	
git i	 ->5	g->1	n->1	
git k	o->1	
git l	a->1	ä->1	
git m	e->3	
git n	y->1	ä->1	å->2	
git o	c->1	m->1	
git p	l->1	å->3	
git s	i->4	k->1	t->3	
git t	i->8	
git u	n->1	p->12	
git v	a->1	i->2	
git ä	n->1	
git å	t->1	
git, 	o->1	ä->1	
git.F	r->2	ö->1	
git.I	 ->1	
git.M	e->1	
gitat	i->1	
gitim	a->6	e->5	i->6	t->1	
gits 	a->3	b->1	f->1	g->1	i->5	m->3	n->1	o->1	p->1	u->3	ä->2	
gits,	 ->2	
gits.	B->1	D->1	S->1	
gium 	a->1	o->1	
gium.	L->1	
givan	d->12	
givar	e->34	k->1	l->1	n->14	p->1	
given	 ->1	h->4	
giver	i->1	
gives	 ->1	
givet	v->25	
givit	 ->7	.->1	s->7	
givli	g->1	
givna	 ->5	
givni	n->6	
gizis	t->5	
giäke	r->1	
giåte	r->1	
giös 	s->1	
giösa	 ->2	
giöst	 ->1	
gjord	a->3	e->38	
gjort	 ->58	,->8	.->6	s->23	
gkras	c->3	
gkult	u->1	
gkörn	i->1	
gla d	e->2	
gla m	å->1	
gla p	r->1	å->3	
glad 	a->12	f->2	o->1	r->1	ö->4	
glada	 ->3	
gladd	e->2	
glade	 ->4	s->1	
gland	e->1	
glar 	i->2	k->1	m->1	o->6	s->2	u->2	v->1	
glar,	 ->3	
glar.	V->1	
glas 	a->1	i->1	p->1	
glas.	K->1	
glash	u->1	
gleda	n->3	
gledn	i->2	
gler 	b->2	f->8	h->1	i->1	n->1	o->10	p->2	s->9	v->1	ä->4	
gler,	 ->10	
gler.	A->1	D->2	E->1	F->1	K->1	
gler?	P->1	
glera	 ->4	d->1	n->1	r->4	s->7	t->2	
gleri	n->15	
glern	a->36	
glesa	 ->1	
glewo	o->2	
glig 	b->1	f->2	k->2	o->1	r->1	u->1	
glig,	 ->1	
glig.	O->1	
gliga	 ->33	,->5	.->5	
glige	n->11	
gligh	e->4	
gligt	 ->14	,->2	.->3	
gling	 ->1	,->1	
gljud	d->1	
globa	l->12	
glups	k->1	
gläde	r->19	
glädj	a->8	e->7	
gläds	 ->6	
gläng	d->1	
glömm	a->14	e->2	
glöms	k->1	
glömt	 ->4	
gm el	l->1	
gmar 	R->1	
gmati	s->3	
gmeta	l->6	
gmärk	e->1	
gmäst	a->2	
gmål,	 ->1	
gn fö	r->3	
gn oc	h->1	
gna a	n->1	t->8	
gna b	e->2	
gna d	e->1	i->1	
gna e	k->2	
gna f	o->1	ö->8	
gna g	i->1	r->1	
gna i	 ->2	d->1	n->6	
gna k	l->1	o->2	
gna l	i->1	ö->1	
gna m	e->5	o->1	y->1	ä->1	
gna n	a->2	e->1	o->1	
gna o	c->2	m->1	p->1	s->2	
gna p	e->3	r->2	å->1	
gna r	e->2	i->1	
gna s	a->1	i->5	k->1	l->1	o->1	p->2	t->1	y->2	ä->2	
gna t	i->1	
gna u	t->1	
gna v	e->1	i->1	ä->1	
gna ä	n->3	
gna å	r->3	t->2	
gna ö	v->1	
gna, 	d->1	e->1	s->1	
gna.D	e->1	
gna.I	 ->1	
gnad 	a->3	f->1	i->1	o->1	
gnad.	H->1	
gnade	 ->5	n->9	
gnads	a->1	p->1	t->1	
gnal 	f->3	o->3	s->1	t->2	
gnale	n->1	r->4	
gnand	e->1	
gnar 	a->1	b->1	d->1	e->1	h->1	j->1	k->1	m->1	o->6	r->1	s->6	ä->2	ö->1	
gnar,	 ->3	
gnar.	D->2	S->2	
gnas 	j->1	å->1	
gnas.	K->1	
gnat 	K->1	a->1	d->1	s->2	
gnati	o->1	
gnats	 ->1	
gne f	r->1	å->1	
gne i	 ->1	
gne o	c->2	
gne s	o->3	
gne-A	r->1	
gnels	e->1	
gnen 	f->1	ä->1	
gner.	D->1	
gnera	t->2	
gnes 	k->1	
gni, 	d->1	
gning	 ->43	,->9	.->9	:->1	?->1	a->58	e->46	s->56	
gnisk	a->1	
gnitu	d->1	
gnivå	g->3	
gnore	r->4	
gnutt	a->2	
gnäll	e->1	
go gr	a->1	
go so	m->1	
go år	s->1	
god a	d->1	n->1	
god b	i->1	
god f	a->1	ö->5	
god i	d->2	n->1	
god j	o->1	
god l	e->1	
god m	i->1	
god t	i->5	r->1	
god u	p->1	
god v	i->1	
god.F	a->1	
goda 	a->4	c->1	e->1	f->8	g->1	h->1	i->1	k->1	l->2	n->1	o->2	p->2	r->4	s->1	t->3	v->3	
goda.	V->1	
godkä	n->89	
godo.	D->1	H->1	O->1	
godos	e->1	
gods 	b->1	i->1	l->1	o->1	p->18	s->4	t->1	v->1	ö->1	
gods,	 ->1	
gods.	 ->1	B->1	D->1	U->1	
gods;	 ->1	
godsN	ä->1	
godse	t->2	
godta	 ->10	.->1	g->17	r->3	s->7	
godto	g->2	
godty	c->6	
gofem	 ->1	
goger	 ->1	
gogi 	-->1	
gogi.	.->1	V->1	
gogis	k->1	
goist	i->2	
golfe	n->4	
golve	t->1	
golyc	k->1	
gom a	t->1	
gom u	p->1	
gom ä	n->1	r->1	
gom.D	e->1	
gomål	 ->2	e->1	
gon a	n->10	r->1	t->1	v->3	
gon b	e->5	i->1	l->1	
gon c	h->1	
gon d	e->3	å->1	
gon e	f->4	n->2	t->1	u->1	
gon f	a->1	ö->3	
gon g	å->7	
gon h	a->1	
gon i	d->1	n->3	
gon j	u->2	
gon k	a->5	l->12	o->8	
gon l	a->1	i->1	y->1	ö->1	
gon m	o->2	å->1	ö->2	
gon n	e->1	y->4	
gon o	f->1	r->2	
gon p	l->2	r->1	å->2	
gon r	e->2	i->2	o->1	ä->3	
gon s	a->2	k->1	o->9	t->3	y->1	å->3	
gon t	a->1	i->3	j->1	r->1	ä->1	
gon u	p->2	t->1	
gon v	e->2	
gon ä	r->2	
gon å	t->1	
gon, 	a->2	e->1	o->2	
gon.A	v->1	
gon.D	e->1	
gon.H	e->1	
gon.I	 ->1	
gon.J	a->1	
gon.V	i->2	
gonbl	i->15	
gonda	g->2	
gonde	 ->1	
gonsi	n->11	
gonst	a->4	
gonti	n->39	
gor -	 ->1	
gor F	r->1	
gor a	l->1	n->1	t->3	v->5	
gor b	e->3	o->1	ö->2	
gor d	e->2	ä->1	
gor e	f->1	l->2	n->1	
gor f	o->1	r->1	ö->2	
gor g	a->1	e->2	ä->1	
gor h	a->5	ö->1	
gor i	 ->7	n->5	
gor k	o->1	
gor l	ö->1	
gor m	e->3	å->1	
gor o	c->29	m->12	
gor p	å->3	
gor s	j->1	k->1	o->50	t->1	å->1	
gor t	i->11	r->1	
gor u	r->1	t->1	
gor v	a->2	e->2	i->2	ä->2	
gor ä	n->1	r->4	
gor) 	o->1	
gor, 	a->1	b->1	e->1	f->2	i->3	m->9	o->5	r->1	s->6	u->4	v->1	ä->4	
gor. 	D->1	
gor..	(->1	
gor.D	e->10	
gor.F	e->1	r->1	ö->2	
gor.H	e->1	
gor.J	a->2	
gor.K	a->1	o->1	
gor.M	y->1	
gor.N	a->1	ä->1	
gor.S	a->1	
gor.V	e->1	i->2	
gor: 	d->1	f->1	o->1	t->1	
gor; 	j->1	
gor?,	 ->1	
gor?Ä	r->1	
gordn	i->52	
gori 	8->2	o->1	
gorie	r->5	
goris	k->1	
gorlu	n->1	
gorna	 ->22	,->4	.->4	s->1	
gors 	i->2	
gorös	 ->1	a->2	t->1	
goskr	i->1	
gosla	v->1	
got E	G->1	
got K	a->1	
got W	a->1	
got a	b->1	n->6	t->4	v->11	
got b	e->1	r->1	ä->1	
got d	i->2	o->1	
got e	l->1	x->2	
got f	e->1	o->1	r->2	ö->11	
got h	i->1	
got i	 ->2	n->2	
got j	a->4	
got k	o->2	
got l	a->1	i->1	y->1	ä->3	
got m	e->3	i->1	y->4	ä->1	å->1	
got o	c->1	k->1	m->8	
got p	a->2	o->2	r->1	
got r	e->2	
got s	k->1	l->3	n->1	o->48	p->1	t->4	v->2	y->1	ä->11	å->3	
got t	a->1	i->3	
got u	p->1	t->1	
got v	a->2	e->3	i->5	
got å	r->1	
got, 	e->2	
got.A	l->1	
got.D	e->2	
got.J	a->1	
got.S	l->1	
got.Ä	n->1	
got?N	e->1	
gott 	a->2	b->1	d->1	e->1	h->1	n->2	o->1	p->1	r->2	s->4	ä->1	
gott.	F->1	
gotte	r->1	
gottg	ö->1	
gou o	c->1	
gplan	 ->1	
gplat	s->3	
gpoli	t->2	
gra -	 ->1	
gra a	l->1	n->1	s->2	v->20	
gra b	e->3	i->1	r->1	
gra d	a->4	e->1	
gra e	n->1	r->1	u->2	x->3	
gra f	a->2	l->1	r->5	å->2	ö->1	
gra g	e->1	o->2	r->3	
gra h	a->2	
gra i	d->2	n->4	
gra k	i->1	o->8	r->1	v->1	
gra l	ä->1	
gra m	e->1	i->2	y->1	å->4	ö->1	
gra n	y->2	ä->1	
gra o	f->1	l->1	m->3	r->2	
gra p	e->2	o->1	r->5	å->1	
gra r	e->2	
gra s	a->2	e->1	i->2	l->1	m->3	o->2	p->1	t->4	y->2	ä->1	å->1	
gra t	a->1	i->4	v->1	y->1	
gra u	n->2	t->1	
gra v	a->2	e->3	i->2	
gra ä	n->3	
gra å	r->6	t->2	
gra ö	g->1	
grad 	a->3	b->1	f->2	k->1	o->2	p->2	s->1	t->2	v->1	ö->1	
grad,	 ->1	
grad.	H->1	K->1	
grade	 ->3	n->2	r->8	s->2	
gradv	i->3	
graf 	o->1	
grafi	 ->1	.->2	n->1	s->10	
grafr	y->2	
gram 	"->1	-->3	D->1	b->1	e->1	f->23	g->1	h->5	i->6	k->1	l->1	m->10	n->3	o->3	p->2	s->10	v->2	ö->1	
gram,	 ->17	
gram.	D->3	F->2	G->2	H->1	J->2	K->1	M->2	N->1	O->1	S->3	V->2	
gram?	J->1	V->1	
grama	n->1	
gramf	ö->1	
gramm	e->108	
gramp	e->3	l->8	
gramr	u->1	
gramu	t->1	
gramv	e->1	
gran 	a->4	u->1	
grand	 ->2	.->1	i->2	
grann	a->4	h->1	l->2	s->1	
grans	k->55	
grant	 ->8	.->2	e->2	
grar 	a->2	h->1	i->1	l->1	
grara	 ->1	
gras 	k->1	
grat 	E->1	b->1	f->1	i->1	
grati	o->24	s->4	
grats	,->1	
gratu	l->36	
grava	 ->1	
grave	r->4	
gravt	 ->1	
gre B	N->1	
gre a	n->1	t->1	
gre b	e->1	o->1	
gre c	h->1	
gre e	l->1	
gre f	i->2	r->3	å->1	
gre g	o->1	r->3	
gre h	a->1	
gre i	 ->3	
gre k	a->4	o->1	u->3	
gre m	y->1	
gre n	i->3	å->2	
gre o	c->2	m->1	r->1	
gre p	e->3	r->2	å->2	
gre r	ä->1	
gre s	i->2	k->3	p->1	t->3	y->1	å->1	
gre t	a->2	i->1	j->3	o->3	y->1	
gre u	t->3	
gre v	a->3	i->1	
gre ä	n->6	r->1	
gre, 	u->1	
gre.D	e->1	
gre.F	ö->1	
gre.I	 ->1	
gre.M	e->1	
gre.N	ä->1	
gre.R	å->1	
gre.S	o->1	
gre.V	i->1	
gre.Ä	v->1	
gredi	e->2	
greke	r->1	
greki	s->6	
grems	-->1	
gren,	 ->1	
grena	r->2	
grens	 ->1	
grep 	m->1	
grepp	 ->10	,->1	a->1	e->11	s->2	
grera	 ->10	d->3	r->1	s->4	
greri	n->6	
gress	 ->1	i->2	
gresu	r->1	
grifi	n->1	
grike	d->1	
gring	 ->1	
gripa	 ->15	,->1	.->1	n->19	s->1	
gripe	n->1	r->15	t->3	
gripi	t->2	
gripl	i->6	
gripn	a->1	
grips	 ->1	
grite	t->3	
grodd	a->1	
grogr	u->1	
grotu	r->1	
group	 ->1	
grov 	f->1	
grund	 ->107	,->1	.->1	?->1	a->24	b->1	e->36	f->4	k->1	l->90	o->1	p->2	s->2	t->1	v->25	
grupp	 ->56	,->9	.->2	?->1	e->107	k->1	o->1	s->4	t->1	u->1	v->1	
gruva	 ->1	
grymt	 ->1	
gräl 	g->1	i->1	
gräl,	 ->1	
gräme	l->1	
gräns	 ->2	a->62	e->34	f->2	k->7	n->12	o->1	p->1	v->1	ö->12	
gräva	 ->2	s->1	
gräve	r->1	
grå v	a->1	
gråzo	n->1	
grödo	r->1	
gröja	r->1	
grön 	v->2	
gröna	 ->12	r->1	s->1	
grönb	o->1	
grönt	 ->1	
grövs	t->1	
gs -,	 ->1	
gs al	l->1	
gs an	s->1	
gs at	t->8	
gs av	 ->4	
gs bo	r->1	
gs br	i->1	
gs da	t->1	
gs de	t->3	
gs di	m->1	
gs em	e->1	
gs en	 ->1	h->1	
gs fa	r->1	s->1	
gs fr	a->6	i->1	
gs fy	s->1	
gs fö	r->5	
gs ge	n->1	
gs hä	l->1	r->1	
gs i 	d->1	g->1	o->2	s->1	ö->1	
gs id	e->1	
gs ig	e->1	
gs in	g->2	r->1	
gs kl	.->2	
gs ku	s->1	
gs me	d->4	
gs må	s->1	
gs nu	 ->1	
gs nä	m->1	
gs oc	h->1	k->1	
gs om	 ->2	v->1	
gs po	l->1	
gs pr	o->1	
gs på	 ->6	t->1	
gs ra	m->1	
gs re	f->1	
gs si	t->1	
gs sk	a->1	u->3	
gs so	m->1	
gs st	a->1	
gs ti	l->1	
gs un	d->2	
gs up	p->3	
gs ut	 ->1	b->1	
gs va	p->1	
gs ve	r->1	
gs vi	d->1	l->1	
gs, 1	2->1	
gs, a	n->1	
gs, f	ö->1	
gs, m	e->1	
gs, u	t->1	
gs- f	ö->1	
gs- o	c->11	
gs.Fö	r->1	
gs.Ja	g->1	
gs.Lå	t->1	
gsakt	e->1	i->2	
gsalt	e->1	
gsam 	b->1	t->1	
gsamh	e->2	
gsamm	a->6	
gsamt	 ->2	.->1	
gsana	l->1	
gsanf	ö->1	
gsanl	ä->4	
gsans	p->1	v->1	
gsarb	e->6	
gsart	i->3	
gsavg	i->1	
gsavt	a->6	
gsavv	e->1	
gsbar	t->2	
gsbed	r->1	
gsbeh	o->1	
gsbel	o->1	
gsbes	t->4	ä->1	
gsbet	o->1	
gsbev	i->4	
gsbid	r->2	
gsbil	d->7	
gsbis	t->2	
gsbol	a->2	
gsbor	d->2	
gsbru	k->6	
gsbud	g->1	
gscen	t->5	
gsche	f->8	
gsdel	.->1	
gsdir	e->2	
gsdok	u->1	
gsdra	b->1	
gseko	n->5	
gsekt	o->1	
gsen 	a->1	o->1	
gsenh	e->1	
gsera	 ->1	
gserb	j->1	
gset 	b->2	e->1	m->1	
gseta	p->1	
gsfak	t->1	
gsfal	l->1	
gsfar	a->2	
gsfas	,->1	e->3	t->1	
gsfel	,->1	e->1	
gsfie	n->30	
gsfin	a->1	
gsfly	g->1	
gsfon	d->21	
gsfor	m->1	
gsfrä	m->2	
gsfrå	g->14	
gsful	l->11	
gsfun	k->1	
gsfäs	t->1	
gsför	d->1	e->4	f->12	h->11	k->1	m->5	o->1	s->200	
gsgiv	a->7	n->1	
gsgra	d->3	
gsgru	p->5	
gshan	d->1	
gsher	r->1	
gshot	a->1	
gsidi	g->3	
gsidk	a->1	
gsikt	i->7	
gsind	u->4	
gsinf	r->1	
gsini	t->1	
gsins	p->1	t->4	
gsint	e->1	
gsjur	i->2	
gskap	i->1	
gskla	r->1	u->1	
gskli	m->1	
gskoa	l->2	
gskol	o->1	
gskom	m->25	
gskon	c->1	f->133	t->1	
gskor	t->2	
gskos	t->8	
gskra	f->6	v->9	
gskri	t->1	
gskur	 ->1	
gskvo	t->1	
gskäl	 ->1	e->1	
gslag	a->1	
gslan	d->1	
gslig	t->1	
gslin	j->2	
gslis	t->47	
gsliv	e->10	
gslog	i->1	
gsläg	e->5	
gslän	d->3	
gslös	 ->2	a->1	t->2	
gsmaj	o->1	
gsmak	t->1	
gsmar	k->2	
gsmed	d->1	e->1	
gsmek	a->2	
gsmet	o->3	
gsmin	i->1	
gsmod	e->2	
gsmom	e->1	
gsmon	o->1	
gsmot	o->1	
gsmäs	s->4	
gsmål	 ->3	e->1	
gsmöj	l->3	
gsmön	s->1	
gsna 	d->2	m->1	o->1	
gsna,	 ->1	
gsnar	k->1	
gsned	l->1	
gsniv	å->5	
gsnor	m->1	
gsnyc	k->1	
gsnät	 ->1	e->1	
gsomr	å->12	
gsorg	a->2	
gspak	e->1	
gspan	e->1	
gspar	t->2	
gsper	i->3	
gspla	n->14	t->3	
gspli	k->6	
gspol	i->22	
gspri	n->1	
gspro	b->5	c->20	g->19	j->1	
gspun	k->11	
gspåf	ö->1	
gsref	o->1	
gsreg	e->3	i->2	l->2	
gsrek	o->5	
gsrep	r->2	
gsres	a->2	o->5	u->1	
gsrik	 ->5	,->1	a->3	t->6	
gsrun	d->1	
gsräd	s->1	
gsrät	t->1	
gsråd	.->1	e->2	
gssam	a->2	
gssed	 ->1	
gssek	t->7	
gssif	f->1	
gssit	u->2	
gsska	d->2	p->1	
gsske	d->3	
gsski	c->1	l->4	
gsskr	i->1	o->7	
gssky	d->1	l->2	
gsspr	i->1	
gssta	d->2	
gsstr	a->9	u->4	ä->2	
gsstå	l->1	
gsstö	d->5	
gssys	t->24	
gssäk	e->1	r->1	
gssäl	l->6	
gssät	t->8	
gst a	k->1	l->1	v->1	
gst b	e->1	
gst f	r->1	
gst g	l->1	
gst k	o->2	
gst o	l->1	
gst p	o->1	å->1	
gst r	i->1	
gst t	r->1	
gst u	p->1	
gst, 	p->1	
gst.V	a->1	
gsta 	a->1	b->1	g->2	i->1	k->1	l->1	m->7	n->1	p->1	s->1	v->1	ä->1	
gstad	g->1	
gstag	a->7	
gstan	k->1	
gsten	 ->2	a->1	d->1	
gstex	t->2	
gstid	n->2	
gstif	t->127	
gstil	l->2	
gstjä	n->5	
gstmä	n->2	
gströ	j->1	
gstäl	l->1	
gstät	h->1	
gsumm	o->1	
gsutr	u->1	y->4	
gsuts	a->1	
gsutö	v->1	
gsver	k->4	
gsvil	l->3	
gsvis	 ->23	,->6	.->1	
gsvän	l->1	
gsvär	d->3	t->2	
gsväv	n->1	
gsvåg	 ->1	
gsvår	d->1	
gsyst	e->2	
gsäga	r->3	
gsänd	r->3	
gsäre	n->1	
gsätt	a->1	
gsåre	t->1	
gsåtg	ä->5	
gsöve	r->1	
gt - 	a->2	f->1	h->1	j->1	o->1	ö->1	
gt 40	0->1	
gt 48	 ->1	
gt : 	P->1	
gt Du	b->1	
gt Eu	r->2	
gt Gr	u->1	
gt In	t->1	
gt Ky	o->1	
gt Ra	p->1	
gt Sc	h->1	
gt Th	e->1	
gt ad	e->1	
gt al	l->3	
gt an	s->4	t->1	
gt ar	b->5	t->9	
gt as	y->1	
gt at	t->197	
gt av	 ->9	f->1	g->2	h->1	s->5	t->1	v->2	
gt ba	k->2	
gt be	g->1	h->2	k->1	r->2	s->9	t->3	v->2	
gt bi	d->1	l->1	n->2	
gt bl	i->1	
gt bo	r->1	
gt br	a->2	i->1	o->1	
gt bä	t->1	
gt bå	d->1	
gt da	n->1	
gt de	 ->5	f->3	m->1	n->3	s->1	t->17	
gt di	r->3	
gt dj	ä->1	
gt dr	a->1	
gt dä	r->2	
gt ed	e->1	
gt ef	f->1	t->9	
gt eg	e->1	
gt el	l->4	
gt en	 ->3	a->1	g->1	k->1	l->1	
gt er	 ->1	k->2	
gt et	t->4	
gt eu	r->1	
gt ex	e->1	p->4	
gt fa	s->2	
gt fe	l->3	
gt fi	n->2	
gt fl	e->2	
gt fo	r->2	
gt fr	a->31	i->1	ä->1	å->5	
gt fu	l->1	
gt få	r->1	
gt fö	r->78	
gt ge	m->2	n->1	
gt go	d->39	t->1	
gt gr	u->2	ö->1	
gt gä	l->1	
gt ha	 ->2	m->1	n->3	r->9	
gt he	l->1	
gt hi	n->1	
gt hj	ä->1	
gt ho	p->1	t->4	
gt hu	r->1	
gt hä	n->2	r->1	
gt hå	l->1	
gt hö	g->3	r->2	
gt i 	F->1	T->1	b->1	d->5	e->1	f->3	h->1	k->3	r->1	s->5	u->2	
gt ic	k->1	
gt if	r->6	
gt in	 ->1	f->4	n->2	o->1	s->9	t->7	
gt ja	 ->2	
gt ju	r->1	
gt ka	m->1	n->3	
gt kl	a->1	
gt kn	y->1	
gt ko	l->1	m->10	n->3	r->2	
gt kr	a->1	i->2	ä->1	
gt kv	a->2	
gt kä	n->2	
gt li	g->1	k->1	t->3	
gt lä	g->4	n->3	
gt lå	n->3	
gt ma	n->1	
gt me	d->28	l->2	r->5	
gt mi	g->2	n->33	s->1	t->2	
gt mo	d->1	t->2	
gt my	c->5	
gt mä	r->1	
gt må	l->2	n->4	s->5	
gt mö	j->3	
gt na	m->1	
gt ne	d->6	r->3	
gt ni	 ->1	
gt no	g->8	
gt nä	r->6	
gt nå	g->1	
gt oa	c->4	
gt ob	e->2	
gt oc	h->56	k->3	
gt of	f->1	t->2	
gt om	 ->2	f->1	r->1	
gt or	d->3	i->2	ä->1	
gt os	s->1	
gt ot	i->1	y->1	
gt pa	r->5	
gt pe	r->1	
gt pl	a->1	
gt po	l->1	s->3	
gt pr	a->1	e->1	i->6	o->11	
gt på	 ->8	p->1	
gt re	f->2	g->3	s->6	
gt ru	m->9	
gt ry	k->1	
gt rä	t->1	
gt sa	d->1	g->2	m->5	t->1	
gt se	 ->1	r->1	t->2	
gt si	g->4	n->2	t->1	
gt sj	ä->1	
gt sk	a->4	e->1	j->1	y->9	
gt sl	å->1	ö->1	
gt sn	a->1	
gt so	m->27	
gt sp	a->1	o->1	
gt st	a->2	e->2	o->7	r->1	ä->1	å->1	ö->23	
gt su	b->1	
gt sv	a->2	å->2	
gt sy	f->1	s->5	
gt sä	g->2	k->1	t->29	
gt så	v->1	
gt ta	 ->3	c->2	l->3	n->2	r->1	
gt te	c->2	
gt ti	d->2	l->12	
gt to	m->1	
gt tv	å->1	
gt ty	d->2	
gt tä	m->1	
gt un	d->6	
gt up	p->10	
gt ur	 ->1	
gt ut	a->1	b->2	n->1	s->1	t->2	v->1	ö->1	
gt va	d->6	
gt ve	t->1	
gt vi	d->1	k->10	l->10	s->8	t->1	
gt vä	l->3	r->2	
gt vå	r->6	
gt yt	t->2	
gt än	d->2	
gt är	 ->14	
gt äv	e->1	
gt åt	 ->1	e->1	g->1	
gt ög	o->1	
gt ön	s->1	
gt öv	e->3	r->1	
gt!Le	d->1	
gt!Me	n->1	
gt, a	t->1	
gt, b	e->2	
gt, d	e->2	j->1	å->1	
gt, e	f->3	n->2	
gt, f	r->1	ö->5	
gt, h	a->2	
gt, i	 ->1	n->3	
gt, j	u->3	
gt, k	a->4	l->1	o->1	
gt, l	i->2	
gt, m	e->5	
gt, n	a->1	å->1	
gt, o	c->10	m->2	
gt, p	e->1	
gt, r	ö->1	
gt, s	a->1	e->2	k->2	t->1	ä->1	å->2	
gt, u	n->1	t->2	
gt, v	i->2	
gt, ä	r->2	v->1	
gt. I	 ->1	
gt.Ar	a->1	
gt.De	n->2	t->9	
gt.Di	r->1	
gt.Ef	t->1	
gt.En	 ->1	
gt.Et	t->1	
gt.Fr	u->1	å->1	
gt.Fö	r->6	
gt.Ge	n->2	
gt.He	r->4	
gt.Hu	r->1	
gt.I 	v->1	
gt.Ja	,->1	g->11	
gt.Lå	n->1	t->1	
gt.Ma	n->1	
gt.Me	d->1	n->4	
gt.Mi	n->3	
gt.Mo	t->1	
gt.Na	t->1	
gt.Nä	r->1	
gt.Of	f->1	
gt.Om	 ->2	
gt.På	 ->1	
gt.Se	d->1	
gt.So	m->1	
gt.St	a->1	ö->1	
gt.Un	d->1	
gt.Va	d->3	r->2	
gt.Vi	 ->9	
gt.Ök	a->1	
gt: d	e->1	
gt; d	e->1	
gt?Av	 ->1	
gtar 	t->1	
gtekn	o->2	
gtera	 ->6	r->1	t->1	
gtext	e->2	
gtgåe	n->11	
gtidl	i->4	
gtids	a->4	
gton 	i->1	o->1	
gton.	 ->1	
gton?	 ->1	
gtons	 ->1	
gtran	s->2	
gts -	 ->2	
gts 8	0->1	
gts a	t->1	v->4	
gts b	ä->1	
gts f	r->17	
gts h	ä->3	
gts i	 ->2	n->1	
gts n	e->1	
gts o	c->1	
gts t	i->1	
gts u	n->1	p->1	
gts, 	i->2	
gtvis	 ->101	,->5	.->2	
gtvät	t->4	
guds 	s->2	
gue, 	v->1	
gueir	a->1	
guer 	h->1	t->1	
guesa	 ->1	
gulde	n->1	
gult 	k->1	
gumen	t->17	
gummi	p->1	
guro,	 ->1	
gusta	a->1	
guver	n->1	
gvari	g->6	
gvatt	n->1	
gverk	 ->1	
gynna	 ->6	d->6	r->4	
gynns	a->3	
gypte	n->2	
gäck 	m->1	
gäld 	å->1	
gälla	 ->9	:->1	n->19	
gälld	e->11	
gälle	r->362	
gälln	i->1	
gällt	 ->2	
gänge	s->1	
gängl	i->23	
gär a	t->2	v->1	
gär b	a->1	
gär d	e->1	
gär e	m->1	n->2	
gär o	c->1	
gär s	n->1	
gär ö	k->1	
gär.V	i->1	
gära 	a->3	d->1	e->2	o->1	ä->2	
gära,	 ->1	
gäran	 ->14	,->3	.->3	?->1	
gäras	 ->3	
gärd 	2->1	a->1	d->1	e->1	f->1	k->1	o->3	s->2	v->2	
gärd,	 ->6	
gärd.	D->2	H->1	I->1	J->1	
gärd;	 ->1	
gärda	 ->1	r->1	s->1	
gärde	 ->3	n->1	r->206	
gärds	 ->1	l->1	o->1	p->7	
gärna	 ->32	
gärni	n->1	
gärs 	f->1	
gärt 	a->1	e->3	i->1	o->2	
gärt,	 ->2	
gärt.	J->1	
gäves	 ->1	
gå Ki	n->1	
gå an	 ->1	
gå at	t->1	
gå be	t->2	
gå de	 ->1	n->1	
gå en	 ->3	
gå et	t->2	
gå fr	a->4	å->2	
gå fö	r->3	
gå gr	u->2	
gå he	m->1	
gå i 	c->1	d->4	e->3	
gå ig	e->4	
gå in	 ->15	
gå la	n->1	
gå lä	n->4	
gå lå	n->1	
gå me	d->3	
gå oc	h->2	
gå of	f->1	
gå på	 ->1	
gå sa	m->1	
gå sn	a->1	
gå so	m->2	
gå så	 ->1	d->1	v->1	
gå ti	l->13	
gå un	d->1	
gå ut	 ->2	,->1	ö->1	
gå vi	d->3	l->1	
gå åt	 ->1	
gå.At	t->1	
gå.Dä	r->1	
gå.Fö	r->1	
gå.Nä	r->1	
gå.Om	 ->1	
gå.So	c->1	
gå.Vi	 ->1	
gåend	e->101	
gång 	-->1	a->7	b->5	d->6	e->5	f->11	h->6	i->5	k->4	m->2	n->1	o->2	p->5	r->2	s->9	t->23	u->6	v->4	ä->4	ö->1	
gång"	.->1	
gång,	 ->8	
gång.	D->5	F->1	H->1	J->1	N->1	O->1	T->1	V->2	
gånga	r->13	
gånge	n->43	r->25	
gångk	ö->1	
gångn	a->2	
gångs	 ->3	b->3	p->15	r->14	s->8	ä->1	
går a	t->8	v->1	
går b	e->3	r->2	
går d	e->10	i->3	ä->1	å->1	
går e	n->3	
går f	e->1	r->5	ö->4	
går g	e->2	
går h	e->2	ä->1	
går i	 ->11	f->2	g->2	n->8	
går j	a->2	
går k	v->1	
går l	y->1	ä->1	å->1	
går m	e->2	o->5	
går n	u->1	ö->1	
går o	c->8	m->1	s->1	
går p	r->1	å->3	
går r	e->1	
går s	n->1	o->1	t->1	ä->1	å->2	
går t	i->17	
går u	t->12	
går v	a->1	i->1	ä->1	
går ä	v->1	
går å	t->2	
går ö	v->1	
går, 	a->1	k->1	o->1	p->1	
går. 	J->1	
går.D	e->1	
går.I	 ->1	
går.J	a->2	
går.V	i->2	å->1	
gård 	t->1	
gårda	g->2	r->2	
gårde	n->1	
gås a	l->1	
gås i	 ->1	g->1	
gås o	c->1	
gås, 	i->1	
gås: 	a->1	
gått 	a->1	e->7	f->2	i->7	m->4	n->2	o->3	s->1	t->2	y->1	
gått.	D->1	I->2	
gåtts	 ->3	
gåvor	 ->1	.->1	
gömma	s->1	
gömme	r->2	
gömts	 ->1	
gör "	K->1	
gör 3	 ->1	
gör 8	1->1	
gör E	u->1	
gör a	l->6	n->4	r->1	t->18	v->1	
gör b	o->1	
gör d	e->52	u->1	ä->3	
gör e	n->14	t->6	
gör f	ö->4	
gör g	e->2	r->3	
gör h	a->1	e->1	u->1	ä->3	
gör i	 ->3	n->2	
gör k	o->1	ä->1	
gör m	a->3	e->2	i->5	ä->1	
gör n	e->1	ä->1	å->5	
gör o	c->2	r->1	s->1	
gör p	o->2	r->1	å->1	
gör r	i->1	
gör s	a->2	i->3	j->1	ä->1	å->1	
gör t	i->2	r->1	v->1	
gör u	n->1	p->1	t->1	
gör v	a->2	i->7	å->1	
gör y	t->1	
gör ä	n->1	r->3	
gör, 	a->1	e->1	
gör.D	e->3	
gör.E	t->1	
göra 	-->1	E->3	a->13	b->3	d->69	e->35	f->20	g->4	h->5	i->9	k->9	l->2	m->27	n->21	o->4	p->2	r->2	s->23	t->5	u->5	v->8	y->1	ä->4	å->1	
göra,	 ->7	
göra.	D->3	E->1	H->1	I->1	J->3	L->1	N->1	P->1	S->1	
göra?	J->1	
göran	d->58	
göras	 ->26	,->1	.->7	
görel	s->5	
görin	g->2	
görli	g->2	
görs 	a->7	e->2	f->3	i->3	m->2	o->1	p->2	ö->1	
görs,	 ->4	
görs.	D->1	J->1	V->1	
h "Ur	b->1	
h "sk	a->1	
h "ti	l->1	
h (A5	-->1	
h - e	f->1	
h - s	o->2	
h -or	g->3	
h 0 p	r->1	
h 1-2	 ->1	
h 10 	m->1	
h 100	 ->1	
h 138	.->1	
h 14 	t->1	
h 16 	p->1	
h 17 	d->1	
h 17.	S->1	
h 19 	p->1	
h 194	.->1	
h 199	2->1	5->1	6->2	7->1	9->6	
h 2 i	 ->1	
h 2, 	v->1	
h 2.D	e->1	
h 20 	n->1	ä->1	
h 200	 ->1	
h 21 	o->2	ä->1	
h 22.	Ä->1	
h 25.	D->1	
h 27 	d->1	
h 29 	m->1	
h 3.I	 ->1	
h 30 	i->1	
h 300	 ->1	
h 33 	a->1	
h 34 	i->1	
h 35.	S->1	
h 3: 	f->1	
h 4.J	a->1	
h 41 	r->1	u->1	
h 45 	a->1	g->1	
h 45,	 ->1	
h 45.	V->1	
h 47 	g->1	
h 48 	g->1	i->1	
h 5 v	i->1	
h 5.E	m->1	
h 53 	p->1	
h 60-	t->1	
h 68 	a->1	
h 7 -	 ->1	
h 7 f	ö->1	
h 7 i	 ->1	
h 7 o	c->1	
h 7, 	d->1	o->1	
h 8 ä	r->1	
h 8, 	s->1	
h 82 	h->1	i->1	
h 82)	 ->1	
h 82,	 ->3	
h 86 	i->2	
h 89 	i->1	
h 9 i	n->1	
h 9 m	i->1	
h 92/	4->1	
h 94 	p->1	
h Alb	a->1	
h Alt	e->1	
h Ams	t->1	
h Ank	a->1	
h BP,	 ->1	
h Bas	s->1	
h Bel	g->1	
h Bra	s->1	
h Bro	k->1	
h Bul	g->1	
h C. 	E->1	
h CEC	A->1	
h Cau	d->1	
h Cyp	e->1	
h Dan	m->2	
h De 	g->1	
h Dem	o->1	
h ELD	R->2	
h EU 	g->2	
h EU-	u->1	
h EUG	F->1	
h Edi	n->1	
h Elm	a->2	
h Emi	l->1	
h Erk	k->1	
h Eti	o->1	
h Eur	o->24	
h FN:	s->1	
h FPÖ	 ->1	
h Fin	l->2	
h Fra	n->10	
h Fru	t->1	
h Gal	i->1	
h Gaz	a->1	
h Gem	e->1	
h Gol	f->1	
h Gra	c->1	
h Gre	k->1	
h Gru	p->1	
h Hel	s->1	
h Hit	l->1	
h Huh	n->1	
h II 	h->1	
h II,	 ->1	
h Ind	i->2	
h Int	e->2	
h Irl	a->2	
h Isr	a->5	
h Ita	l->1	
h Jac	k->1	
h Jör	g->1	
h Kas	p->1	
h Kin	a->2	n->3	
h Kir	g->1	
h Kou	c->1	
h Kul	t->1	
h Lan	g->3	
h Lei	n->5	
h MAR	P->1	
h Mad	a->1	e->2	
h Med	e->1	
h Nor	g->1	
h Nya	 ->1	
h OLA	F->1	
h One	s->1	
h PPE	 ->1	
h PSE	-->2	
h Pac	k->1	
h Pak	i->3	
h Pal	a->1	e->3	
h Par	i->1	
h Pet	r->1	
h Por	t->3	
h Prí	n->1	
h Raf	a->2	
h Rap	k->1	
h Sam	m->10	
h Sch	r->1	u->1	
h Sim	p->1	
h Sjö	s->1	
h Soc	i->1	
h Spa	n->1	
h Sto	r->2	
h Swo	b->1	
h Syd	o->1	
h Syr	i->7	
h Tad	z->1	
h Tai	w->1	
h Tam	m->2	
h Tsa	t->1	
h Tur	k->1	
h Tys	k->2	
h Uzb	e->1	
h Vit	o->1	
h Väs	t->1	
h Wye	-->1	
h X o	c->1	
h abs	o->1	
h acc	e->1	
h adm	i->1	
h adv	o->1	
h age	r->2	
h akt	i->2	u->1	ö->1	
h ald	r->2	
h all	a->4	m->1	r->1	t->10	
h amb	i->4	
h ana	l->3	
h and	a->1	r->26	
h ang	e->1	r->1	å->1	
h ann	a->2	o->1	
h anp	a->2	
h ans	e->4	l->1	t->3	v->4	
h ant	a->2	i->3	
h anv	ä->3	
h apr	o->1	
h arb	e->14	
h art	i->1	
h ass	o->1	
h asy	l->3	
h att	 ->148	,->2	
h av 	E->2	a->1	c->1	d->6	e->1	f->1	s->1	u->1	
h avd	e->1	
h avg	i->1	ö->2	
h avl	ä->1	
h avr	a->1	e->1	
h avs	e->2	i->1	k->1	l->1	t->1	
h avt	a->3	
h avv	e->1	i->1	
h bad	 ->1	
h bag	a->1	
h bal	a->3	
h ban	k->1	
h bar	a->3	n->3	t->1	
h bea	k->1	
h bed	r->4	ö->4	
h bef	o->5	r->1	ä->1	
h beg	r->2	
h beh	o->2	å->1	ö->4	
h bek	r->2	y->1	ä->1	
h bel	o->1	y->1	ö->2	
h bem	ö->1	
h ber	 ->1	i->1	ä->1	
h bes	l->1	t->3	v->1	
h bet	a->1	y->2	ä->3	
h bev	i->4	
h bid	r->6	
h bil	i->2	l->2	
h bl.	a->2	
h bla	n->2	
h bli	 ->1	r->2	
h blu	n->1	
h bor	d->2	
h bos	t->1	ä->1	
h bot	t->1	
h bra	n->1	
h bri	n->1	s->1	
h bro	d->2	
h bru	k->2	
h brä	n->3	
h brå	d->5	
h bud	g->3	
h byr	å->2	
h bäs	t->2	
h bät	t->2	
h båt	a->1	
h bör	 ->3	j->3	
h cal	v->1	
h can	n->1	
h cen	t->6	
h che	f->1	
h cho	c->1	
h dag	 ->1	e->1	
h dam	m->1	
h dat	o->1	
h de 	1->1	a->4	b->1	d->1	e->2	f->6	g->1	h->5	i->5	k->8	l->7	m->8	n->2	o->2	p->4	s->16	t->1	u->1	v->2	y->2	å->2	ö->2	
h deb	a->2	
h dec	e->1	
h del	a->1	s->4	t->2	v->1	
h dem	o->10	
h den	 ->98	n->10	
h der	a->12	
h des	s->34	t->1	
h det	 ->166	,->1	a->2	s->1	t->38	
h dia	l->1	
h dio	x->1	
h dir	e->3	
h dis	k->4	
h dit	 ->2	
h dju	p->1	r->2	
h djä	r->1	
h dom	a->1	s->8	
h dra	 ->1	b->1	
h dri	c->1	v->1	
h duk	t->1	
h dyr	t->1	
h där	 ->11	,->1	e->2	f->33	i->10	m->25	v->1	
h då 	a->1	b->3	d->1	h->2	i->4	k->1	m->2	o->1	r->3	s->1	t->1	v->1	ä->1	
h då,	 ->1	
h dål	i->1	
h döt	t->1	
h eff	e->16	
h eft	e->18	
h ege	n->1	
h ej 	b->1	
h eko	n->21	s->1	
h ele	k->1	
h en 	a->1	b->4	d->1	e->6	f->4	g->7	h->3	i->3	k->4	m->3	n->2	o->2	p->3	r->3	s->17	t->1	u->2	v->3	ö->1	
h en,	 ->1	
h ena	t->1	
h end	a->2	
h ene	r->2	
h eng	a->2	
h enh	e->4	ä->1	
h enk	l->1	
h enl	i->2	
h ens	t->1	
h ent	y->2	
h env	i->1	
h er 	s->2	
h er.	K->1	
h era	 ->2	
h erb	j->2	
h erf	a->3	
h erh	å->1	
h erk	ä->2	
h ers	ä->3	
h ert	 ->1	
h eti	s->1	
h ett	 ->32	
h eur	o->9	
h exa	k->1	m->1	
h exp	e->1	
h ext	r->1	
h fak	t->2	
h fal	l->1	s->1	
h far	l->2	v->1	
h fas	t->1	
h fat	t->5	
h fau	n->1	
h fed	e->1	
h fel	a->1	
h fem	t->1	
h fie	n->1	
h fin	a->6	n->2	
h fir	a->1	
h fis	k->2	
h fle	r->2	x->6	
h flo	d->1	
h fly	k->1	
h fod	e->1	
h fol	k->2	
h for	s->1	t->3	
h fra	m->23	n->2	
h fre	d->2	
h fri	 ->1	h->4	v->1	
h fro	d->2	
h fru	k->4	
h frä	m->34	
h frå	g->7	n->3	
h ful	l->5	
h fun	g->1	k->1	
h fus	i->2	
h fyr	a->1	
h fys	i->1	
h fäl	t->1	
h få 	d->1	e->1	p->1	t->1	
h fåg	e->1	
h får	 ->4	k->1	
h fåt	t->2	
h föl	j->5	
h för	 ->55	a->4	b->8	d->6	e->13	f->4	h->7	i->1	k->2	l->2	m->5	n->1	o->1	p->1	r->1	s->40	t->3	v->9	
h gag	n->1	
h gar	a->6	
h ge 	d->4	f->1	k->1	r->2	t->1	u->1	
h gem	e->6	
h gen	e->3	o->15	t->2	
h geo	g->1	
h ger	 ->3	
h ges	 ->3	
h giv	e->4	
h gjo	r->1	
h gla	s->1	
h glo	b->1	
h glä	d->1	
h god	k->1	
h got	t->1	
h gra	n->2	
h gru	n->3	p->2	
h grä	n->2	
h grö	n->1	
h gäl	l->1	
h gå 	o->1	v->1	
h går	 ->1	d->1	
h gör	 ->6	a->11	
h ha 	e->1	r->1	
h ham	n->1	
h han	 ->4	d->9	s->10	t->4	
h har	 ->16	
h hel	a->4	s->1	t->2	
h hen	n->4	
h her	r->43	
h hit	t->1	
h hjä	l->4	
h hob	b->1	
h hon	 ->1	
h hop	p->5	
h hot	 ->1	a->3	
h hum	a->1	
h hun	d->1	
h hur	 ->11	
h hus	ö->1	
h huv	u->1	
h hyg	i->1	
h hyl	l->1	
h häl	s->1	
h här	 ->6	m->1	t->1	
h hål	l->16	
h hög	e->3	r->1	
h höj	a->1	e->1	
h i G	r->1	
h i M	e->1	
h i N	e->1	
h i S	t->1	
h i T	h->1	y->1	
h i a	l->1	
h i b	u->1	
h i d	e->13	
h i e	n->3	
h i f	a->1	r->2	ö->2	
h i g	a->1	e->1	o->1	r->1	
h i h	ä->1	
h i i	c->1	
h i j	u->1	
h i k	o->1	
h i l	i->1	
h i m	e->1	
h i n	å->1	
h i o	r->1	
h i p	a->1	r->1	
h i r	a->1	
h i s	a->1	e->1	k->1	t->5	y->6	å->2	
h i u	t->2	
h i v	i->6	ä->2	
h i ö	r->1	v->3	
h ibl	a->3	
h ick	e->2	
h ide	e->2	
h idr	o->3	
h ifr	å->1	
h ikr	a->1	
h ill	v->1	
h ima	g->1	
h imm	a->1	
h ind	i->1	u->5	
h inf	o->5	ö->6	
h ing	a->1	e->4	r->2	
h inh	ä->1	
h ini	t->2	
h ink	o->1	
h inl	e->1	
h inn	e->3	
h ino	m->7	
h inp	r->1	
h inr	e->1	i->9	ä->2	
h ins	a->2	e->1	p->1	t->5	y->3	
h int	a->1	e->69	r->2	
h inv	a->5	e->1	
h irl	ä->1	
h isr	a->2	
h jag	 ->149	
h jor	d->5	
h jur	i->3	
h jus	t->4	
h jäm	s->1	
h kab	i->1	
h kam	p->1	
h kan	 ->7	d->1	s->6	
h kap	i->1	
h kar	a->1	t->1	
h kat	a->1	o->1	
h kin	e->1	
h kla	r->3	
h klo	k->1	
h knu	t->1	
h koh	e->1	
h kol	l->2	
h kom	m->57	p->4	
h kon	c->4	f->1	k->12	s->25	t->13	v->2	
h kor	r->4	t->1	
h kos	t->3	
h kra	f->2	v->3	
h kre	a->1	
h kri	m->1	s->2	t->3	
h kry	p->1	
h krä	n->1	v->3	
h krå	n->1	
h kul	t->3	
h kun	n->3	s->1	
h kva	l->2	
h kvi	c->1	n->7	
h käl	l->1	
h käm	p->1	
h kär	a->2	n->2	
h kör	 ->1	
h lag	a->2	e->1	s->3	
h lan	d->9	s->1	
h lar	m->1	
h led	a->8	e->3	n->2	
h leg	i->1	
h lem	.->1	
h lev	a->1	e->1	
h lik	a->2	n->3	v->2	
h lit	t->1	
h liv	s->3	
h lju	d->1	
h loc	k->1	
h lok	a->4	
h los	s->1	
h lov	 ->1	a->2	
h luk	t->1	
h lyc	k->3	
h läc	k->1	
h läg	e->1	g->5	
h läm	p->2	
h län	g->1	
h lär	o->1	
h lät	 ->1	t->2	
h lån	g->11	
h lås	e->1	
h låt	 ->4	a->3	
h lös	a->1	e->1	
h mak	t->1	
h man	 ->17	d->1	
h mar	k->1	
h mat	e->1	
h med	 ->67	,->3	b->6	d->2	e->35	f->1	l->6	v->2	
h mek	a->1	
h mel	l->3	
h men	a->1	i->1	
h mer	 ->14	a->1	
h met	o->1	
h mig	.->1	
h mil	i->1	j->16	l->1	
h min	 ->6	a->2	d->4	i->1	o->1	s->3	
h mis	s->3	
h mod	e->4	
h mon	e->4	o->1	t->1	
h mor	a->1	d->2	
h mot	 ->3	i->1	o->2	s->4	t->1	
h mus	s->1	
h myc	k->7	
h myn	d->1	
h män	 ->3	.->2	n->6	
h mär	k->1	
h måh	ä->1	
h mål	 ->3	,->2	s->1	
h mån	a->2	g->8	
h mås	t->5	
h möj	l->8	
h mör	d->1	
h nat	i->4	u->7	
h ned	s->1	
h neg	a->1	
h neo	n->1	
h nep	o->4	
h neu	t->1	
h ni 	b->1	h->2	m->1	s->2	v->1	ä->1	
h niv	å->1	
h nog	g->3	
h nor	d->1	
h not	e->1	
h nu 	E->1	a->1	b->2	d->1	e->1	k->1	p->1	s->2	å->1	
h nya	 ->4	n->1	
h nye	t->1	
h nyl	i->3	
h nyn	a->2	
h nyt	t->2	
h näm	n->1	
h när	 ->12	i->2	
h nät	s->1	t->1	
h någ	o->4	r->1	
h nöd	v->6	
h oac	c->4	
h obe	r->1	s->1	
h och	 ->2	
h ock	s->8	
h ode	l->1	
h oeg	e->1	
h oek	o->1	
h off	e->2	i->1	
h oft	a->2	
h ofö	r->1	
h ojä	m->1	
h okl	a->3	
h okr	ä->1	
h oli	k->5	
h olj	e->1	
h oly	c->2	
h om 	P->1	a->1	b->1	d->7	i->1	k->2	n->2	o->1	r->1	s->2	v->3	
h omb	u->2	
h ome	d->3	
h omf	a->5	
h omg	e->1	i->1	å->1	
h omr	i->1	ö->1	
h oms	o->2	t->2	
h ont	.->1	
h ope	r->1	
h opp	o->1	
h ord	a->1	f->2	
h org	a->2	
h ori	g->1	
h ors	a->1	
h orä	t->1	
h oss	 ->2	
h ost	r->1	
h osä	k->2	
h otv	e->1	
h oum	b->1	
h oun	d->1	
h out	n->1	
h pap	p->1	
h par	l->20	t->3	
h pas	s->1	
h pek	a->2	
h per	 ->2	m->1	s->4	
h pla	c->1	
h pli	k->2	
h pol	i->15	
h pos	i->1	t->1	
h pra	g->1	
h pre	c->1	s->2	
h pri	c->1	n->4	o->3	
h pro	b->3	c->2	d->6	g->6	p->1	t->1	
h prä	g->1	
h på 	a->2	d->2	e->2	f->2	g->2	h->1	m->3	s->6	t->1	v->1	
h påm	i->1	
h påp	e->1	
h pås	k->1	t->1	
h påt	a->1	
h påv	e->1	i->1	
h rap	p->1	
h ras	i->4	
h rat	i->2	
h rec	i->1	
h red	o->2	
h ref	o->4	
h reg	e->11	i->19	l->4	
h rej	ä->1	
h rek	o->2	
h rel	e->2	i->1	
h ren	a->1	o->1	t->3	
h rep	r->1	
h res	i->1	p->8	u->2	
h rev	i->2	
h rig	o->1	
h rik	a->1	t->5	
h rin	g->1	
h ris	:->1	
h rol	l->1	
h rom	e->3	
h rut	i->1	
h räd	d->1	
h räk	n->1	
h rät	t->59	
h råd	 ->1	e->36	f->1	s->1	
h rös	t->1	
h sam	a->10	f->1	h->3	l->3	m->9	o->2	r->2	t->10	
h san	k->1	s->2	
h se 	o->1	t->4	v->1	
h sed	a->9	
h sek	r->2	t->1	
h sel	e->1	
h sen	a->1	
h ser	 ->2	i->2	v->1	
h set	t->1	
h sex	i->1	u->1	v->1	
h sif	f->1	
h sin	 ->3	
h sis	t->3	
h sit	t->1	u->2	
h sju	k->1	
h sjä	l->3	
h sjö	f->1	n->1	
h ska	l->4	p->9	t->1	
h ski	l->1	
h sko	g->1	
h skr	o->1	
h sku	l->3	
h sky	d->2	l->2	
h skä	r->2	
h skö	n->1	t->3	
h sla	m->1	
h slu	s->1	t->19	
h slä	c->1	p->2	
h smu	t->1	
h små	,->1	
h sna	b->3	
h snå	r->1	
h soc	i->40	
h sol	i->2	
h som	 ->89	,->3	
h spa	r->1	
h spe	c->4	
h spr	i->2	å->2	
h sta	b->2	r->1	t->9	
h sti	m->1	
h sto	l->1	r->2	
h str	a->9	i->1	u->6	ä->2	å->1	
h stä	d->1	l->3	m->1	r->2	
h stå	 ->1	l->3	n->1	
h stö	d->13	r->1	
h suc	c->1	
h suv	e->4	
h sva	g->2	r->2	
h svå	g->1	r->7	
h syf	t->2	
h syn	l->1	
h syr	i->1	
h sys	s->11	t->1	
h säg	:->1	a->3	e->3	
h säk	e->12	
h sän	d->1	
h sär	s->11	
h sät	t->2	
h så 	a->3	l->4	m->1	s->4	v->9	
h såd	a->4	
h sål	e->2	
h sås	o->1	
h söd	r->1	
h sör	j->1	
h t.o	.->1	
h ta 	f->1	h->1	o->1	u->2	
h tac	k->6	
h tak	t->1	
h tal	a->3	m->1	
h tan	k->1	
h tar	 ->1	
h tas	 ->2	
h tek	n->2	
h tel	e->4	
h the	 ->1	
h tid	i->1	p->2	
h tig	g->1	
h til	l->52	
h tin	g->2	
h tis	d->1	
h tit	t->1	
h tjo	c->1	
h tjä	n->3	
h tog	 ->1	
h tol	e->2	k->1	
h top	p->1	
h tot	a->1	
h tra	g->1	n->8	
h tre	 ->1	d->1	
h tro	 ->1	l->1	r->1	t->2	
h trå	d->1	n->1	
h tun	g->1	
h tur	i->14	
h tus	e->2	
h två	 ->2	n->1	
h tyd	l->13	
h tyv	ä->1	
h täm	l->1	
h tän	k->1	
h täp	p->1	
h und	a->2	e->14	v->1	
h ung	d->5	e->1	
h uni	o->1	v->1	
h upp	b->1	e->3	f->5	h->1	l->3	m->4	r->5	s->2	
h uta	n->5	
h utb	i->4	
h ute	s->1	
h utf	o->2	
h utg	i->1	ö->3	
h uti	f->1	
h utl	ä->1	
h utn	y->2	
h uto	m->1	
h utr	i->2	
h uts	e->1	k->1	l->2	
h utt	a->2	ö->1	
h utv	e->22	i->1	ä->3	
h utö	v->1	
h vad	 ->10	
h val	b->1	f->1	t->1	u->10	
h van	 ->3	s->1	
h vap	e->3	
h var	 ->7	a->3	f->4	j->6	n->1	s->1	
h vek	h->1	
h vem	 ->2	
h ver	k->9	
h vet	e->10	t->1	
h vi 	a->4	b->13	d->1	f->9	g->2	h->15	i->1	k->9	l->2	m->10	r->1	s->5	t->2	u->3	v->7	ä->2	
h via	 ->1	
h vid	 ->4	g->1	t->1	
h vik	t->3	
h vil	k->9	l->4	
h vin	s->1	
h vis	 ->2	,->1	a->5	s->4	t->1	
h väd	j->1	
h väg	a->1	r->1	
h väl	 ->3	f->3	j->2	k->2	m->1	s->1	
h vän	l->1	s->1	
h väp	n->1	
h vär	d->3	l->1	
h väx	t->4	
h vål	d->1	
h vår	 ->4	a->4	t->3	
h vör	d->1	
h yng	s->1	
h yrk	e->1	
h ytl	i->1	
h ytt	e->3	r->1	
h ÖVP	 ->1	
h Öst	e->6	
h äga	n->1	
h ägn	a->1	
h än 	e->1	m->3	
h änd	a->1	r->2	å->2	
h änn	u->3	
h är 	b->1	e->3	k->2	n->1	o->1	r->1	
h äre	n->1	
h äve	n->31	
h å a	n->4	
h åkl	a->1	
h åsa	m->1	
h åsi	k->1	
h åst	a->1	
h åte	r->26	
h åtg	ä->3	
h öka	d->3	
h öms	e->1	
h öns	k->1	
h öpp	e->11	n->2	
h öre	g->1	
h öst	e->3	u->1	
h öve	r->16	
h övr	i->4	
h! Ur	s->1	
h)Det	 ->1	
h, at	t->1	
h, de	t->1	
h, fr	a->1	
h, fö	r->2	
h, he	r->1	
h, i 	a->1	
h, nå	g->1	
h, or	d->1	
h, re	n->1	
h, sl	u->1	
h, so	m->3	
h, tr	o->1	
h, ut	a->1	
h-Beh	r->7	
h-avt	a->1	
h.Det	 ->1	
h.Eft	e->1	
h.För	u->1	
h.Jag	 ->1	
h.Vi 	m->1	
h/ell	e->1	
h: Ve	m->1	
h?Fru	 ->1	
hI ok	t->1	
hII. 	f->1	
ha an	s->2	v->1	
ha ar	b->1	
ha at	t->1	
ha be	g->1	h->2	v->1	
ha br	u->1	
ha de	n->2	s->1	t->4	
ha di	s->1	
ha dr	u->1	
ha dö	t->1	
ha eg	n->1	
ha en	 ->36	
ha er	b->1	
ha et	t->17	
ha fr	a->1	i->2	
ha fu	n->1	
ha fö	r->2	
ha ge	n->2	
ha gj	o->2	
ha gr	ä->1	
ha ha	f->1	n->1	
ha hi	t->1	
ha hö	g->3	r->1	
ha i 	å->1	
ha in	 ->1	r->1	
ha kl	a->1	
ha ko	m->3	n->2	
ha ku	n->2	
ha kv	a->1	
ha kä	r->1	
ha ly	s->3	
ha lä	s->1	
ha ma	j->1	t->1	
ha me	d->2	
ha mi	n->1	
ha mo	d->2	
ha my	c->2	
ha mö	j->3	
ha ne	d->1	
ha ny	t->1	
ha nå	g->7	t->1	
ha oc	h->1	
ha of	f->1	
ha pr	e->1	o->1	
ha rä	t->2	
ha rå	d->1	
ha sa	g->1	m->2	t->1	
ha se	t->1	
ha sj	u->1	
ha sk	a->2	e->1	
ha st	o->1	u->2	
ha su	t->1	
ha sy	n->1	
ha ta	g->1	
ha ti	l->4	
ha tr	e->1	
ha tv	å->3	
ha ty	d->2	
ha un	d->2	
ha up	p->1	
ha ut	t->1	v->1	
ha va	r->7	
ha ve	l->1	
ha vi	s->3	
ha vä	g->1	r->1	v->1	
ha yt	t->1	
ha äg	t->1	
ha än	d->1	
ha ås	t->1	
ha ön	s->2	
ha öv	e->1	
ha, e	t->1	
ha.Al	l->1	
habil	i->1	
hablo	n->1	
hade 	a->4	b->5	d->1	e->3	f->7	g->4	h->3	i->4	j->2	k->9	m->3	n->2	o->2	p->2	r->2	s->6	t->5	v->17	ä->1	ö->2	
hade?	J->1	
haft 	a->3	b->1	d->1	e->3	f->5	i->1	m->4	n->2	o->1	p->2	s->6	t->2	u->1	v->1	ä->1	
haft,	 ->2	
haft.	V->1	
hagli	g->2	
hakat	 ->1	
hall"	,->1	
halt 	v->1	
halv 	d->1	t->2	
halva	 ->4	
halvh	j->1	
halvm	i->1	
halvo	f->1	
halvt	 ->2	i->3	
halvv	ä->2	
halvå	r->5	
halvö	,->1	.->1	n->1	
hambu	r->1	
hamel	s->1	
hamma	r->1	
hamn 	i->1	m->2	p->1	
hamn.	D->1	
hamna	 ->3	d->1	r->22	v->2	
hamnb	e->1	
hamne	n->2	
hamni	n->1	
hamnk	o->2	
hampa	g->1	
han a	n->3	r->1	t->1	v->1	
han b	e->3	
han d	r->1	å->1	
han e	l->1	
han f	ä->1	å->1	ö->3	
han g	e->1	j->1	ö->1	
han h	a->20	e->1	u->1	
han i	 ->5	b->1	n->8	
han j	u->2	
han k	a->1	o->6	
han l	a->4	ä->1	
han m	o->1	å->1	
han n	y->2	ä->1	
han o	c->2	r->1	
han p	r->1	å->2	
han s	a->3	i->2	k->3	t->1	v->1	ä->2	
han t	a->2	o->1	y->1	ä->1	
han u	t->3	
han v	i->6	
han ä	n->1	r->7	v->1	
han ö	n->1	
han, 	e->1	v->1	
han; 	J->1	
hand 	a->3	b->2	d->3	h->3	i->1	k->1	l->1	m->1	n->2	o->13	p->3	s->5	t->2	u->1	v->2	ä->4	
hand,	 ->4	
hand.	A->1	D->2	
hand?	F->1	
handa	 ->3	h->43	
hande	 ->1	l->29	n->6	
handf	u->1	
handi	c->1	k->3	
handl	a->165	i->182	ä->1	
hands	a->4	b->1	k->12	
handu	p->2	
hang 	b->1	e->1	f->2	g->2	h->1	j->1	k->1	m->1	o->2	s->4	ä->4	
hang,	 ->6	
hang.	.->1	D->4	J->1	O->1	Ä->1	
hange	n->2	t->11	
hanka	r->1	
hans 	a->10	b->11	e->5	f->15	g->1	h->1	i->4	k->7	l->2	o->2	p->5	r->1	s->6	u->9	v->2	å->1	
hanse	n->4	r->2	
hante	r->41	
hantv	e->2	
hapea	u->1	
happy	 ->1	
har -	 ->2	
har 1	3->1	7->1	
har 4	0->1	
har A	l->1	
har B	N->1	
har E	u->7	
har G	o->1	
har L	o->2	
har P	a->1	
har S	o->1	
har a	c->2	g->1	k->1	l->19	n->34	r->4	t->12	v->12	
har b	a->3	e->42	i->8	l->15	o->1	r->4	y->2	ä->1	ö->2	
har c	i->1	o->1	
har d	e->72	i->7	o->2	r->7	ä->7	å->1	ö->1	
har e	f->3	g->1	k->1	m->3	n->50	r->4	t->32	x->4	
har f	a->8	e->2	l->6	o->5	r->30	u->7	ä->1	å->28	ö->84	
har g	a->3	e->16	i->3	j->45	l->2	o->8	r->3	å->11	ö->1	
har h	a->19	e->7	i->8	o->1	ä->9	å->5	ö->12	
har i	 ->27	d->3	n->71	s->1	
har j	a->25	u->14	
har k	a->2	l->2	o->35	u->12	v->1	ä->1	ö->2	
har l	a->36	e->9	i->5	o->4	u->1	y->17	ä->12	å->3	ö->4	
har m	a->23	e->20	i->5	o->6	y->4	å->3	ö->6	
har n	a->2	i->2	o->4	u->13	y->3	ä->9	å->28	ö->2	
har o	b->1	c->18	f->4	l->2	m->3	r->2	
har p	a->4	e->3	l->1	r->9	å->20	
har r	a->4	e->27	y->1	ä->14	å->2	ö->5	
har s	a->34	e->13	i->4	j->3	k->24	l->4	m->1	o->3	p->6	t->28	v->1	y->1	ä->4	å->5	
har t	a->30	e->2	i->25	o->1	r->6	v->3	y->3	ä->2	
har u	n->14	p->22	t->18	
har v	a->31	e->9	i->87	u->1	ä->9	å->3	
har ä	g->4	n->13	r->2	v->2	
har å	l->1	s->1	t->2	
har ö	k->6	s->1	v->5	
har" 	m->1	
har, 	a->1	d->1	e->1	f->1	l->2	o->3	s->3	u->1	ä->1	
har.D	e->1	
har.T	a->1	
har: 	d->1	
har?N	i->1	
harad	e->1	
haras	 ->1	
hard 	C->1	
hard-	a->1	
harm 	e->4	
harm-	e->1	
harma	c->1	
harmo	n->18	
hartr	a->1	
has b	e->1	
hasta	d->1	r->1	t->1	
hasti	g->1	
hat o	c->1	
hatet	 ->1	,->1	
hatis	k->1	
hatte	n->1	
hauss	e->1	
hav f	ö->1	
hav o	c->1	
hav, 	o->1	
havan	d->1	
havar	e->1	n->2	
haven	 ->2	,->1	.->1	
haver	e->1	i->6	
havet	 ->10	,->1	.->3	s->2	
havs 	h->2	m->1	v->1	
havs,	 ->4	
havs.	A->1	D->1	R->1	V->1	
havs?	T->1	
havsf	o->1	ö->1	
havsl	ä->1	
havsm	i->2	
havso	m->1	
havsv	a->1	
he Ba	n->1	
he Ro	y->1	
he ci	v->1	
he im	p->1	
he oc	h->1	
he, L	i->1	
head-	k->1	
heato	 ->8	.->1	b->1	s->11	
hebre	i->1	
heck 	i->1	
heder	 ->1	s->1	v->1	
hedra	 ->2	d->1	n->1	r->1	
heer 	o->1	s->2	
heer,	 ->4	
heerJ	a->1	
heerb	e->3	
heers	 ->3	
hef h	a->1	
hefen	 ->1	
hefer	 ->4	,->2	.->1	n->8	
heik.	D->1	
heikh	 ->1	-->1	.->2	
hejda	s->1	t->1	
hekta	r->2	
hel b	e->1	
hel d	e->6	
hel k	v->1	
hel p	e->1	
hel r	a->1	ä->1	
hela 	9->1	B->1	E->19	M->1	a->1	b->2	d->17	e->3	f->7	g->3	h->2	i->3	k->7	l->1	m->1	o->1	r->3	s->5	t->11	u->8	v->5	å->3	
helge	n->1	
helhe	t->21	
helhj	ä->8	
helig	a->1	
hell 	o->1	s->1	
helle	r->47	
hellr	e->6	
helms	h->1	
helsi	k->1	
helst	 ->35	,->7	.->4	
helt 	a->4	b->1	d->1	e->24	f->5	g->2	h->2	i->8	k->23	l->2	m->3	n->4	o->24	p->2	r->11	s->6	t->3	u->2	v->2	ä->1	å->2	ö->3	
helt,	 ->1	
helt.	 ->1	D->1	E->1	
heltä	c->4	
hem e	f->1	
hem f	ö->1	
hem o	c->2	
hem t	i->1	
hem ä	r->1	
hem. 	H->1	
hem.N	i->1	
hema 	g->1	
hemby	g->1	
hemfö	r->1	
hemla	n->3	
hemli	g->5	
hemlä	n->1	x->1	
hemlö	s->5	
hemma	 ->7	,->1	p->1	
hemme	t->1	
hemsk	 ->1	a->4	
hemvi	s->1	
hen f	ö->3	
hen h	a->1	
hen i	 ->1	
hen s	j->1	
hen v	i->1	
hen, 	j->1	
hen.F	r->1	
hen; 	d->1	
henge	n->10	
henne	 ->7	.->1	s->19	
hens 	b->2	
hephe	r->3	
her i	n->1	
her o	c->1	
her v	e->1	
her" 	s->1	
heran	s->1	
herar	,->1	
herds	t->3	
heren	s->1	
hern 	f->3	s->1	t->1	
hern,	 ->3	
herna	 ->1	.->1	
heroi	s->1	
herr 	B->8	C->3	E->2	F->1	G->1	H->2	J->1	K->6	L->1	M->1	N->1	P->6	R->1	S->4	f->4	g->1	k->70	l->10	m->1	o->2	p->1	r->7	t->28	v->3	
herra	r->45	
hes i	 ->1	
het -	 ->1	
het 1	9->1	
het D	a->1	
het R	a->1	
het S	t->1	
het a	l->1	t->54	v->8	
het b	e->6	l->1	o->1	u->1	ö->1	
het d	e->9	o->1	ä->2	
het e	f->3	l->11	n->2	
het f	i->3	o->1	r->3	u->2	ö->48	
het g	e->3	
het h	a->5	e->1	o->1	ä->2	ö->1	
het i	 ->51	n->16	
het k	o->7	r->1	u->1	ä->1	
het l	a->1	i->2	
het m	e->61	i->1	o->3	å->5	
het n	a->1	ä->5	
het o	c->117	m->7	
het p	å->16	
het r	i->1	ä->1	ö->3	
het s	k->5	o->35	t->2	y->1	ä->3	å->3	
het t	i->15	ä->1	
het u	n->4	p->1	t->2	
het v	a->6	i->7	
het ä	g->1	r->16	v->2	
het å	r->1	t->7	
het!K	u->1	
het" 	(->1	g->1	m->1	
het, 	a->2	b->1	d->8	e->3	f->8	h->3	i->5	j->2	k->3	l->2	m->8	n->4	o->12	p->1	r->2	s->37	u->7	v->6	ä->1	ö->1	
het. 	D->2	E->1	M->1	
het.(	F->1	
het.A	t->1	v->1	
het.B	e->1	
het.D	e->23	ä->4	
het.E	n->2	t->1	u->2	
het.F	r->4	ö->4	
het.H	a->3	e->3	
het.I	 ->6	
het.J	a->12	
het.L	a->1	i->1	
het.M	a->2	e->5	
het.N	i->3	u->2	ä->1	
het.O	c->1	m->2	r->1	
het.P	a->1	å->1	
het.R	a->1	e->1	
het.S	o->2	t->1	å->1	
het.T	a->2	h->1	r->1	
het.V	a->1	i->8	ä->1	
het.Å	r->1	
het: 	F->1	
het; 	f->1	
het? 	R->1	
het?A	t->1	
het?K	o->1	
het?N	i->1	
het?S	k->1	
het?V	i->1	
hetJa	g->1	
heta 	i->1	
heten	 ->219	)->1	,->27	.->45	s->32	
heter	 ->222	,->31	.->37	?->1	n->111	s->2	
hetet	e->1	
hetli	g->36	
hets 	o->1	s->1	
hets-	 ->2	
hetsa	k->1	n->1	s->3	v->1	
hetsb	a->1	e->1	u->1	
hetsc	e->1	h->3	
hetse	n->4	
hetsf	l->15	r->8	å->1	ö->2	
hetsg	a->2	r->3	
hetsk	a->1	o->2	r->2	
hetsl	a->3	
hetsm	y->8	
hetsn	i->2	o->2	ä->1	
hetso	m->4	
hetsp	e->1	o->5	r->58	
hetsr	a->2	i->1	ä->1	å->18	
hetss	i->2	k->1	t->3	y->3	
hetst	i->5	ä->2	
hetsu	t->5	
hetsv	a->1	e->1	
hetså	t->2	
hett 	e->1	
hetta	.->1	
hette	 ->1	
heuge	n->2	
hez t	o->1	
hhofe	r->1	
hiel 	v->1	
hiera	r->4	
hies 	a->1	r->1	
high 	l->1	
hill 	o->1	
hinde	r->34	
hindr	a->49	e->3	
hingt	o->3	
hinna	 ->2	
hip m	e->1	
hiqui	t->1	
histi	s->2	
histo	r->34	
hit m	e->2	
hit o	c->1	
hit s	o->1	
hit, 	e->1	
hitta	 ->12	d->1	r->3	t->1	
hitti	l->41	
hjamo	,->1	
hjäl 	d->1	
hjälp	 ->48	,->2	.->5	a->41	e->5	l->1	s->1	t->3	v->1	
hjärt	a->20	l->7	
hler 	t->1	
hler,	 ->1	
hler.	F->1	
hlers	 ->1	
hne, 	d->1	
hner 	f->1	k->1	u->1	
hner,	 ->3	
hners	 ->6	
ho fö	r->1	
ho på	p->1	
ho so	m->1	
ho vä	l->1	
ho. D	e->1	
hobby	,->1	b->1	
hoc-d	i->1	
hoc-t	r->1	
hock 	f->1	
hocka	d->1	
hocke	r->2	
hoek 	s->1	
hofer	,->1	
hokla	d->1	
hol, 	t->1	
holka	 ->2	s->2	
holm 	d->1	
holm,	 ->1	
holm.	H->1	
hom P	o->3	
homof	o->1	
homog	e->2	
homos	e->1	
hon a	l->1	
hon f	o->1	ö->3	
hon h	a->4	
hon i	 ->1	n->3	
hon j	u->1	
hon k	a->1	o->1	
hon l	a->1	
hon p	å->2	
hon s	e->1	k->3	
hon t	a->1	i->1	
hon u	n->1	
hon v	i->1	
hon ä	r->2	
honom	 ->22	,->2	.->4	
hop a	l->1	
hop d	e->1	
hop f	ö->1	
hop p	e->1	
hop s	i->1	
hop t	i->1	
hop u	t->1	
hop ä	n->1	
hop, 	e->1	o->1	
hop.D	e->1	
hop.I	n->1	
hop.J	a->1	
hopp 	f->1	
hoppa	 ->1	d->1	s->95	
hoppe	t->1	
hoppl	ö->1	
hoppn	i->12	
hord 	k->1	
horde	r->1	
horis	o->3	
hormo	n->1	
hos D	a->1	
hos E	G->1	u->1	
hos F	P->1	
hos R	E->1	
hos a	l->2	v->1	
hos b	e->1	l->1	
hos d	e->12	
hos e	n->2	
hos f	a->1	ö->2	
hos i	n->1	
hos k	o->6	
hos m	e->2	ä->1	å->1	
hos o	r->1	s->3	
hos p	r->2	
hos r	å->1	
hos s	i->2	
hos t	i->1	
hos v	u->1	å->1	
hospi	c->1	
hot -	 ->1	
hot f	r->1	
hot m	o->6	
hot o	m->1	
hot p	å->1	
hot s	p->1	
hota 	f->1	
hotad	.->2	e->4	
hotan	d->1	
hotar	 ->6	
hotas	 ->3	.->1	
hotat	 ->1	
hotbi	l->1	
hotel	s->1	
hotet	 ->7	
hotfu	l->1	
hov a	v->15	
hov i	 ->1	
hov k	o->1	
hov o	c->4	
hov s	o->1	y->1	
hov t	i->8	
hov, 	a->1	n->1	
hov.A	v->1	
hov.H	e->1	
hov.U	p->1	
hoven	 ->4	.->1	
hovet	 ->34	
hovsm	a->2	ä->3	
how t	i->1	
hrend	t->7	
hreye	r->3	
hrkop	 ->1	
hroed	t->14	
hröde	r->1	
hs i 	o->1	
ht ka	n->1	
ht me	d->1	
ht oc	h->1	
ht ti	l->1	
ht.De	n->1	
htala	t->1	
hters	k->2	
htför	d->3	
htid 	i->1	
hts.A	n->1	
hu oc	h->1	
hud B	a->2	
hugg 	p->3	
hulda	 ->1	
hulz 	e->1	s->2	
human	 ->1	i->5	
humle	n->1	
humör	 ->2	
hun s	a->1	
hund.	N->1	
hundr	a->19	
hur E	G->1	u->1	
hur a	l->1	n->2	r->1	v->1	
hur b	e->2	i->1	r->3	u->1	
hur d	e->41	i->1	
hur e	n->2	t->1	
hur f	a->1	o->1	r->1	ö->2	
hur g	o->1	å->1	
hur h	a->2	o->1	ö->1	
hur i	n->1	
hur k	l->3	o->7	ä->1	
hur l	e->1	i->1	ä->2	å->5	
hur m	a->18	e->1	i->1	ä->1	å->3	
hur n	i->3	u->2	
hur o	c->1	f->1	
hur p	a->3	e->1	r->2	
hur r	i->1	
hur s	a->1	k->4	m->1	n->1	o->4	t->10	v->4	ä->1	
hur t	i->1	r->1	u->1	
hur u	n->2	p->1	r->1	t->3	
hur v	i->28	ä->2	å->1	
hur.K	o->1	
hur.R	å->1	
huruv	i->14	
hus 1	9->1	
hus h	a->1	
hus o	c->2	
hus s	o->1	
hus u	n->1	
hus, 	e->1	f->1	h->1	m->2	
hus.E	u->1	
hus.G	e->1	
hus.H	e->1	
husef	f->3	
huset	 ->3	
husga	s->4	
hushå	l->1	
huslä	k->1	
husöv	e->1	
huvud	 ->9	a->5	d->2	e->1	f->4	l->1	r->3	s->21	u->1	
hwarz	w->1	
hweiz	,->1	
hwitz	.->1	
hy oc	h->1	
hyckl	a->2	e->3	
hygie	n->2	
hylla	n->1	
hylln	i->1	
hypot	e->2	
hyrd 	a->1	
hyreg	i->1	
hysa 	f->1	m->1	ä->1	
hyser	 ->5	
hysse	n->5	
hyste	r->1	
häfta	t->1	
häfti	g->1	
häler	i->1	
hälft	e->3	
hälle	 ->10	n->5	s->2	t->25	
hälli	g->32	
hälls	e->3	m->1	o->1	s->1	v->1	
hälsa	 ->15	,->3	.->1	n->4	r->1	
hälsn	i->2	
hälso	-->1	e->1	r->2	s->1	v->3	
hämma	d->1	n->2	r->1	
hämna	s->1	
hämni	n->1	
hämta	 ->3	n->1	r->1	s->1	t->1	
hämtn	i->1	
hän; 	d->1	
hända	 ->16	.->1	?->1	
hände	 ->7	.->1	l->25	r->28	
hänfö	r->1	
hänga	 ->1	n->2	r->3	
hängb	r->1	
hänge	r->12	t->1	
hängi	g->2	
hänse	e->8	
hänsy	n->72	
hänt 	a->2	t->1	u->2	
hänt.	V->1	
hänt:	 ->1	
hänta	.->1	
hänvi	s->35	
här -	 ->6	
här D	o->1	
här a	k->1	l->1	n->2	t->1	v->1	
här b	e->6	l->1	u->1	ö->1	
här c	i->1	
här d	e->8	i->1	
här e	n->2	t->1	
här f	a->10	i->2	o->1	r->18	ö->10	
här g	å->4	
här h	a->6	
här i	 ->45	d->1	n->13	
här k	a->3	o->4	v->1	
här l	a->2	i->1	å->2	
här m	a->1	ä->1	å->1	
här n	y->1	ä->1	
här o	c->6	l->1	m->7	
här p	a->3	e->1	l->3	o->1	r->5	u->2	å->1	
här r	e->3	u->1	ö->1	
här s	a->3	i->3	k->1	l->2	n->2	o->3	t->1	v->1	ä->2	
här t	e->2	i->2	y->11	
här u	n->2	p->2	t->1	
här v	e->4	i->6	ä->1	
här y	p->1	t->1	
här ä	r->8	
här å	r->2	
här ö	v->2	
här, 	a->3	d->2	f->1	i->1	m->4	n->1	o->1	u->1	
här. 	i->1	
här.D	e->3	
här.E	f->1	
här.F	ö->1	
här.K	o->1	
här.V	i->3	
här; 	v->1	
här?D	e->1	
härda	 ->1	r->1	
härdi	g->1	
härdl	i->3	
häref	t->1	
härig	e->2	
härja	d->2	
härle	d->1	
härme	d->3	
härrö	r->4	
härti	l->1	
härvi	d->1	
häste	n->1	
häva 	a->1	i->1	s->1	
hävas	 ->4	
hävda	 ->7	d->3	r->12	t->5	
hävdv	u->1	
häver	 ->1	
hävs.	E->2	
hävts	.->1	
håg I	r->1	
håg a	t->8	
håg d	e->3	
håg r	e->1	
håg s	i->1	
håg ä	r->1	
håg.E	u->1	
hågor	 ->1	?->1	
hål i	 ->2	
hål, 	s->1	
hål: 	V->1	
hålen	 ->1	
håll 	a->1	f->2	h->1	i->3	k->2	o->3	r->1	s->4	t->1	v->1	
håll,	 ->5	
håll.	D->2	F->1	I->1	J->2	V->1	
håll:	 ->1	
håll?	.->1	
hålla	 ->85	,->1	n->84	s->11	
hållb	a->25	
hålle	n->1	r->93	t->27	
hålli	t->23	
hålln	a->1	i->66	
hålls	 ->4	,->1	.->1	a->2	l->2	m->2	r->2	t->7	v->1	
hån m	o->1	
hånar	 ->1	
hård 	g->1	k->1	p->1	
hård,	 ->1	
hårda	 ->7	r->3	s->2	
hårdn	a->2	
håret	 ->1	
hårkl	y->1	
hårt 	a->3	d->2	l->1	r->1	
hårt,	 ->1	
hårt.	M->1	
håvar	 ->1	
hône-	A->1	
hög a	r->1	
hög b	e->1	
hög f	e->1	
hög g	r->6	
hög i	n->1	
hög k	v->1	
hög n	i->2	
hög p	r->2	
hög s	e->1	k->1	o->1	t->2	y->1	
hög, 	d->1	
höga 	f->1	g->1	k->3	n->1	p->1	r->2	s->1	t->2	å->2	
höga,	 ->1	
höga.	M->1	
högak	t->1	
höge 	k->1	r->1	
höger	 ->2	,->1	e->5	m->1	n->19	p->1	v->1	
höghe	t->2	
höglj	u->1	
högni	v->3	
högra	 ->1	
högre	 ->18	.->1	
högsk	o->1	
högst	 ->11	,->1	a->16	
högt 	f->1	i->2	p->3	s->1	u->1	v->1	
högt,	 ->1	
högt.	S->1	
högte	k->2	
högti	d->4	
höja 	J->1	d->1	f->1	l->1	
höjan	d->1	
höjas	.->1	
höjd 	-->1	a->1	g->1	s->1	u->1	
höjde	 ->1	n->1	r->3	
höjdp	u->2	
höjer	 ->1	
höjni	n->2	
höjs 	t->1	
höjts	 ->1	
höll 	K->1	a->3	d->1	e->4	i->1	m->1	n->1	s->1	ö->1	
hölls	 ->4	
höna 	h->1	
hör a	l->1	t->5	
hör b	l->1	
hör d	e->1	ä->1	
hör e	n->2	t->1	
hör f	r->1	
hör h	e->5	ä->1	
hör i	h->2	n->2	
hör j	a->1	
hör n	u->1	å->2	
hör s	a->1	ä->1	
hör t	i->7	
hör v	i->2	
hör. 	E->1	
höra 	a->5	d->2	e->1	f->1	k->1	m->2	n->2	o->2	p->4	t->1	v->3	
höra,	 ->1	
höra.	D->1	E->1	
höran	d->2	
hörar	l->1	
höras	 ->1	,->1	
hörd 	k->1	m->1	
hörd.	D->1	
hörda	 ->1	
hörde	 ->4	
hörig	 ->2	a->2	h->15	
hörli	n->1	
hörn 	d->1	f->1	
hörns	t->1	
hört 	-->1	D->1	d->2	e->3	f->2	i->2	m->3	o->1	p->2	s->3	t->2	u->1	v->1	
hört,	 ->1	
hört.	J->1	
hörts	 ->1	
höst 	p->1	
höva 	a->1	e->1	f->1	g->3	k->2	l->1	p->2	r->1	u->2	ö->1	
hövas	.->1	
hövde	 ->2	
höver	 ->96	,->1	.->2	
hövli	g->1	
hövs 	d->3	e->6	f->2	i->3	m->1	n->1	o->1	p->1	s->2	
hövs,	 ->2	
hövs.	D->1	F->1	I->1	S->2	
hövt 	s->1	t->1	
hövts	 ->1	
hüsse	l->4	
i "ge	n->1	
i - C	a->1	
i - a	t->1	v->2	
i - d	e->1	
i - e	n->1	
i - j	a->1	
i - n	ä->1	
i - r	å->1	
i - s	o->1	
i - v	ä->1	
i 15 	s->1	
i 196	7->1	
i 199	3->1	5->1	7->3	8->2	9->7	
i 20 	å->1	
i 200	 ->2	0->8	2->2	
i 55 	m->1	
i 8 b	e->1	
i 8 o	c->1	
i ABB	-->1	
i Ada	n->1	
i Adr	i->1	
i Afr	i->3	
i Akk	u->1	ö->1	
i Als	a->1	
i Ams	t->17	
i Asi	e->1	
i Auv	e->1	
i Avi	a->1	
i BNI	 ->1	
i Bel	g->2	
i Ber	e->1	g->1	l->7	
i Bis	c->5	
i Bor	d->1	
i Bra	n->2	
i Bre	t->2	
i Bry	s->7	
i Bud	a->1	
i CEN	:->1	
i Cav	a->1	
i Cen	t->5	
i Cer	m->1	
i Cus	í->1	
i DDR	.->1	
i Dan	m->9	
i Dub	l->4	
i ECH	O->1	
i EG-	d->1	f->7	
i EKS	G->3	
i EMU	-->1	
i EU 	m->1	o->1	
i EU,	 ->1	
i EU-	b->1	f->2	l->2	
i EU:	s->7	
i Eko	f->1	
i Eti	o->1	
i Eur	o->173	
i Fac	t->1	
i Fei	r->1	
i Fin	l->2	
i Fol	k->1	
i Fra	n->11	
i För	b->2	e->12	
i GUE	/->1	
i Gaz	a->2	
i Gen	è->2	
i Gol	a->2	
i Gre	k->2	
i Gru	p->2	
i Gua	t->1	
i Gul	f->1	
i Hai	d->1	
i Hel	s->14	
i ICE	S->2	
i Ind	i->1	
i Int	e->1	
i Irl	a->10	
i Isr	a->1	
i Ist	a->1	
i Ita	l->6	
i Jon	c->1	
i Kar	l->1	
i Kau	k->2	
i Kfo	r->1	
i Kin	a->3	
i Kos	o->34	
i Kou	c->1	
i Kyo	t->1	
i Kär	n->1	
i Köl	n->1	
i Lam	a->7	
i Lan	g->1	k->3	
i Lap	p->2	
i Lea	d->1	
i Lib	y->1	
i Lii	k->2	
i Lil	l->1	
i Lis	s->5	
i Lom	é->1	
i Lon	d->4	
i Lor	r->1	
i Lut	t->1	
i Lux	e->4	
i Maa	s->2	
i Mac	a->1	
i Mad	r->2	
i McN	a->1	
i Med	e->1	
i Mel	l->14	
i Mex	i->1	
i Mit	r->1	
i Mon	t->2	
i Mos	k->1	
i Ned	e->4	
i New	 ->1	
i Nor	g->1	
i OLA	F->1	
i Oma	g->1	
i PPE	 ->1	-->2	
i Pad	d->1	
i Par	i->1	
i Pay	s->1	
i Pek	i->1	
i Por	t->5	
i Pro	d->1	
i Rap	k->1	
i Rom	-->1	
i Rys	s->2	
i Sai	n->1	
i San	 ->1	t->1	
i Sch	e->1	r->1	w->2	
i Sea	t->3	
i Sha	r->1	
i She	p->3	
i Sko	t->2	
i Sri	 ->3	
i Sto	c->2	r->9	
i Str	a->4	
i Sve	r->2	
i Syd	a->1	o->1	
i Syr	i->2	
i TV-	p->1	
i Tad	z->2	
i Tam	m->14	
i Tau	e->1	
i Tex	a->1	
i The	a->4	
i Thy	s->1	
i Tib	e->5	
i Tur	k->7	
i Tys	k->5	
i UEN	-->1	
i USA	 ->2	,->1	
i Urb	a->1	
i Van	 ->1	
i Vat	a->1	
i Ven	e->1	
i Vär	l->1	
i Wal	e->3	
i Was	h->1	
i Wie	n->1	
i Yas	s->1	
i a) 	b->1	
i abs	o->4	
i acc	e->2	
i age	r->3	
i aid	s->1	
i akt	 ->4	u->1	
i ald	r->1	
i all	 ->3	a->64	e->1	m->10	r->1	s->1	t->14	v->1	
i ana	 ->1	l->2	
i and	r->15	
i anl	e->1	
i ann	a->5	
i anp	a->1	
i ans	e->29	l->4	p->2	v->3	å->3	
i ant	a->1	
i anv	ä->13	
i arb	e->29	
i art	i->14	o->1	
i att	 ->78	
i avf	a->1	
i avg	e->4	ö->1	
i avh	ä->1	
i avl	a->1	
i avs	i->2	k->1	l->2	n->1	t->2	
i avt	a->2	
i avv	a->4	i->2	
i bal	a->1	
i bar	a->5	
i beb	å->1	
i bed	r->1	ö->3	
i bef	i->11	
i beg	r->4	
i beh	a->4	o->3	ö->48	
i bek	l->3	r->2	ä->1	
i ben	ä->1	
i ber	 ->3	e->2	ä->2	ö->3	
i bes	l->11	t->2	v->2	
i bet	a->2	e->1	o->3	r->2	v->1	y->1	ä->14	
i bev	i->2	
i bib	e->1	
i bid	r->3	
i bil	-->1	a->5	d->2	e->1	i->2	p->1	
i bio	s->2	
i bla	n->1	
i ble	v->1	
i bli	r->5	
i bok	s->1	
i bor	d->10	t->1	
i bra	 ->1	
i bri	s->1	
i bro	t->1	
i bru	k->2	
i bry	t->1	
i brä	s->1	
i brå	d->1	
i bud	g->9	
i byg	g->1	
i bät	t->2	
i båd	a->2	e->1	
i böc	k->1	
i bör	 ->32	,->1	.->1	j->9	
i cen	t->2	
i cir	k->1	
i dag	 ->109	,->25	.->22	:->1	e->5	l->1	o->2	s->1	
i dan	s->1	
i dat	a->1	
i de 	1->1	2->3	a->4	b->2	c->1	d->1	e->8	f->13	g->3	h->3	i->1	j->1	k->2	l->3	m->5	n->3	o->10	p->3	r->6	s->1	t->1	u->2	y->1	ö->3	
i deb	a->10	
i dec	e->7	
i del	a->2	s->1	t->2	
i dem	 ->1	.->1	o->2	
i den	 ->106	.->1	n->103	
i der	a->1	
i des	s->28	
i det	 ->106	,->3	.->3	a->5	t->97	
i dia	l->2	
i dir	e->16	
i dis	c->1	k->22	
i doc	k->1	
i dok	u->1	
i dom	i->1	s->3	
i dra	r->1	
i dri	c->1	f->1	
i där	e->1	f->3	i->1	m->2	
i då 	2->1	a->1	g->1	o->3	t->1	v->1	ä->1	
i eff	e->3	
i eft	e->13	
i ege	n->14	t->1	
i eko	n->6	
i eme	l->5	
i en 	a->16	b->3	d->7	e->9	f->6	h->3	i->1	k->6	l->4	m->17	n->3	o->2	p->10	r->11	s->16	t->3	u->3	v->6	å->2	
i ena	s->1	
i enh	ä->1	
i eni	g->1	
i enk	l->1	
i enl	i->28	
i ens	t->1	
i er 	s->1	u->1	v->2	
i era	 ->4	
i erb	j->1	
i erf	a->1	
i erk	ä->3	
i ert	 ->7	
i ett	 ->82	
i eur	o->6	
i eve	n->1	
i exa	k->1	
i exp	a->1	e->1	
i f.d	.->1	
i fak	t->6	
i fal	l->3	
i far	a->1	m->1	t->2	
i fas	t->4	
i fat	t->5	
i feb	r->7	
i fem	 ->2	t->1	
i fic	k->4	
i fin	a->1	n->2	
i fjo	l->2	
i fle	r->6	x->1	
i fok	u->1	
i fol	k->4	
i for	m->12	s->3	t->26	
i fra	m->62	
i fre	d->8	
i fri	h->1	
i fro	n->1	
i frä	m->1	
i frå	g->76	n->5	
i ful	l->4	
i fun	d->1	k->1	
i fyr	a->2	
i fär	d->2	s->1	
i fäs	t->1	
i få 	b->1	t->2	v->1	
i får	 ->23	,->1	
i fåt	t->5	
i föl	j->3	
i för	 ->31	b->16	d->40	e->18	f->7	g->3	h->25	k->3	l->6	m->3	o->3	p->1	r->11	s->46	t->1	v->17	
i gan	s->1	
i gar	a->2	
i ge 	a->1	e->1	k->1	u->1	
i gem	e->14	
i gen	a->1	d->1	e->1	g->1	o->13	
i ger	 ->7	
i gic	k->1	
i gjo	r->6	
i gla	d->1	s->1	
i glä	d->2	
i glö	m->1	
i god	 ->7	k->5	t->1	
i got	t->1	
i gra	t->2	
i gru	n->9	
i gäl	l->1	
i gär	n->2	
i gån	g->6	
i går	 ->13	,->2	.->2	
i gör	 ->18	.->1	a->6	s->1	
i ha 	e->2	t->1	u->1	ö->1	
i had	e->11	
i haf	t->3	
i ham	n->6	
i han	 ->1	d->6	s->7	t->2	
i har	 ->239	,->3	m->1	
i hav	 ->1	e->5	s->1	
i hel	a->20	g->1	h->3	t->5	
i hem	m->2	
i hen	n->1	
i her	r->1	
i hie	r->1	
i his	t->1	
i hit	t->5	
i hjä	l->1	r->2	
i hop	p->10	
i huv	u->7	
i hys	e->1	
i hän	d->9	s->1	v->2	
i här	 ->13	
i häv	d->2	
i hål	l->10	
i hån	a->1	
i hår	e->1	
i hög	 ->3	n->2	r->2	s->1	
i höl	l->1	
i hör	t->1	
i hös	t->1	
i i E	U->1	u->3	
i i G	U->1	r->1	
i i I	t->1	
i i L	i->1	
i i M	o->1	
i i P	P->1	
i i S	t->1	
i i T	u->1	
i i a	l->1	
i i d	a->13	e->11	
i i e	f->1	g->1	n->3	
i i f	r->1	
i i g	å->1	
i i j	u->1	
i i k	a->3	r->1	
i i m	e->1	o->5	y->1	
i i o	c->1	
i i p	a->2	
i i s	j->2	l->1	t->4	y->1	å->1	
i i t	r->1	
i i v	å->3	
i i Ö	s->1	
i i å	r->1	
i iak	t->1	
i ibl	a->2	
i ick	e->2	
i ige	n->1	
i igå	n->1	
i inb	e->1	
i ind	u->1	
i inf	o->1	r->1	ö->3	
i ing	e->4	i->1	å->3	
i inh	ä->1	
i ini	t->1	
i ink	o->2	
i inl	e->9	ä->2	
i inn	a->1	e->1	
i ino	m->2	
i inr	i->1	ä->1	
i ins	e->11	i->1	k->1	t->5	
i int	e->116	
i inv	a->1	
i ita	l->1	
i jag	a->1	
i jan	u->1	
i jor	d->1	
i ju 	o->2	v->1	
i jul	i->5	
i jun	i->6	
i jus	t->12	
i jäm	f->1	s->2	
i kab	i->1	
i kal	l->2	
i kam	m->19	p->2	
i kan	 ->90	,->1	d->1	s->5	
i kap	i->2	p->1	
i kat	o->1	
i ked	j->1	
i kla	r->7	v->1	
i kni	p->1	
i kny	t->1	
i koa	l->1	
i kom	 ->1	m->95	p->1	
i kon	c->3	f->2	k->10	s->7	t->3	v->2	
i kos	t->1	
i kra	f->24	
i kri	g->1	s->1	t->1	
i kry	p->1	
i krä	v->11	
i kul	i->1	t->1	
i kun	d->2	n->7	
i kur	s->2	
i kva	r->1	
i kvä	l->4	
i kän	n->13	
i lad	e->2	
i lag	.->1	e->1	s->9	t->2	
i lan	d->6	
i led	a->1	e->1	n->1	
i lev	a->1	t->1	
i lib	e->1	
i lid	e->1	
i lik	a->2	g->1	h->9	
i lin	j->5	
i lit	a->5	
i liv	e->1	
i lju	s->5	
i lov	a->2	
i lyc	k->3	
i lys	s->3	
i läg	g->8	
i läm	n->2	
i län	d->1	
i lär	d->1	
i lät	 ->1	t->1	
i låt	 ->1	a->1	e->1	
i löp	e->1	
i lös	g->1	
i maj	 ->2	,->1	.->2	
i mak	r->1	
i man	d->1	t->1	
i mar	k->2	s->1	
i mas	s->1	
i med	 ->23	b->4	d->1	g->2	i->1	l->31	v->2	
i mel	l->2	
i men	a->8	
i mer	 ->5	a->2	
i mig	 ->2	
i mil	j->6	
i min	 ->11	a->2	d->3	i->4	n->2	o->1	
i mis	s->2	
i mit	t->18	
i mju	k->1	
i mod	e->1	
i mor	g->32	
i mot	 ->3	i->1	s->8	t->1	
i myc	k->7	
i myn	d->1	
i män	n->1	
i mål	 ->5	-->1	
i mån	a->1	d->2	g->14	
i mås	t->145	
i möb	l->1	
i möj	l->3	
i nat	i->2	u->5	
i niv	å->4	
i nor	r->2	
i nov	e->5	
i nu 	b->1	d->3	e->1	g->3	h->4	i->1	k->2	m->3	r->1	s->1	t->1	v->1	ä->1	
i nul	ä->1	
i nya	 ->1	
i nyh	e->1	
i nyl	i->2	
i näm	n->7	
i när	 ->8	a->1	h->4	i->1	m->3	
i näs	t->1	
i nå 	å->1	
i någ	o->10	r->3	
i nöd	e->1	v->1	
i nöj	d->1	
i obj	e->1	
i obl	i->1	
i och	 ->70	
i ock	s->30	
i off	e->3	r->1	
i oft	a->1	
i ofö	r->1	
i okt	o->2	
i oli	k->4	
i olj	e->1	
i oly	c->1	
i om 	a->1	d->1	e->1	h->1	n->1	s->1	
i omf	o->1	
i omr	å->16	ö->1	
i ons	d->1	
i ord	 ->4	a->1	f->2	
i oro	a->2	
i oss	 ->10	
i oty	d->1	
i oun	d->1	
i oöv	e->1	
i par	l->40	
i pek	a->1	
i pen	g->1	
i per	i->3	
i pla	c->1	n->4	s->1	
i ple	n->4	
i plå	n->1	
i plö	t->1	
i pol	i->6	
i por	t->2	
i pos	i->2	
i pra	k->10	
i pre	c->1	j->1	s->4	
i pri	n->12	
i pro	b->2	c->3	g->4	j->1	p->2	t->3	
i pun	k->2	
i på 	I->1	a->1	b->1	d->2	e->2	l->2	m->1	n->2	t->1	v->1	
i påb	ö->1	
i pås	t->1	
i rad	e->1	i->1	
i ram	p->1	
i rap	p->8	
i rat	i->2	
i rea	g->1	l->5	
i red	a->11	
i ref	o->2	
i reg	e->6	i->12	l->3	
i rel	a->2	
i res	o->4	p->6	u->1	
i ret	o->1	
i rik	t->6	
i rim	l->1	
i rin	g->1	
i ris	k->1	
i rop	a->1	
i rul	l->1	
i rus	a->2	
i räk	n->4	
i rät	t->12	
i råd	e->35	
i rör	l->8	
i rös	t->8	
i sad	e->13	
i sak	e->2	
i sam	a->8	b->35	f->1	h->2	m->9	t->5	
i sat	t->1	
i se 	a->1	i->2	r->1	t->6	u->1	v->1	
i sen	a->2	
i sep	t->12	
i ser	 ->15	
i sex	 ->1	
i sid	o->1	
i sig	 ->16	.->2	;->1	
i sik	t->3	
i sin	 ->40	a->15	o->1	
i sis	t->2	
i sit	t->21	u->3	
i sju	 ->1	k->1	
i sjä	l->28	
i ska	 ->1	l->69	p->4	
i ske	p->1	
i ski	c->3	
i sko	g->2	
i skr	e->2	
i sku	g->1	l->21	
i sky	d->1	h->1	n->1	
i sli	p->2	
i slu	t->21	
i slö	s->1	
i små	 ->1	f->1	
i sna	b->2	r->9	
i soc	i->6	
i sol	i->1	
i som	 ->37	l->1	
i sor	g->1	
i spe	l->2	
i spä	n->1	
i sta	r->4	t->1	
i ste	r->1	
i sti	c->1	l->1	
i sto	r->12	
i str	a->1	i->9	u->1	ä->2	
i sty	r->2	
i stä	d->6	l->48	n->4	r->1	v->1	
i stå	n->4	r->7	
i stö	d->14	r->13	
i sub	v->1	
i sva	n->1	r->2	
i sve	n->1	
i svå	r->2	
i syd	v->1	
i syf	t->8	
i sym	p->1	
i syn	l->1	n->45	
i sys	s->4	t->1	
i säg	e->9	
i säk	e->4	
i säm	r->1	s->1	
i sän	d->1	
i sär	s->2	
i sät	t->2	
i så 	a->3	f->2	m->1	s->3	
i såd	a->7	
i såg	 ->1	
i sål	e->1	
i såv	ä->1	
i söd	r->1	
i t.e	x->2	
i ta 	d->1	h->1	
i tac	k->3	
i tag	i->3	
i tak	t->3	
i tal	a->20	m->1	
i tan	k->2	
i tar	 ->11	
i tem	p->1	
i tex	t->1	
i tid	 ->3	.->1	e->5	i->3	n->2	
i til	l->28	
i tit	t->1	
i tjä	n->1	
i tol	k->3	
i top	p->3	
i tor	n->1	
i tra	f->3	n->1	
i tre	 ->2	d->3	
i tro	d->1	l->1	r->6	t->1	
i trä	f->1	n->1	
i trå	d->1	
i tve	k->2	
i tvi	v->1	
i tvu	n->3	
i tvä	r->1	
i två	 ->5	
i tyc	k->7	
i tyd	l->1	
i tys	k->1	
i tyv	ä->2	
i tän	k->6	
i tät	e->2	
i und	e->11	r->1	v->1	
i ung	e->1	
i uni	o->31	
i upp	 ->3	d->3	e->1	l->3	m->7	n->7	r->4	s->3	
i ur 	k->1	
i urs	p->1	
i urv	a->1	
i uta	n->3	
i utb	y->2	
i ute	s->1	
i utf	o->3	ö->1	
i utg	ö->1	
i utk	a->1	
i utl	a->1	å->1	
i utn	ä->1	
i uto	m->1	
i uts	k->24	t->1	
i utt	a->2	r->2	
i utv	e->8	i->2	ä->1	
i utö	v->1	
i vac	k->1	
i vad	 ->3	
i vak	s->1	
i val	u->1	
i van	 ->5	l->1	
i var	 ->8	a->8	d->1	j->14	k->2	m->1	n->2	t->1	
i vec	k->1	
i vel	a->1	
i vem	s->1	
i ver	k->18	
i vet	 ->28	,->7	a->2	e->1	
i vid	 ->2	t->2	
i vik	t->1	
i vil	j->2	k->17	l->66	
i vin	d->1	
i vis	a->4	s->23	
i vit	b->13	
i väg	e->3	
i väl	d->1	f->1	j->1	k->4	
i vän	d->3	l->1	s->1	t->9	
i vär	l->12	
i väs	e->1	
i våg	a->1	
i vår	 ->22	a->20	t->22	
i yrk	e->2	
i ytt	e->2	r->1	
i zon	 ->1	e->1	
i ÖVP	 ->1	
i Öst	e->37	
i äga	n->1	
i ägn	a->4	
i äkt	e->1	
i ämn	e->3	
i än 	e->1	
i änd	r->10	å->3	
i änn	u->6	
i är 	a->5	b->7	d->5	e->4	f->4	h->1	i->9	j->1	k->1	m->11	n->4	o->2	p->1	s->5	t->2	u->1	v->2	ä->1	ö->5	
i äre	n->1	
i äve	n->6	
i ålä	g->1	
i år 	2->1	k->1	u->1	v->1	
i år,	 ->3	
i år.	D->1	F->1	H->1	K->1	
i åra	t->1	
i årt	i->1	
i åst	a->1	
i åta	n->1	
i åte	r->7	
i åtg	ä->1	
i åtm	i->1	
i öka	r->1	
i öns	k->7	
i öpp	e->1	
i öre	g->1	
i öst	 ->1	e->1	r->1	
i öve	r->17	
i övr	i->5	
i! Ja	g->1	
i! Jo	n->1	
i! Up	p->1	
i!Her	r->1	
i!Jag	 ->1	
i" so	m->1	
i, Mi	t->1	
i, be	t->1	
i, br	i->1	
i, de	 ->2	n->1	t->2	
i, då	l->1	
i, ef	t->1	
i, en	 ->3	
i, fr	u->3	
i, fö	r->1	
i, gi	v->1	
i, he	r->4	
i, in	o->1	t->1	
i, ja	 ->1	g->1	
i, ju	s->1	
i, ka	n->2	
i, ku	l->1	
i, la	n->1	
i, li	k->3	
i, lj	u->1	
i, me	d->3	n->6	
i, mi	n->1	s->1	
i, ne	p->1	
i, nä	r->1	
i, ob	e->1	
i, oc	h->7	
i, om	 ->2	
i, or	d->1	
i, pr	e->1	
i, se	d->1	
i, si	s->1	
i, sk	r->1	u->1	
i, so	m->5	
i, så	 ->1	s->1	
i, t.	e->2	
i, ti	l->1	
i, tr	o->1	
i, ut	r->1	v->1	
i, va	d->1	
i, vi	c->1	l->1	
i, än	d->1	
i, är	 ->1	
i, äv	e->2	
i- oc	h->10	
i-, t	r->1	
i-gem	e->1	
i-irl	ä->1	
i-ras	i->1	
i.(Pa	r->1	
i.. (	F->1	
i...(	T->1	
i.All	a->1	t->1	
i.Anl	e->1	
i.Båd	a->1	
i.De 	p->1	
i.Den	 ->2	
i.Det	 ->8	
i.Där	f->1	
i.Eft	e->1	
i.En 	ö->1	
i.Ett	 ->1	
i.Eur	o->1	
i.Fol	k->1	
i.For	s->1	
i.Fru	 ->1	
i.För	 ->1	
i.Hai	d->1	
i.Her	r->1	
i.Hur	 ->1	
i.Här	 ->1	
i.I k	o->1	
i.Jag	 ->3	
i.Kan	s->1	
i.Kul	t->1	
i.Lik	r->1	
i.Man	 ->2	
i.Min	 ->1	
i.När	 ->1	
i.Sed	a->1	
i.Som	 ->1	
i.Så 	ä->1	
i.Utv	i->1	
i.Vi 	a->1	f->1	s->1	
i.Vid	 ->1	
i.Vil	l->1	
i.Vår	 ->1	
i: fr	å->1	
i; ma	n->1	
i? Oc	h->1	
i?.He	r->1	
ia - 	r->1	s->1	
ia Br	y->1	
ia Eu	r->1	
ia Pa	l->1	
ia Ro	t->1	
ia al	l->2	
ia at	t->2	
ia bi	l->1	
ia da	 ->1	
ia de	 ->1	t->1	
ia en	s->1	
ia fr	å->1	
ia fu	n->1	
ia ha	r->1	
ia i 	E->1	
ia in	k->1	
ia ko	m->1	
ia ma	r->1	
ia oc	h->2	
ia om	 ->1	b->1	
ia rö	r->10	
ia sa	m->1	
ia sk	u->1	
ia so	m->2	
ia st	r->2	
ia ti	l->2	
ia ty	p->1	
ia un	i->1	
ia va	l->3	
ia vä	r->1	
ia åt	e->1	
ia, d	e->1	
ia, e	n->1	
ia, o	b->1	
ia, r	e->1	
ia-Ro	m->1	
ia.De	t->1	
ia.Än	t->1	
iagen	t->1	
iaktt	a->8	
ial -	 ->1	
ial b	e->1	
ial d	u->2	
ial f	r->2	
ial i	 ->1	
ial k	a->1	
ial m	e->1	
ial n	o->1	
ial o	c->6	
ial r	ä->2	
ial s	a->7	e->1	o->3	t->2	y->1	
ial t	i->1	r->3	
ial u	t->8	
ial, 	a->1	d->1	t->1	
ial- 	o->1	
ial.D	e->2	
ial.F	ö->2	
ial.J	a->1	
ial.S	j->1	
iala 	E->1	a->1	b->2	d->5	e->5	f->5	i->2	k->2	m->4	o->19	p->8	r->2	s->14	t->1	u->5	v->1	ä->1	
ialbe	s->2	
ialde	m->15	
ialdo	m->1	
ialen	,->1	
ialet	 ->1	,->2	
ialfo	n->15	r->2	
ialfr	å->5	
ialfö	r->6	
ialin	r->1	
ialis	e->5	m->2	t->34	
ialog	 ->15	,->1	.->7	e->8	
ialpo	l->4	
ialpr	o->1	
ialt 	a->4	h->5	m->1	p->2	r->3	s->1	
ialt,	 ->1	
ialt.	D->1	
ialut	b->1	
ian 1	9->1	
iane 	o->2	
iane,	 ->1	
iano 	u->1	
ians 	m->2	s->1	
ianse	n->3	r->1	
iansp	r->1	
ianvä	n->6	
iarit	e->21	
ias f	r->3	
ias o	c->1	
iasm 	f->1	p->1	s->1	
iat f	ö->1	
iat h	o->1	
iat.M	e->1	
iatis	k->4	
iativ	 ->42	,->7	.->7	a->1	b->1	e->16	f->1	r->5	
iatäc	k->1	
ibakt	e->1	
ibane	s->1	
ibano	n->5	
ibbig	a->1	
ibedr	ä->1	
ibehå	l->11	
ibekä	m->4	
ibel 	l->1	o->1	u->1	
ibel,	 ->1	
ibel.	V->1	
ibelt	 ->6	
ibera	l->31	
iberi	s->1	
ibesp	a->3	
ibest	ä->2	
ibet 	F->1	d->1	h->1	m->1	o->3	s->2	t->1	u->2	
ibet"	 ->1	,->1	
ibet,	 ->3	
ibet-	f->1	
ibet.	E->1	V->1	
ibet?	J->1	
ibeta	n->10	
ibi n	ä->1	
ibili	t->11	
ibla 	a->1	f->1	o->1	
ibla.	D->1	
iblan	d->25	
iblar	e->2	
iblio	t->2	
ibuti	o->1	
ibyen	s->1	
ic - 	o->1	
ic Br	a->1	
ic i 	d->1	
ical 	c->1	
icant	e->1	
icap 	ä->1	
ice d	e->4	
ice f	ö->1	
ice n	a->1	
ice o	r->11	
ice t	a->2	
ice.A	l->1	
ice.J	a->1	
ice.O	f->1	
ice.S	t->1	
iceko	r->1	
icekv	a->1	
icen,	 ->1	
icens	i->1	
icent	r->1	
icera	 ->4	d->25	n->3	r->5	s->1	t->9	
iceri	n->10	
ichar	d->1	
icher	 ->1	
ichie	l->1	
icht 	m->1	o->1	
icht.	D->1	
ichte	r->2	
ichtf	ö->3	
ichyr	e->1	
iciel	l->7	
icien	,->2	t->1	
icine	r->1	
icio 	S->1	
icit.	F->1	
icite	t->2	
ick -	 ->1	
ick K	i->1	
ick a	t->1	
ick b	a->2	e->1	
ick d	e->3	
ick e	f->1	m->1	n->2	t->1	
ick f	r->1	ö->1	
ick h	ö->2	
ick i	 ->3	n->3	
ick j	a->3	u->2	
ick k	ä->1	
ick m	e->1	i->1	y->1	ö->1	
ick n	e->1	å->2	
ick o	c->2	s->2	
ick s	e->1	n->1	t->1	
ick t	i->3	
ick u	p->1	
ick v	a->1	i->3	
ick, 	1->1	f->1	n->1	
ick.A	v->1	
ick.D	e->1	
ick.H	e->1	
ick.K	o->1	
ick.Ä	v->1	
icka 	e->1	n->1	p->1	u->2	v->1	
icka,	 ->1	
ickad	e->2	
ickar	 ->3	
ickas	 ->1	
ickat	 ->2	
ickba	r->5	
icke 	b->1	e->2	f->2	i->1	k->2	l->2	o->1	s->1	t->1	v->1	ö->1	
icke-	a->2	d->3	f->1	m->1	s->12	
icken	 ->1	
icker	 ->2	
icket	 ->6	,->2	.->1	;->1	m->1	
ickfr	i->1	
ickli	g->1	
ickni	n->1	
ickor	n->1	s->1	
ickpr	o->3	
icks.	P->1	
icksi	l->3	
icksv	a->1	
icy, 	s->1	
icyav	t->1	
icyde	l->1	
icyfö	r->1	
id 12	 ->1	
id 70	0->1	
id By	r->3	
id EG	-->3	
id EU	-->1	
id Eu	r->4	
id Ge	n->1	
id Ha	i->1	
id Ky	o->1	
id La	n->1	
id Me	d->1	
id Pa	d->1	
id a)	 ->1	
id al	l->3	
id an	d->3	l->1	t->3	v->1	
id ar	t->1	
id at	t->27	
id av	 ->3	
id ba	r->1	
id be	d->1	h->6	s->1	t->1	
id bl	i->2	
id br	a->1	
id bä	t->1	
id bö	r->5	
id ca	.->1	
id da	g->1	
id de	 ->5	n->17	r->1	s->5	t->13	
id do	m->2	
id dr	o->1	
id dä	r->1	
id då	 ->3	
id ef	f->1	t->1	
id el	l->1	
id en	 ->9	d->1	
id et	t->12	
id ev	e->1	
id fa	l->1	s->1	
id fi	n->2	
id fl	e->5	y->1	
id fr	a->3	å->2	
id fu	n->1	
id fy	s->1	
id få	r->1	t->1	
id fö	r->20	
id gj	o->2	
id go	t->1	
id gr	a->1	ä->1	
id gö	r->1	
id ha	 ->1	l->1	n->2	r->11	
id he	l->1	
id hi	t->1	
id hj	ä->1	
id hä	v->1	
id hö	j->1	r->2	
id i 	E->1	d->4	e->1	v->1	
id in	g->1	s->1	t->8	
id ja	g->1	
id jo	r->1	
id jä	m->1	
id ka	n->5	
id kl	i->1	
id ko	m->6	
id kr	i->1	ä->1	
id ku	l->1	s->1	
id kä	r->1	
id la	g->1	
id li	v->1	
id lu	n->1	
id lä	g->1	t->1	
id ma	n->1	
id me	d->8	n->1	
id mi	l->1	n->2	
id mo	t->2	
id my	c->1	
id mä	n->1	
id må	s->2	
id mö	t->3	
id na	t->3	
id no	t->1	
id nu	v->1	
id ny	p->1	
id nä	m->1	s->1	
id nå	g->2	
id oc	h->6	k->1	
id oe	r->1	
id of	f->1	
id om	 ->1	r->5	s->1	
id op	t->1	
id or	d->1	
id pa	r->1	s->1	
id pl	a->1	e->1	
id pr	i->2	o->1	
id pu	n->2	
id på	 ->4	
id re	g->4	
id rä	t->2	
id rå	d->1	
id sa	m->3	
id se	 ->1	
id si	d->8	
id sj	ä->1	ö->1	
id sk	a->4	u->1	
id sl	u->1	ö->1	
id so	m->4	
id st	a->1	o->1	r->1	ä->1	å->1	ö->1	
id sy	f->1	
id sä	g->1	k->1	
id så	 ->2	
id ta	 ->1	l->2	
id te	m->1	
id ti	d->1	l->7	
id to	p->2	
id tr	a->3	e->1	
id tv	å->2	
id un	d->2	
id up	p->3	
id ut	a->4	b->1	f->1	g->1	n->1	s->1	v->2	
id va	c->1	l->2	r->3	
id vi	 ->1	k->2	l->2	s->2	
id vå	r->1	
id yr	k->1	
id än	 ->1	n->1	
id är	 ->8	
id äv	e->1	
id år	e->1	t->1	
id åt	 ->1	e->2	
id öv	e->2	
id, a	t->2	
id, d	e->1	
id, e	n->1	
id, f	ö->1	
id, h	a->1	e->1	
id, i	 ->1	n->1	
id, m	e->1	
id, o	c->3	m->1	
id, p	l->1	
id, v	a->2	i->1	
id, ä	r->1	
id.. 	(->1	
id.De	 ->2	n->1	t->2	
id.En	 ->1	
id.Fö	r->1	
id.Ha	n->1	
id.Ja	g->1	
id.Ko	m->1	
id.Ma	n->1	
id.Nä	r->1	
id.Om	 ->1	
id.So	m->1	
id.Ta	c->1	
id.Ti	l->1	
id.Vi	 ->1	
id: d	e->1	
ida E	U->1	
ida G	o->1	
ida a	t->2	
ida b	e->2	i->2	
ida d	e->10	i->1	
ida e	k->1	u->1	
ida f	i->1	o->1	r->1	ö->2	
ida g	ö->1	
ida h	ö->1	
ida i	 ->3	n->4	
ida k	o->4	r->1	
ida m	e->1	o->2	
ida n	i->1	å->1	
ida o	c->2	
ida p	r->1	
ida r	e->1	
ida s	c->1	e->1	i->1	k->2	o->1	
ida t	i->2	r->1	u->1	
ida u	n->1	
ida v	a->2	i->1	
ida å	t->1	
ida, 	b->1	f->2	i->1	o->2	s->2	v->1	
ida.D	e->1	
ida.F	r->1	
ida.H	e->1	
ida.I	b->1	
ida.J	a->1	
ida.O	c->1	
ida.V	i->1	
ida.Ä	v->1	
ida?I	n->1	
idag,	 ->1	
idaki	s->2	
idan 	a->7	b->3	d->1	e->1	f->5	h->4	k->3	l->1	m->1	o->6	r->1	s->1	t->2	v->3	ä->3	ö->1	
idan,	 ->2	
idan.	J->1	
idand	e->15	
idare	 ->29	.->7	?->1	b->3	u->4	
idari	s->2	t->29	
idas 	ö->1	
idat 	s->1	
idate	r->1	
idatl	a->1	i->1	ä->10	
idd b	ö->1	
idd h	ä->1	
idd m	o->1	
idd o	c->1	
idd ä	n->1	
idd.J	a->1	
iddag	 ->4	,->2	.->1	e->2	s->4	
iddel	h->1	
idden	 ->1	
ide W	e->1	
ideal	,->1	a->1	e->2	i->1	
ideel	l->2	
idemo	k->1	
iden 	2->1	a->5	b->3	f->11	g->4	h->5	i->3	k->8	l->1	m->2	n->1	o->5	p->3	r->1	s->9	t->2	v->5	ä->4	ö->3	
iden,	 ->7	
iden.	A->1	D->7	E->5	H->1	I->1	J->1	K->2	M->3	N->3	P->1	S->2	U->1	V->3	
iden:	 ->1	
iden?	D->1	V->1	
idens	 ->3	
ident	 ->5	,->1	e->4	i->20	
ideol	o->5	
ider 	a->5	d->3	e->2	f->2	g->1	h->1	i->5	k->3	l->1	m->4	o->5	p->1	r->1	s->7	t->3	u->3	ä->1	
ider,	 ->5	
ider.	.->1	C->1	D->2	S->1	
idera	 ->5	d->1	s->2	
ideri	n->13	
iders	 ->19	
ides 	b->1	m->1	
idga 	E->2	d->4	f->1	g->1	k->1	m->2	o->1	u->2	
idga?	D->1	
idgad	 ->4	e->1	
idgar	 ->3	
idgas	 ->5	,->2	.->6	
idgat	 ->2	
idgni	n->71	
idhål	l->4	
idhöl	l->1	
idiar	i->21	
idig 	e->1	f->1	h->1	i->1	r->2	t->1	
idiga	 ->3	r->81	
idigh	e->1	
idigt	 ->77	.->1	
idisk	 ->7	a->14	t->10	
idit 	a->1	f->2	
idits	 ->1	
idiär	,->1	
idkar	e->1	
idlag	 ->1	
idlan	d->1	
idlig	a->1	e->1	t->3	
idmak	t->1	
idnap	p->1	
idnin	g->22	
idoef	f->1	
idor 	f->1	h->1	o->1	
idor.	D->1	
idore	r->2	
idorn	a->2	
idosk	o->2	
idpun	k->10	
idra 	m->3	s->1	t->31	
idra,	 ->1	
idrag	 ->28	.->2	:->1	e->3	i->9	s->9	
idrar	 ->20	
idrog	 ->3	
idrot	t->4	
ids i	 ->1	
ids m	e->1	
ids p	å->1	
ids t	i->1	
ids u	t->1	
ids ä	n->1	
ids, 	o->1	
ids-s	i->1	
idsar	b->4	
idsbe	d->1	s->1	
idsdi	r->3	
idsdu	g->1	
idsfr	i->10	
idsfö	r->1	
idsgr	ä->1	
idsin	r->1	s->1	
idsmä	s->2	
idsor	i->1	
idspa	t->2	
idspe	n->6	r->4	
idspl	a->5	
idsra	m->5	
idsry	m->2	
idssk	ä->1	
idssy	s->1	
idstr	ä->1	
idsål	d->2	
idsåt	g->1	
idsöd	a->1	
idta 	d->2	e->6	f->9	g->1	k->1	l->1	m->3	n->1	o->1	p->2	s->1	å->5	
idtab	e->6	
idtag	i->5	n->1	
idtal	a->1	
idtar	 ->8	
idtas	 ->10	,->2	.->2	
idtog	 ->1	s->1	
idual	i->1	
iduel	l->7	
iduer	,->1	
iduts	l->1	
idé -	 ->1	
idé a	t->2	
idé j	a->1	
idé k	o->1	
idé o	m->1	
idé s	o->3	
idé ä	r->1	
idé, 	m->1	
idéer	 ->6	,->1	n->1	
idén 	a->6	b->3	m->1	o->2	v->1	
idén,	 ->1	
ie Cu	r->1	
ie Re	p->1	
ie av	 ->1	
ie oc	h->1	
ie, h	ö->1	
ie- o	c->1	
ie-st	i->1	
ieben	g->1	
iebes	ö->1	
iebör	s->1	
ieck 	h->1	
ied (	a->1	
ied.K	o->1	
iedep	a->2	
ieffe	k->6	
iefin	g->1	
iefus	i->1	
iekti	v->1	
iel v	a->1	
ielan	d->4	
ielft	e->1	
iell 	b->1	d->1	f->1	g->1	i->1	k->1	n->2	o->2	p->1	r->1	t->1	å->1	ö->1	
iell,	 ->1	
iella	 ->60	,->1	
iellt	 ->41	,->1	
ielse	 ->2	n->5	
ielso	n->5	
iemin	i->3	
ien 9	0->1	
ien a	t->3	
ien b	e->1	
ien d	ä->1	
ien e	f->1	l->2	
ien f	i->1	ö->2	
ien h	a->8	o->1	
ien i	 ->2	n->1	
ien j	u->1	
ien m	å->1	
ien n	ä->1	
ien o	c->21	
ien s	k->2	o->6	å->1	
ien t	i->3	
ien ä	n->1	r->5	
ien, 	B->1	I->1	K->1	P->1	S->1	T->1	b->1	d->1	e->2	f->1	j->1	m->1	o->2	s->1	t->2	u->1	v->2	Î->1	ä->1	
ien.D	e->1	ä->1	
ien.E	t->1	
ien.F	ö->1	
ien.H	e->1	
ien.I	 ->1	
ien.M	ä->1	
ien.O	z->1	
ien.P	l->1	
ien.S	a->1	t->1	
ien.U	t->1	
ien.V	i->1	
ien?E	f->1	
ien?V	i->1	
iende	,->1	
ienfr	å->1	
ienne	 ->1	
iens 	g->2	i->1	k->1	p->1	r->1	s->1	t->2	u->1	
iense	r->2	
iensk	 ->1	a->12	e->2	t->2	
ient 	i->1	
iente	n->1	r->9	
ienti	f->1	l->1	
ientl	i->33	
iepro	g->1	
ier -	 ->6	
ier D	u->1	
ier a	t->2	v->1	
ier e	l->2	
ier f	i->1	r->1	ö->11	
ier g	e->1	
ier h	a->3	
ier i	 ->1	
ier k	a->1	o->3	
ier m	e->3	å->1	
ier o	c->17	m->4	
ier p	å->2	
ier r	e->1	ö->2	
ier s	a->1	k->2	o->14	
ier t	o->1	
ier u	p->1	t->1	
ier ä	n->1	
ier ö	k->1	
ier, 	a->2	d->1	f->1	h->1	m->3	o->3	s->3	t->1	u->1	
ier..	H->1	
ier.A	l->1	
ier.D	e->4	
ier.K	o->1	v->1	
ier.L	å->1	
ier.M	e->2	
iera 	E->1	b->1	d->1	e->2	f->1	i->1	o->3	s->2	v->4	
ierad	 ->5	e->11	
ierar	 ->3	k->4	
ieras	 ->8	,->2	.->1	
ierat	 ->8	,->1	.->2	s->1	
ierba	r->2	
ierdo	 ->1	
ierin	g->43	
ierna	 ->36	,->2	.->4	s->2	
iers 	u->2	
ies a	n->1	
ies r	ä->1	
ies v	a->1	
ieski	f->2	
iesmi	t->1	
iestr	a->1	
iet (	F->1	S->1	Ö->1	
iet D	e->1	
iet I	 ->1	
iet a	t->2	
iet d	å->1	
iet e	n->1	t->1	
iet f	ö->1	
iet h	a->6	e->1	
iet i	 ->1	n->2	
iet m	å->1	
iet n	u->1	ä->1	
iet o	c->7	
iet p	l->1	
iet r	e->1	
iet s	o->3	ö->1	
iet t	i->1	
iet v	i->1	
iet ä	r->3	
iet".	E->1	
iet) 	p->1	
iet),	 ->2	
iet).	D->1	
iet, 	H->1	b->3	h->1	s->4	
iet.A	v->1	
iet.D	e->2	
iet.H	e->1	
iet.M	e->1	
iet.O	m->1	
iet.V	a->1	i->2	
ietni	s->3	
iets 	a->1	f->2	g->12	k->2	m->1	p->2	s->1	v->1	
iety 	ä->1	
ieuro	p->1	
ieäga	r->2	
ifall	 ->2	,->1	a->1	i->1	
ifart	e->2	
ifasc	i->3	
ifera	 ->3	.->1	
iferi	n->1	
ifert	.->1	
ifest	a->1	
iffer	e->5	
iffra	 ->4	,->3	
iffro	r->15	
ifice	r->38	
ifici	e->2	
ifier	a->22	b->2	i->3	
ifik 	o->1	s->1	å->1	
ifika	 ->17	t->5	
ifikt	 ->7	
ifin-	r->1	
ifina	n->1	
ifiqu	e->1	
ifolk	l->1	
ifond	e->2	
iform	e->1	
ifråg	a->22	o->4	
ifrån	 ->31	,->2	.->2	
ift a	t->2	v->1	
ift d	e->1	
ift e	r->1	
ift f	r->1	ö->2	
ift i	 ->2	
ift k	o->1	
ift m	e->1	
ift o	c->1	m->1	
ift p	å->1	
ift r	e->1	
ift s	k->1	o->4	
ift t	i->1	
ift v	i->1	
ift ä	r->3	
ift!H	e->1	
ift, 	i->1	o->1	
ift. 	D->1	
ift.A	t->1	
ift.D	e->1	
ift.E	f->1	
ift.J	a->1	
ift.O	m->1	
ift.V	i->1	
ift: 	d->1	
ifta 	f->1	i->1	l->1	p->1	
iftan	d->5	
iftar	 ->4	n->2	
iftat	 ->1	
ifte 	u->1	
ifte,	 ->1	
ifte.	V->1	
iften	 ->7	.->1	
ifter	 ->32	,->6	.->5	:->1	n->20	
iftet	 ->2	.->1	
iftig	a->3	
iftli	g->8	
iftni	n->113	
ifts-	 ->1	
iftsf	ö->2	
iftsl	ä->2	
iftsm	å->1	
iftsp	o->1	r->1	
iftss	e->1	
iftst	a->1	
iftsä	k->1	
ifull	a->1	
iförb	r->1	
iförr	å->1	
iförs	ö->2	
ig - 	a->1	
ig -,	 ->1	
ig Eu	r->1	
ig OL	A->1	
ig ac	c->1	
ig al	d->1	l->4	
ig an	 ->2	d->1	g->1	l->2	s->2	v->2	
ig ar	a->1	b->2	t->1	
ig as	s->2	
ig at	t->63	
ig av	 ->12	e->1	s->2	
ig ba	k->4	r->6	
ig be	f->1	g->1	h->2	r->2	s->6	t->1	v->1	
ig bi	l->1	
ig bl	a->1	i->1	
ig bo	r->1	
ig br	a->2	o->1	
ig by	r->2	
ig bä	r->2	
ig bö	r->1	
ig da	g->1	
ig de	b->8	l->10	m->2	n->6	s->2	t->7	
ig di	a->2	r->1	s->1	
ig dj	u->1	
ig do	c->2	
ig dä	r->3	
ig dö	d->1	r->1	
ig ef	f->2	t->2	
ig ek	o->1	
ig el	l->5	
ig em	e->1	o->3	
ig en	 ->8	d->1	h->1	s->1	
ig er	 ->1	
ig et	t->6	
ig eu	r->1	
ig ex	a->1	p->1	
ig fa	k->1	
ig fi	n->1	
ig fo	r->1	
ig fr	a->3	e->4	i->1	å->21	
ig fu	l->1	n->3	
ig få	r->2	
ig fö	r->86	
ig ga	r->1	
ig ge	 ->1	n->1	
ig gi	v->2	
ig gl	o->1	
ig gr	a->2	u->8	
ig gä	l->1	r->1	
ig gö	r->2	
ig ha	 ->1	n->4	r->5	
ig he	l->2	m->1	
ig hi	e->1	s->1	
ig hj	ä->3	
ig hu	r->2	v->1	
ig hä	n->5	
ig i 	D->1	E->3	K->1	S->1	Y->1	b->1	d->9	e->8	f->1	h->1	k->3	m->1	o->1	r->1	s->3	t->1	u->2	v->1	
ig i.	S->1	
ig ih	o->1	
ig in	 ->8	f->10	g->1	o->2	r->2	s->3	t->10	
ig iv	ä->1	
ig jo	n->1	
ig ju	 ->1	r->1	s->1	
ig jä	m->1	
ig ka	n->2	p->1	r->2	t->2	
ig kl	a->1	
ig kn	a->1	
ig ko	m->7	n->9	r->1	s->3	
ig kr	i->1	
ig ku	l->2	n->1	
ig kv	a->1	
ig kä	r->1	
ig la	g->3	r->1	
ig le	d->2	g->1	
ig li	t->1	
ig lä	n->1	s->1	x->1	
ig lö	s->5	
ig ma	j->1	k->3	n->4	r->1	x->1	
ig me	d->14	l->1	n->3	r->7	s->1	
ig mi	l->2	n->2	
ig mo	t->8	
ig my	c->9	n->1	
ig mä	r->1	
ig må	n->3	s->1	
ig mö	j->2	
ig na	i->1	t->1	
ig ne	d->3	
ig ni	v->3	
ig no	g->2	
ig nu	 ->1	
ig ny	n->1	
ig nä	r->6	s->1	
ig nå	g->1	
ig nö	d->1	
ig ob	e->2	
ig oc	h->46	k->7	
ig oe	r->1	
ig of	f->2	
ig om	 ->36	e->1	f->1	p->1	s->1	
ig on	d->1	ö->1	
ig or	i->1	o->1	
ig pa	r->1	
ig pe	r->4	
ig po	l->6	s->1	
ig pr	a->1	e->1	o->2	
ig pu	n->7	
ig på	 ->31	,->1	m->2	p->1	v->2	
ig ra	m->2	p->1	
ig re	a->2	d->1	f->4	g->3	l->1	s->3	v->1	
ig ri	k->1	s->2	
ig ro	l->8	
ig ru	m->1	
ig ry	k->1	
ig rä	t->2	
ig rå	d->2	
ig sa	g->1	k->1	m->6	
ig se	g->1	k->3	m->1	r->1	
ig si	g->3	m->1	t->4	
ig sj	ä->11	
ig sk	a->2	i->1	u->1	y->1	
ig sl	u->2	
ig so	l->2	m->9	
ig st	a->3	r->4	ä->1	ö->2	
ig su	b->1	
ig sv	a->1	
ig sy	n->1	s->1	
ig sä	g->2	k->2	n->1	r->3	t->1	
ig så	 ->1	l->1	
ig t.	e->1	
ig ta	 ->1	c->1	
ig te	k->2	
ig ti	d->8	l->42	
ig to	l->1	
ig tr	a->1	
ig tv	e->1	i->1	
ig ty	d->1	
ig un	d->5	
ig up	p->7	
ig ut	 ->3	a->2	b->4	e->2	f->3	g->2	m->2	s->6	v->2	ö->1	
ig va	d->3	k->1	r->14	
ig ve	t->1	
ig vi	 ->2	d->1	l->3	
ig vä	g->1	l->2	r->1	
ig yr	k->1	
ig yt	t->1	
ig än	d->3	
ig är	 ->9	
ig äv	e->2	
ig å 	P->1	
ig åk	l->1	
ig ås	i->3	
ig åt	 ->16	,->1	g->2	s->1	
ig ök	n->1	
ig öv	e->8	n->1	
ig!".	D->1	
ig!Ha	n->1	
ig".E	u->1	
ig, a	n->1	t->2	v->1	
ig, b	l->1	å->1	
ig, d	e->3	
ig, e	f->2	n->2	
ig, f	ö->2	
ig, g	r->1	ö->1	
ig, h	a->1	e->4	
ig, i	r->1	
ig, l	å->1	
ig, m	e->2	i->1	å->1	
ig, n	ä->4	
ig, o	c->3	m->1	t->1	
ig, p	å->1	
ig, s	k->1	n->1	o->1	t->1	ä->2	å->2	
ig, u	t->1	
ig, v	i->3	
ig. F	ö->1	
ig. S	å->1	
ig.Av	 ->1	
ig.Br	i->1	
ig.De	 ->2	n->3	t->5	
ig.Em	e->1	
ig.En	 ->1	
ig.Er	i->1	
ig.Eu	r->1	
ig.Ge	n->1	
ig.Gr	u->1	
ig.He	r->2	
ig.I 	n->1	
ig.Ja	g->13	
ig.Ko	n->1	
ig.Ma	n->1	r->1	
ig.Me	d->1	n->1	
ig.Na	t->1	
ig.Oc	h->3	
ig.Pr	o->1	
ig.Sa	m->1	
ig.Ta	c->1	
ig.Un	d->1	
ig.Va	r->1	
ig.Vi	 ->4	
ig.Är	 ->1	
ig: d	e->1	i->1	
ig: h	a->1	
ig; d	e->1	
ig?De	t->1	
ig?Hu	r->1	
ig?Jo	,->1	
ig?Va	d->1	
iga "	A->1	
iga -	 ->5	
iga 3	7->1	
iga E	U->1	u->3	
iga H	a->1	
iga a	d->2	g->2	k->1	l->1	n->3	p->2	r->7	t->12	v->4	
iga b	a->1	e->32	i->10	l->1	r->6	u->4	å->1	
iga c	h->1	
iga d	e->17	i->3	o->2	å->1	
iga e	f->3	g->1	k->1	l->4	n->5	r->1	t->2	u->2	x->1	
iga f	a->5	e->1	i->4	o->5	r->56	å->1	ö->66	
iga g	a->3	e->4	i->3	n->1	r->11	
iga h	a->6	i->1	o->1	y->1	ä->5	
iga i	 ->13	.->1	a->1	d->1	f->1	m->1	n->24	r->1	
iga k	a->3	l->1	o->30	r->5	v->1	ä->1	
iga l	a->2	e->1	i->9	o->1	ä->8	ö->4	
iga m	a->3	e->22	i->6	o->5	y->1	ä->2	å->7	ö->1	
iga n	a->2	e->1	i->1	o->1	y->2	ä->2	
iga o	c->57	f->1	m->11	r->15	s->1	
iga p	a->3	e->2	l->2	o->6	r->17	u->2	å->5	
iga r	a->6	e->25	i->3	o->1	ä->38	å->5	
iga s	a->7	c->1	e->7	i->3	k->5	l->1	o->5	p->3	t->64	u->1	v->4	y->5	ä->3	å->2	
iga t	a->5	e->5	i->6	j->3	r->3	u->2	
iga u	n->1	p->7	t->10	
iga v	a->3	e->5	i->3	r->2	ä->8	å->1	
iga y	t->1	
iga ä	m->12	n->6	r->3	v->1	
iga å	k->1	s->1	t->11	
iga ö	a->1	n->1	p->1	v->6	
iga, 	a->2	e->4	f->2	i->2	k->2	m->2	n->1	o->8	p->4	r->1	u->1	v->4	ä->1	
iga. 	M->1	
iga.(	T->1	
iga.A	l->1	v->2	
iga.D	e->3	
iga.E	n->1	
iga.F	ö->3	
iga.H	e->2	
iga.I	 ->3	n->1	
iga.J	a->1	
iga.M	a->1	e->1	
iga.N	i->2	
iga.O	m->1	
iga.P	å->2	
iga.S	å->1	
iga.V	i->4	
iga/h	a->1	
iga; 	v->1	
iga?F	ö->1	
igad,	 ->1	
igad.	D->1	K->1	
igade	 ->7	s->1	
igand	e->11	
igant	i->5	
igar 	a->1	e->2	k->1	
igare	 ->152	,->7	.->6	l->1	
igas 	a->1	d->1	f->1	ä->1	
igas,	 ->2	
igast	 ->1	,->1	e->50	
igat 	a->4	f->1	s->3	
igat,	 ->2	
igat.	D->1	
igato	r->14	
igats	 ->2	
igdom	 ->3	,->2	.->1	/->1	e->4	s->1	
ige i	 ->1	
ige o	c->3	
ige p	i->1	
ige s	o->1	
ige. 	D->1	
ige.J	a->1	
igen 	-->1	1->1	E->1	F->1	J->1	K->1	W->1	a->44	b->33	d->12	e->26	f->40	g->18	h->39	i->36	k->35	l->7	m->26	n->6	o->12	p->14	r->12	s->32	t->23	u->8	v->28	ä->19	å->2	ö->3	
igen"	,->1	
igen,	 ->27	
igen.	C->1	D->3	F->1	H->1	I->1	J->1	M->1	R->1	S->1	V->1	
igen:	 ->2	
igena	r->3	
igenk	ä->1	
igeno	m->37	
igens	e->1	k->1	
igent	 ->3	a->1	
iger 	5->1	i->1	
iger.	H->1	
igera	r->1	
igern	 ->1	
iges 	a->1	
iget 	-->1	1->1	o->1	p->1	s->1	
iget.	E->1	J->1	P->1	
igets	 ->4	
igga 	b->1	h->1	i->2	k->1	p->1	s->1	t->4	u->1	v->1	
iggan	d->10	
igger	 ->81	,->3	.->2	;->1	
iggjo	r->13	
iggör	 ->5	a->12	s->4	
igh l	e->1	
ighet	 ->216	!->1	"->1	,->33	.->38	?->1	e->459	s->81	
ight 	k->1	t->1	
ights	.->1	
ighål	l->2	
igier	a->1	
igina	l->1	
igine	l->1	
igit 	m->1	
igit.	F->1	
igiös	 ->1	a->2	t->1	
igjor	d->1	
iglan	d->1	
iglig	 ->3	t->1	
igmat	i->1	
igna 	o->1	
ignal	 ->9	e->5	
ignel	s->1	
igner	a->1	
ignor	e->4	
igorö	s->4	
igott	e->1	
igou 	o->1	
igra 	o->1	s->1	
igran	t->2	
igrat	i->8	
igrer	a->1	
igsek	t->1	
igshe	r->1	
igssk	a->1	
igstä	l->1	
igt -	 ->6	
igt :	 ->1	
igt D	u->1	
igt E	u->2	
igt G	r->1	
igt I	n->1	
igt K	y->1	
igt R	a->1	
igt S	c->1	
igt T	h->1	
igt a	d->1	l->1	n->5	r->14	s->1	t->185	v->19	
igt b	e->19	i->4	l->1	r->4	ä->1	
igt d	a->1	e->24	i->3	j->1	r->1	
igt e	f->10	g->1	l->4	n->7	r->3	t->3	u->1	x->5	
igt f	a->2	e->3	i->2	l->1	o->2	r->7	u->1	å->1	ö->75	
igt g	e->3	o->40	r->3	ä->1	
igt h	a->14	e->1	i->1	o->5	u->1	ä->3	å->1	ö->5	
igt i	 ->20	c->1	n->20	
igt j	a->1	u->1	
igt k	a->4	l->1	n->1	o->16	r->4	ä->2	
igt l	i->5	ä->7	å->3	
igt m	a->1	e->30	i->37	o->3	y->5	å->11	ö->2	
igt n	a->1	o->8	ä->5	
igt o	a->4	b->2	c->58	f->3	m->4	r->6	s->1	t->2	
igt p	a->5	e->1	l->1	o->4	r->16	å->8	
igt r	e->11	y->1	ä->1	
igt s	a->8	e->4	i->2	j->1	k->15	l->2	o->23	p->2	t->36	u->1	v->4	y->6	ä->32	å->1	
igt t	a->11	e->2	i->14	o->1	y->2	ä->1	
igt u	n->5	p->8	r->1	t->8	
igt v	a->6	e->1	i->29	ä->3	å->6	
igt y	t->2	
igt ä	n->2	r->13	v->1	
igt å	t->3	
igt ö	g->1	n->1	v->3	
igt!L	e->1	
igt!M	e->1	
igt, 	a->1	b->2	d->4	e->5	f->6	h->1	i->4	j->3	k->5	l->2	m->5	n->2	o->10	r->1	s->8	u->2	ä->1	
igt.A	r->1	
igt.D	e->10	i->1	
igt.E	f->1	n->1	t->1	
igt.F	r->2	ö->6	
igt.G	e->2	
igt.H	e->4	u->1	
igt.I	 ->1	
igt.J	a->11	
igt.L	å->2	
igt.M	a->1	e->4	i->3	o->1	
igt.N	a->1	ä->1	
igt.O	f->1	m->2	
igt.P	å->1	
igt.S	o->1	t->2	
igt.U	n->1	
igt.V	a->4	i->9	
igt.Ö	k->1	
igt: 	d->1	
igt; 	d->1	
igt?A	v->1	
igtvi	s->108	
igvat	t->1	
igå d	e->1	
igåen	d->4	
igång	 ->4	.->1	k->1	s->1	
igås 	i->1	
igör 	h->1	
igöra	 ->2	n->1	s->1	
igörs	 ->1	
ihan;	 ->1	
ihand	e->2	
ihet 	1->1	a->6	b->1	e->2	f->14	i->3	n->1	o->10	s->2	u->1	ä->2	å->1	
ihet,	 ->38	
ihet.	D->1	F->1	I->1	J->1	V->1	
ihet:	 ->1	
ihet;	 ->1	
ihete	n->20	r->5	
ihets	k->1	r->1	
ihjäl	 ->1	
ihop 	a->1	d->1	f->1	p->1	s->1	t->1	u->1	ä->1	
ihop,	 ->1	
ihop.	D->1	I->1	J->1	
ihärd	i->1	
ihåg 	I->1	a->8	d->3	r->1	s->1	ä->1	
ihåg.	E->1	
iikan	e->3	
iimpo	r->1	
iinne	h->1	
iintr	e->1	
iis-J	ø->2	
ij-va	n->1	
ijs o	c->1	
ijs.(	E->1	
ik - 	d->2	
ik De	t->1	
ik Jö	r->1	
ik an	t->1	
ik av	 ->4	
ik eg	e->1	
ik el	l->2	
ik en	 ->1	
ik et	a->1	
ik fi	n->1	
ik fr	ä->1	
ik få	r->1	
ik fö	r->16	
ik ha	r->3	
ik hu	v->1	
ik hö	r->1	
ik i 	E->1	a->1	f->1	n->1	o->1	s->2	v->2	
ik in	d->1	t->1	
ik ka	n->2	
ik ku	n->1	
ik me	d->4	l->1	
ik mi	g->1	
ik mo	d->1	t->2	
ik må	s->3	
ik mö	j->1	
ik nä	r->3	
ik oc	h->28	
ik om	 ->2	
ik or	i->1	
ik po	l->2	
ik på	 ->3	
ik re	k->1	
ik rö	r->1	
ik sa	m->1	
ik sk	ö->1	
ik so	m->31	
ik st	r->1	
ik så	 ->1	
ik ti	l->1	
ik un	d->1	
ik up	p->1	
ik ut	g->1	
ik va	r->1	
ik vi	 ->1	l->1	
ik är	 ->5	
ik åt	e->1	
ik öv	e->1	
ik!Om	 ->1	
ik" o	c->1	
ik, d	e->3	v->2	å->1	
ik, e	n->2	
ik, f	r->1	ö->1	
ik, h	a->1	
ik, i	n->2	
ik, m	o->1	
ik, n	e->1	ä->1	å->1	
ik, o	c->1	
ik, s	a->2	o->1	
ik, t	r->10	
ik, u	t->1	
ik, v	a->2	i->1	
ik- o	c->2	
ik..(	F->1	
ik.By	g->1	
ik.De	 ->1	n->1	t->7	
ik.Dä	r->1	
ik.Då	 ->1	
ik.En	 ->1	
ik.Eu	r->1	
ik.Fa	k->1	
ik.Fr	å->2	
ik.Fö	r->1	
ik.Ge	n->1	
ik.Ha	n->2	
ik.Hi	t->1	
ik.Hä	r->1	
ik.I 	d->1	
ik.Ja	g->1	
ik.Me	n->1	
ik.Re	f->1	
ik.Ri	k->1	
ik.Tv	ä->1	
ik.Vi	 ->3	
ik.Äv	e->1	
ik: v	i->1	
ik?He	r->1	
ik?Va	d->1	
ika E	U->1	
ika a	l->1	r->2	t->7	v->1	
ika b	e->11	i->1	r->2	y->1	
ika d	e->8	j->1	o->1	u->1	y->1	ä->1	
ika e	f->1	n->3	t->2	u->2	
ika f	a->4	o->4	r->3	ö->12	
ika g	e->3	i->1	r->3	ä->2	
ika h	a->2	i->1	u->1	å->1	ö->1	
ika i	 ->2	n->11	
ika k	a->4	o->3	u->3	
ika l	i->1	o->2	ä->6	ö->1	
ika m	e->8	i->2	y->2	å->3	ö->3	
ika n	a->8	o->1	å->1	
ika o	b->1	c->4	f->1	
ika p	a->3	l->2	o->5	r->2	u->1	
ika r	a->1	e->11	i->1	ä->1	ö->1	
ika s	a->1	i->1	j->2	k->3	l->2	p->1	t->6	v->1	y->1	ä->4	
ika t	a->1	e->2	i->2	o->1	y->3	
ika u	p->1	t->6	
ika v	a->4	e->1	i->9	ä->3	
ika ä	n->7	r->1	
ika å	t->4	
ika ö	p->1	v->2	
ika, 	e->1	f->3	o->2	s->2	v->1	
ika-o	l->1	
ika.D	e->1	
ika.I	 ->1	
ika.J	a->3	
ika.P	å->1	
ika.V	a->1	e->1	
ikabe	h->1	k->1	
ikada	n->2	
ikafr	å->1	
ikal 	f->1	o->1	p->1	
ikala	 ->8	.->1	
ikale	r->1	
ikali	e->5	s->1	
ikalt	 ->3	,->1	.->1	
ikaly	d->1	
ikan 	o->1	
ikand	e->6	
ikane	n->3	r->10	
ikans	k->11	
ikapa	c->1	
ikapi	t->1	
ikapp	,->1	.->1	a->3	
ikapr	o->1	
ikar 	m->1	r->1	s->1	v->1	
ikare	 ->3	,->1	
ikarn	a->5	
ikart	a->2	
ikas 	h->3	k->1	o->3	ä->2	ö->1	
ikas.	D->1	H->1	
ikasm	u->1	
ikast	e->3	
ikaså	 ->4	
ikat 	f->1	o->3	s->2	
ikat,	 ->1	
ikati	o->18	
ikato	r->5	
ike (	f->1	
ike -	 ->3	
ike a	g->1	t->2	
ike b	a->1	e->1	l->1	
ike d	å->1	
ike e	l->3	t->1	
ike f	ö->2	
ike g	e->2	
ike h	a->2	
ike i	 ->3	n->1	
ike k	o->3	
ike m	e->1	i->1	å->2	
ike n	a->1	
ike o	c->9	m->1	
ike s	o->6	ä->1	
ike t	i->1	
ike v	i->2	
ike ä	r->3	
ike, 	B->1	S->1	b->1	d->2	f->1	g->1	h->2	i->1	k->1	n->1	o->1	v->2	
ike. 	D->1	
ike..	 ->1	(->1	
ike.D	e->4	ä->1	
ike.F	r->1	ö->2	
ike.I	 ->1	
ike.J	a->2	
ike.M	e->1	
ike.N	i->1	
ike.O	m->1	
ike.V	i->3	
ike.Ö	s->1	
ike: 	i->1	
ikeEn	 ->1	
ikeFr	u->1	
ikeNä	s->1	
ikedo	m->10	
ikel 	1->16	2->13	3->8	4->8	5->6	6->12	7->8	8->16	9->3	s->2	ä->1	
ikel,	 ->2	
ikels	e->5	
iken 	(->1	-->2	1->2	J->1	K->3	S->2	T->3	b->1	e->3	f->14	g->1	h->4	i->12	k->4	l->1	m->8	n->2	o->10	p->2	r->1	s->8	t->2	v->2	y->1	Ö->1	ä->2	å->3	ö->1	
iken,	 ->21	
iken.	 ->1	A->1	B->1	D->9	E->3	F->2	H->1	I->1	J->5	K->1	P->1	S->1	V->1	
iken?	F->1	V->1	
ikenH	e->1	
ikens	 ->19	
iker 	a->4	b->3	d->1	f->3	h->2	i->1	k->1	m->2	o->3	p->1	s->2	v->1	ä->1	
iker,	 ->4	
iker.	B->1	
ikern	a->12	
ikers	 ->1	
ikes 	a->1	b->1	d->2	f->9	i->2	k->1	n->1	o->3	p->1	r->2	s->2	v->1	
ikes-	 ->4	
ikesf	r->4	
ikesh	a->4	
ikesm	i->9	
ikesp	o->3	
iket 	a->1	f->1	o->1	s->3	t->1	
iket,	 ->3	
iket.	M->1	S->1	
ikets	 ->6	
ikgil	t->2	
ikh h	a->1	
ikh-a	v->1	
ikh.D	e->1	
ikh.F	ö->1	
ikhet	 ->28	.->1	e->6	
ikisk	 ->5	a->42	e->2	
ikist	a->5	
ikit 	a->1	
ikiti	n->2	
iklar	,->3	.->1	n->11	
ikled	 ->1	
iklig	,->1	.->1	a->3	e->1	
ikmet	e->2	
ikna.	V->1	
iknan	d->19	
iknar	 ->2	
iknin	g->44	
iko, 	A->1	
ikolo	n->1	
ikomm	i->1	
ikomr	å->6	
ikont	r->2	
ikonv	e->1	
ikraf	t->4	
ikrat	i->1	
ikrav	 ->1	e->1	
ikrik	t->4	
ikrof	ö->1	
ikrok	r->2	
ikros	t->1	
ikryp	t->2	
iks m	å->1	
iksom	 ->55	
ikstä	l->2	
ikt -	 ->2	
ikt F	l->1	
ikt a	t->25	
ikt b	e->2	l->1	ä->1	
ikt d	a->1	e->1	ä->1	
ikt e	k->1	l->1	n->1	t->1	
ikt f	i->1	ö->4	
ikt g	å->1	ö->1	
ikt h	a->5	
ikt i	n->4	
ikt k	a->5	o->3	u->1	
ikt l	a->1	e->1	y->1	ä->1	
ikt m	e->4	o->1	
ikt o	c->7	m->6	
ikt p	å->2	
ikt r	e->1	
ikt s	a->1	k->4	o->6	t->1	ä->2	
ikt v	e->1	i->9	
ikt ä	m->1	n->1	r->5	v->2	
ikt ö	v->1	
ikt, 	d->1	e->2	g->1	i->1	l->1	m->2	o->2	t->1	v->1	ä->1	
ikt.B	å->1	
ikt.D	e->3	
ikt.I	 ->1	
ikt.J	a->1	
ikt.K	o->1	
ikt.O	c->1	m->2	
ikt.R	e->1	
ikt.V	a->1	
ikt; 	å->1	
ikta 	d->1	e->4	f->1	g->1	k->4	r->3	u->5	
ikta,	 ->1	
ikta.	J->1	
iktad	 ->5	.->2	e->12	
iktan	d->1	
iktar	 ->5	e->4	
iktas	 ->3	
iktat	 ->8	,->2	.->1	o->1	s->2	u->2	
ikte,	 ->2	
ikte.	F->1	
iktel	s->13	
ikten	 ->30	,->4	.->9	s->1	
ikter	 ->19	,->3	.->2	a->2	n->5	
iktfö	r->1	
iktig	 ->79	,->7	.->8	?->1	a->147	h->57	t->155	
iktio	n->9	
iktiv	 ->1	
iktli	g->4	n->74	
iktni	n->55	
iktpu	n->2	
iktsf	o->1	ö->2	
iktsm	e->1	
iktsp	l->1	
ikväl	 ->4	
ikvär	d->5	
ikäll	a->2	o->35	
il - 	f->1	
il -,	 ->1	
il 19	9->1	
il Po	l->1	
il el	l->3	
il en	e->1	
il fö	r->2	
il gr	a->1	u->1	
il i 	g->1	
il ko	s->1	
il me	d->2	
il nä	r->1	
il oc	h->1	
il so	c->1	m->4	
il sä	k->2	
il ut	a->2	
il ve	t->1	
il, s	i->1	
il, t	å->1	
il- o	c->2	
il-De	l->1	
il-Ro	b->1	
il-pr	o->1	
il. E	n->1	
il.De	n->1	t->1	
il.Ja	g->1	
il.Ly	n->1	
il.Tr	o->1	
ila b	l->1	r->2	
ila s	a->3	
ilaga	 ->1	.->1	n->2	
ilago	r->2	
ilags	t->1	
ilank	e->1	
ilar 	-->1	b->1	d->2	e->1	f->1	g->1	h->2	i->6	k->1	l->1	m->1	n->1	o->4	p->1	s->16	t->1	u->1	ä->2	å->1	
ilar,	 ->14	
ilar.	D->4	I->3	J->3	M->1	V->2	
ilar?	N->1	
ilarb	e->1	
ilare	 ->1	
ilarn	a->10	
ilate	r->9	
ilbef	o->2	
ilbes	t->1	
ilbra	n->1	
ild a	v->2	
ild b	e->3	
ild f	r->1	u->1	
ild i	n->1	
ild k	l->1	o->1	u->1	
ild m	a->1	e->1	
ild o	c->1	
ild p	e->1	
ild r	e->1	o->1	
ild t	a->1	o->1	
ild u	p->2	
ild, 	o->1	
ild.D	e->1	
ild.F	ö->1	
ild.N	u->1	
ilda 	b->1	d->2	e->4	f->5	i->3	k->2	l->2	m->4	n->1	p->2	r->3	s->7	t->1	v->1	ä->1	å->3	
ildad	e->3	
ildan	d->5	
ildar	 ->6	
ildas	 ->4	,->1	.->1	?->1	t->1	
ildat	 ->1	s->2	
ilde 	j->1	m->1	
ilde,	 ->1	
ilde.	E->1	
ildel	a->3	
ilden	 ->2	
ilder	 ->1	n->1	
ildni	n->66	
ildra	 ->3	r->1	t->2	
ileda	r->1	
ilege	.->1	?->1	
ilegi	e->3	u->1	
ilemm	a->3	
ilen 	b->1	i->1	u->1	
ilen,	 ->2	
ilen.	J->1	K->1	
ilera	s->1	
ilför	s->2	
ilhel	m->1	
ilia-	R->1	
ilien	.->1	
iligi	e->1	
ilikn	a->1	
ilind	u->30	
ilis 	f->1	
ilisa	t->1	
ilise	r->11	
ilism	.->1	
ilist	e->1	
ilita	r->2	
ilite	r->1	t->26	
ilitä	r->6	
ilj L	i->1	
ilja 	-->1	M->1	a->16	b->18	c->1	e->4	f->22	g->16	h->10	k->3	l->3	m->1	n->2	o->1	p->8	r->4	s->27	t->25	u->13	v->7	y->1	ö->1	
ilja,	 ->2	
ilja.	.->1	J->1	
iljad	e->3	
iljak	t->4	
iljan	 ->10	d->9	
iljar	 ->5	.->1	d->15	
iljas	 ->6	.->3	
iljat	 ->5	s->3	
ilje-	 ->1	
iljed	o->1	
iljef	a->1	ö->1	
iljej	o->3	
iljel	i->1	
iljem	ä->1	
iljer	 ->13	,->2	
iljes	t->1	
iljeå	t->1	
iljon	 ->1	e->63	t->1	
iljt 	u->1	
iljö 	f->2	i->1	k->1	m->1	s->2	v->1	
iljö!	D->1	
iljö,	 ->11	
iljö-	 ->2	
iljö.	D->3	M->1	U->1	V->1	
iljöa	n->3	v->1	
iljöb	e->3	r->1	
iljöd	e->1	i->1	
iljöe	r->4	
iljöf	a->2	r->4	ö->4	
iljöi	n->1	
iljök	a->11	o->6	r->8	v->1	
iljöl	a->1	
iljöm	i->1	ä->11	å->3	
iljön	 ->15	!->1	,->9	.->10	o->2	s->2	
iljöo	m->4	v->1	
iljöp	e->1	o->8	r->4	å->1	
iljör	å->1	ö->2	
iljös	e->1	i->1	k->15	t->1	y->6	
iljöu	t->1	
iljöv	ä->9	
ilka 	a->1	b->2	d->7	e->3	f->8	g->5	i->2	j->1	k->16	l->4	m->5	n->2	o->4	p->4	r->1	s->11	t->3	u->3	v->5	ä->9	å->7	ö->1	
ilkas	 ->2	
ilken	 ->54	,->1	
ilket	 ->180	
ilkon	s->1	
ilkyr	k->1	
ilköp	a->2	
ill "	M->1	
ill -	 ->2	
ill 1	0->1	5->1	9->3	
ill 2	 ->1	,->2	5->1	
ill 3	 ->1	0->1	
ill 4	 ->1	
ill 5	0->1	
ill 7	,->1	0->1	7->1	
ill 8	3->1	5->1	
ill 9	 ->1	1->1	4->2	
ill A	l->1	
ill B	a->1	o->2	r->2	
ill C	h->1	o->1	
ill D	i->1	
ill E	G->2	U->6	f->1	u->23	
ill F	r->3	ö->4	
ill G	e->1	r->1	
ill I	r->1	
ill K	a->2	i->2	o->8	u->1	
ill L	o->2	
ill M	c->1	i->1	o->2	
ill N	i->2	
ill O	L->1	
ill P	P->1	a->3	u->1	
ill R	a->1	
ill S	c->1	o->3	t->2	y->1	
ill T	h->1	i->1	r->1	y->2	
ill V	e->1	
ill W	a->2	i->1	u->1	
ill a	b->1	l->29	n->16	r->8	t->271	v->8	
ill b	a->11	e->35	i->3	l->1	o->4	r->4	u->1	y->2	ä->2	å->2	ö->10	
ill c	a->1	
ill d	a->1	e->253	i->22	o->4	r->2	ä->11	
ill e	f->2	g->3	k->1	l->1	m->3	n->104	r->13	t->30	u->1	x->45	
ill f	a->5	e->1	i->3	l->3	o->5	r->30	u->5	ä->2	å->1	ö->110	
ill g	a->4	e->15	i->1	l->1	o->7	r->17	ä->7	å->3	ö->4	
ill h	a->46	e->10	j->2	o->1	u->5	ä->3	ö->5	
ill i	 ->11	c->1	d->1	n->27	s->1	
ill j	a->97	o->1	u->3	ä->2	
ill k	a->6	l->3	n->1	o->56	r->3	u->1	v->1	ä->1	ö->1	
ill l	a->3	e->3	i->6	u->1	y->1	ä->3	å->2	
ill m	a->13	e->25	i->24	o->4	y->6	ä->1	å->4	ö->3	
ill n	a->9	i->2	o->1	u->1	y->9	ä->9	å->10	ö->2	
ill o	a->1	c->48	f->1	i->1	j->1	l->5	m->9	p->1	r->6	s->4	
ill p	a->8	e->5	i->1	l->1	r->13	u->1	å->11	
ill r	a->1	e->25	i->3	ä->8	å->19	ö->1	
ill s	a->8	e->7	i->32	j->6	k->21	l->15	m->2	n->1	o->3	p->2	t->56	u->5	v->2	y->6	ä->43	å->5	
ill t	a->34	e->2	i->10	o->1	r->7	u->1	v->6	y->1	
ill u	-->1	n->5	p->8	r->2	t->21	
ill v	a->22	e->10	i->39	o->1	ä->6	å->14	
ill y	r->2	t->3	
ill Ö	s->1	
ill ä	n->15	r->4	v->2	
ill å	r->2	t->10	
ill ö	k->2	n->1	s->1	v->1	
ill!H	e->1	
ill, 	a->1	d->1	e->2	f->1	h->1	i->2	k->1	m->3	n->2	o->6	r->1	s->1	u->1	v->1	å->1	
ill.A	v->1	
ill.D	e->4	ä->1	
ill.E	t->1	
ill.F	ö->1	
ill.H	e->2	
ill.I	 ->2	
ill.J	a->1	
ill.R	e->1	
ill.S	å->1	
ill.V	i->1	
ill: 	j->1	
ill?D	a->1	
ill?H	u->1	
ill?J	a->1	
illa 	b->1	d->1	k->1	m->2	o->4	
illa,	 ->2	
illar	 ->1	
illav	a->1	
illba	k->52	
illbr	i->4	
illde	l->12	
illdr	a->1	
ille 	a->1	f->3	g->1	h->1	p->1	t->1	u->1	v->3	
illeg	a->8	
illen	n->7	
iller	k->3	
illes	 ->1	
illfi	n->1	
illfo	g->6	
illfr	e->27	
illfä	l->97	
illfö	r->13	
illgo	d->1	
illgr	i->2	
illgä	n->21	
illgå	n->25	
illha	n->43	
illhe	t->2	
illhö	r->8	
illi!	J->1	
illig	 ->3	a->15	h->1	s->1	t->7	
illin	g->1	
illko	m->6	r->64	
illkä	n->9	
illmä	t->2	
illmö	t->3	
illna	d->44	
illni	n->1	
illnä	r->6	
illob	b->2	
illoj	a->2	
illol	j->1	
illor	 ->1	
illrä	c->75	t->2	
ills 	C->1	a->2	b->2	d->2	h->11	i->8	k->1	m->1	o->1	s->1	t->2	v->7	ä->2	å->1	
ills,	 ->2	
ills.	D->2	H->1	
ills?	V->1	
illsa	m->30	t->3	
illse	 ->13	
illsk	a->1	o->1	r->2	y->1	
illsl	u->1	
illst	å->22	
illsv	a->3	
illsä	t->4	
illta	 ->1	g->1	l->1	
illtr	o->1	ä->7	
illva	l->1	
illve	r->86	
illvi	d->1	l->1	
illvä	g->8	n->1	x->20	
illäg	g->18	n->2	
illäm	p->177	
illåt	 ->10	a->13	e->20	l->3	n->6	s->3	
ilmen	 ->1	
ilmer	 ->1	
ilmär	k->1	
ilo g	å->1	
ilo m	å->1	
ilo o	c->1	
ilo, 	s->1	
ilobb	y->1	
ilome	t->1	
iloso	f->5	
ilot 	i->1	
ilote	n->1	
ilotp	r->2	
ilovo	 ->1	
ilpar	k->6	
ilpro	d->1	
ilreg	e->1	
ilrät	t->1	
ils l	i->2	
ilse 	g->1	
ilsek	t->1	
ilsel	e->2	
ilska	 ->2	n->1	
ilskr	o->2	
ilsky	d->2	
ilskö	p->1	
ilspr	i->1	
ilsto	l->1	
ilt E	U->2	
ilt S	t->1	u->1	
ilt a	k->1	l->1	t->1	
ilt b	e->6	r->1	u->1	ö->1	
ilt d	e->7	
ilt e	f->1	n->1	t->1	
ilt f	a->2	r->2	ä->1	å->1	ö->8	
ilt g	e->2	l->1	ä->2	
ilt h	a->1	e->1	ä->1	
ilt i	 ->7	l->1	m->1	n->2	
ilt j	o->1	u->1	
ilt k	ä->3	
ilt l	y->1	
ilt m	e->7	y->1	ä->1	å->2	
ilt n	ä->4	ö->1	
ilt o	m->1	r->1	
ilt p	u->2	å->6	
ilt s	e->1	k->1	o->1	p->1	ä->2	
ilt t	a->2	i->6	r->1	y->3	
ilt u	p->3	t->1	
ilt v	a->4	i->11	å->2	
ilt ä	n->1	r->1	
ilt å	t->1	
ilt, 	o->1	
iltib	e->1	
iltig	 ->3	a->7	h->12	t->4	
iltil	l->17	
ilton	.->1	
iltre	r->1	
ilure	s->1	
ilver	 ->2	,->1	
ilvra	k->6	
iläga	r->1	
iläng	d->1	
ilåte	r->1	
ilöne	r->1	
ima f	r->1	
ima i	 ->1	
ima o	r->2	
ima s	t->1	
ima, 	m->1	
ima.H	e->1	
image	 ->1	
imagi	n->1	
imal 	e->1	f->1	s->1	
imala	 ->3	y->1	
imali	s->1	
imalt	 ->2	.->1	
imang	 ->1	e->2	
imat 	s->1	
imat.	D->1	
imate	t->7	
imatf	ö->4	
imatp	r->1	
imatu	m->1	
imbus	 ->1	
imen 	i->1	
imen.	J->1	
imens	 ->1	i->13	
iment	e->1	
imera	 ->3	r->3	s->1	y->1	
imeri	n->1	
imete	r->1	
imibe	s->2	
imifi	n->1	
imiin	n->1	
imika	p->1	
imiko	n->1	
imikr	a->2	
imilä	n->1	
imilö	n->1	
imina	l->4	
imine	l->3	r->23	
imini	v->1	
imino	r->2	
iminä	r->3	
imire	f->2	g->3	
imis-	n->1	
imist	i->6	
imite	t->6	
imiti	v->1	
imitr	a->5	
imixe	n->1	
imiål	d->1	
imlig	 ->4	a->6	e->1	t->12	
imma 	ä->1	
immar	 ->6	,->1	
immat	e->1	
imme 	e->1	o->2	s->2	
immig	r->6	
immun	i->1	
imoru	m->1	
imple	m->1	
impon	e->3	
impop	u->1	
impor	t->6	
impso	n->1	
impul	s->6	
imsav	t->2	
imsbe	t->2	
imsol	l->1	
imspa	r->1	
imsrå	d->2	
imsåt	g->1	
imt i	n->1	
imt o	m->2	
imt, 	f->1	
imula	n->4	t->2	
imule	r->7	
imum 	-->1	a->1	m->1	p->1	
imus-	b->1	
imynd	i->1	
imål,	 ->1	
imöge	l->1	
in - 	t->1	
in 19	4->1	
in 26	 ->1	
in Eu	r->1	
in Fr	a->1	
in ab	s->1	
in ak	t->1	
in an	d->5	s->2	
in ar	b->2	
in at	t->4	
in av	s->4	
in ba	k->1	
in be	d->2	f->3	h->1	r->1	s->1	u->1	
in bi	d->1	l->5	
in bl	a->1	
in br	o->1	ä->1	
in bu	d->2	
in da	g->2	
in de	l->7	m->1	n->2	t->3	
in dj	u->2	
in do	m->1	
in dr	a->1	
in eg	e->10	
in ek	o->3	
in en	d->1	e->2	
in er	f->2	
in et	t->2	
in ex	a->1	i->1	
in fa	k->1	
in fo	r->1	
in fr	e->1	u->1	å->17	
in fu	n->1	
in fy	r->1	
in få	r->1	
in fö	d->1	r->20	
in ge	m->1	
in gl	ä->2	
in go	d->1	
in gr	u->30	
in ha	d->1	r->5	
in he	l->10	m->2	
in hu	n->1	
in hä	n->1	v->1	
in hö	j->2	
in i 	E->2	H->1	K->1	M->1	a->3	b->1	d->4	e->5	f->4	h->1	i->1	o->1	r->1	t->3	u->1	v->1	ä->1	å->1	
in i,	 ->1	
in in	i->1	o->2	s->1	t->1	v->1	
in ka	m->1	n->1	t->1	
in ko	l->25	m->4	n->3	
in kr	ä->1	
in kä	r->1	
in li	k->1	n->2	v->1	
in lö	p->1	
in ma	k->2	r->1	s->1	
in me	d->3	n->15	r->2	
in mo	r->1	t->2	
in må	n->3	
in na	t->5	
in nu	v->2	
in ny	n->1	
in nä	r->2	
in ob	e->1	
in oc	h->34	
in or	d->4	g->1	o->1	
in os	s->1	
in pa	r->1	
in pe	n->1	r->3	
in pl	a->3	i->1	
in po	l->3	t->1	
in pr	e->1	o->1	
in på	 ->23	:->1	s->1	
in ra	p->2	
in re	a->1	g->3	s->2	
in ri	s->2	
in ro	l->6	
in rä	t->5	
in rö	s->6	
in se	d->1	
in si	g->2	n->1	s->3	t->1	
in sj	ä->2	
in sk	a->2	u->2	
in sl	u->2	
in so	 ->1	l->4	m->13	
in sp	e->2	o->1	
in st	a->1	o->2	r->1	ä->3	å->1	
in su	v->1	
in sy	n->2	
in sä	k->1	t->1	
in så	 ->2	n->1	
in ti	d->1	l->3	
in tr	e->3	
in tu	r->6	
in un	d->4	
in up	p->19	
in ut	a->1	b->2	f->2	k->1	v->1	
in va	l->2	r->2	
in ve	t->1	
in vi	l->3	t->1	
in vu	n->1	
in vä	g->1	n->1	
in vå	r->2	
in we	b->1	
in yt	t->1	
in än	d->1	
in är	 ->2	
in ås	i->12	
in ön	s->4	
in!He	r->1	
in", 	d->1	
in, d	å->1	
in, e	f->1	
in, f	l->1	ö->2	
in, g	e->1	j->1	
in, h	a->2	
in, m	e->2	i->1	
in, o	c->6	m->1	
in, p	u->1	å->1	
in, r	a->1	
in, s	o->4	å->1	
in, t	.->1	
in, u	t->1	
in, v	i->2	
in-rå	d->3	
in. D	e->1	
in. M	e->1	
in.Al	l->1	
in.Be	d->1	
in.Ce	n->1	
in.De	t->5	
in.Dä	r->1	
in.Fö	r->2	
in.He	l->1	r->1	
in.In	g->1	
in.Ja	g->3	
in.Li	v->1	
in.Lå	t->1	
in.Me	n->1	
in.Nä	r->1	
in.Om	 ->2	
in.Sa	m->1	
in.Sc	h->1	
in.St	å->1	
in.Va	r->1	
in.Vi	 ->4	
in: e	n->1	
in?Pa	r->1	
ina a	f->1	k->1	n->3	r->1	t->3	v->1	
ina b	a->1	e->4	i->2	r->1	
ina d	a->38	o->2	
ina e	g->15	k->1	l->1	r->1	
ina f	a->3	e->1	i->2	o->1	r->2	ö->9	
ina g	a->2	o->1	r->6	
ina h	a->1	e->1	ä->2	å->3	
ina i	n->9	
ina j	o->1	
ina k	o->24	ä->5	
ina l	a->1	i->1	o->1	ä->1	ö->1	
ina m	e->6	i->1	å->1	
ina n	a->3	
ina o	c->5	f->1	l->1	m->1	r->1	
ina p	r->1	
ina r	a->1	e->8	i->2	ä->1	å->2	ö->2	
ina s	e->2	k->3	l->4	o->3	p->1	t->3	y->2	ö->1	
ina t	a->3	e->1	i->2	j->2	r->1	
ina u	n->2	p->6	t->2	
ina v	a->1	e->1	i->1	ä->4	
ina y	r->1	
ina ä	n->2	r->1	
ina å	r->1	t->2	
ina ö	g->1	n->1	v->1	
ina, 	o->1	
ina-I	s->1	
ina.H	e->1	
ina.U	n->1	
inafl	y->1	
inafr	å->1	
inal 	i->1	
inale	r->3	
inali	s->4	t->1	
inalp	o->1	
inalv	e->1	
inans	 ->1	d->1	e->2	i->79	m->1	
inarb	e->1	
inari	u->1	
inas 	l->1	r->1	
inati	o->8	
inavi	s->1	
inban	a->1	
inbeg	r->12	
inbju	d->6	
inbjö	d->1	
inbla	n->14	
inbur	g->1	
inbyg	g->1	
incid	e->1	
incip	 ->28	,->3	.->4	e->150	i->8	s->1	
incit	a->8	
ind o	c->1	
inda 	b->1	p->1	ö->1	
inda.	D->1	I->1	
indan	d->12	
inde 	o->1	
indel	a->2	n->1	s->15	
inden	 ->1	
inder	 ->32	,->3	.->7	
indfä	l->4	
indik	a->6	
indir	e->7	
indis	k->1	
indiv	i->14	
indra	 ->29	d->3	n->2	r->9	s->7	t->3	
indre	 ->51	.->1	?->1	n->3	
indrä	n->2	
indus	t->113	
ine d	i->1	
ine f	ö->1	
ine h	a->1	
ine n	ä->1	
ine q	u->2	
ine, 	d->1	
ineff	e->3	
inell	 ->1	a->3	
inen 	f->2	h->1	i->1	
inen,	 ->3	
inens	 ->2	
inent	,->1	.->1	a->2	e->1	
iner 	b->1	f->1	g->1	i->2	n->1	o->1	ä->1	
inera	 ->7	d->3	n->5	s->2	
ineri	e->1	n->30	
inern	a->1	
inese	r->2	
inesi	s->7	
inett	 ->1	.->1	e->1	
inez 	a->1	
infek	t->2	
infil	t->1	
infin	i->1	n->1	
infly	t->12	
infor	d->2	m->90	
infra	s->15	
infri	a->1	
infrå	g->1	
inför	 ->71	,->1	.->2	:->1	a->55	d->3	l->19	s->6	t->6	
ing (	1->1	E->1	a->2	r->1	å->1	
ing -	 ->10	,->1	
ing 1	7->1	9->1	
ing 2	0->2	
ing 3	7->1	
ing 6	0->1	8->1	
ing 8	0->2	
ing D	e->1	
ing E	c->1	u->1	
ing F	ä->1	
ing I	V->2	
ing T	a->1	
ing V	I->1	
ing a	l->2	n->7	t->26	v->324	
ing b	a->2	e->2	i->1	l->3	o->1	r->1	ö->4	
ing d	e->5	y->1	ä->6	
ing e	.->1	f->2	l->8	n->4	t->5	x->2	
ing f	i->4	o->1	r->27	u->1	å->1	ö->77	
ing g	a->1	e->6	j->1	r->1	å->1	
ing h	a->17	o->3	ä->1	å->1	
ing i	 ->85	a->1	n->30	
ing k	a->5	n->1	o->14	r->2	u->1	
ing l	e->1	i->4	ä->2	å->1	
ing m	a->4	e->43	i->2	o->10	å->11	
ing n	e->1	i->2	r->2	u->1	ä->3	ö->1	
ing o	c->137	f->2	m->34	
ing p	l->1	r->1	å->51	
ing r	a->1	e->1	ä->2	ö->2	
ing s	a->2	e->1	i->1	k->16	o->104	t->4	y->1	ä->2	å->4	
ing t	a->5	i->44	r->2	y->1	
ing u	n->4	t->8	
ing v	a->8	e->2	i->15	
ing ä	g->1	n->6	r->31	v->2	
ing å	t->4	
ing ö	v->2	
ing!J	a->1	
ing" 	a->1	o->1	
ing",	 ->2	
ing".	J->1	
ing) 	i->2	o->2	
ing).	V->1	
ing)N	ä->1	
ing, 	O->1	a->5	b->3	d->13	e->13	f->24	g->2	h->4	i->12	k->5	l->3	m->17	n->7	o->19	p->6	r->1	s->28	t->4	u->8	v->13	ä->4	å->3	ö->1	
ing-P	M->1	
ing. 	D->2	E->1	M->1	
ing.(	A->1	
ing..	 ->1	(->1	
ing.A	l->3	n->1	v->4	
ing.D	a->1	e->58	o->2	ä->4	
ing.E	f->1	n->4	t->1	u->1	
ing.F	l->1	r->4	ö->10	
ing.G	e->2	
ing.H	a->1	e->12	ä->1	
ing.I	 ->12	n->2	
ing.J	a->29	
ing.K	a->1	o->8	
ing.L	i->1	å->2	
ing.M	a->6	e->4	y->1	å->2	
ing.N	a->1	i->3	u->1	ä->1	å->1	
ing.O	c->4	f->1	m->8	
ing.P	P->1	a->1	r->1	å->2	
ing.R	e->1	
ing.S	a->1	e->1	l->4	å->1	
ing.T	a->1	i->2	
ing.V	a->1	i->15	å->1	
ing.Ä	r->2	
ing: 	e->1	f->1	i->1	
ing:D	e->1	
ing; 	d->1	e->1	f->2	
ing?D	e->2	
ing?H	ä->1	
ing?J	a->1	
ing?O	l->1	
ing?T	y->1	
ing?Ä	r->1	
inga 	a->1	b->3	d->3	f->2	g->1	i->1	k->2	m->4	n->2	o->3	p->1	r->5	s->5	t->1	u->2	v->3	ä->1	
inga.	V->1	
ingad	e->6	
ingal	u->3	
ingan	d->8	
ingar	 ->295	!->1	"->1	)->1	,->46	-->1	.->74	:->7	;->1	n->142	s->3	
ingas	 ->10	.->1	
ingat	 ->3	s->1	
ingdy	r->1	
ingel	ä->1	
ingen	 ->682	"->1	,->71	.->90	:->4	;->2	?->7	j->2	s->21	t->21	
inger	 ->2	,->1	
inget	 ->33	
ingfl	ö->1	
ingfo	n->1	r->20	
inggå	 ->1	s->1	
ingiv	i->6	
ingom	 ->3	.->1	
ingpo	l->2	
ingra	 ->2	
ingre	d->2	p->5	s->1	
ingri	n->1	p->9	
ings 	b->1	d->1	h->1	p->1	v->1	
ings-	 ->12	
ingsa	k->3	l->1	n->7	r->5	v->6	
ingsb	a->2	e->7	i->11	o->3	
ingsc	e->5	h->8	
ingsd	i->2	o->1	r->1	
ingse	n->1	r->1	t->1	
ingsf	a->7	e->2	i->30	l->1	o->22	r->15	u->11	ö->232	
ingsg	r->6	
ingsh	a->1	o->1	
ingsi	d->1	n->10	
ingsk	a->1	l->3	o->170	r->14	u->1	v->1	
ingsl	a->1	i->58	o->1	ä->6	ö->5	
ingsm	a->4	e->7	i->1	o->5	ä->2	å->4	ö->4	
ingsn	i->5	o->1	y->1	
ingso	m->10	r->2	
ingsp	a->4	l->23	o->21	r->45	å->1	
ingsr	e->18	u->1	ä->2	å->1	
ingss	a->2	e->4	i->2	k->14	p->1	t->18	y->22	ä->9	
ingst	a->7	e->1	j->5	ä->1	
ingsu	m->1	t->6	
ingsv	e->4	i->33	ä->7	å->1	
ingsä	r->1	
ingså	r->1	t->5	
ingsö	v->1	
ingto	n->5	
ingtv	ä->4	
ingå 	e->1	i->5	s->2	
ingå.	A->1	
ingåe	n->5	
ingån	g->1	
ingår	 ->11	.->2	
ingåt	t->6	
inhem	s->2	
inho 	f->1	p->1	s->1	v->1	
inho.	 ->1	
inhos	 ->1	
inhäm	t->6	
inier	a->12	i->1	n->4	
inifr	å->1	
inima	l->1	
inime	r->1	
inimi	b->2	f->1	i->1	k->4	l->2	n->3	r->5	s->1	
inimo	r->1	
inimu	m->4	s->1	
ining	s->1	
inion	 ->2	e->1	s->1	
inipe	n->1	
inire	f->1	
inist	e->55	i->3	r->41	
initi	a->77	e->2	o->14	v->9	
initu	m->1	
inivå	,->1	
inje 	(->1	m->5	o->1	s->4	
inje.	G->1	J->1	
injen	 ->2	.->1	
injer	 ->36	"->1	,->5	.->3	:->1	n->31	
inkel	 ->6	.->3	n->2	
inkla	r->1	
inklu	d->4	s->17	
inkom	p->3	s->10	
inkon	s->1	v->2	
inkri	s->1	
inkrä	k->1	
inkte	r->1	
inkti	o->1	v->1	
inköp	 ->1	s->1	
inkör	s->1	
inlan	d->6	
inled	a->31	d->10	e->6	n->8	s->5	
inlet	t->13	
inlig	h->1	
inläg	g->18	
inläm	n->5	
inlän	d->5	
inlås	t->1	
inlåt	a->1	
inlöp	a->1	
inmäs	s->1	
inna 	-->1	a->1	b->1	d->4	e->9	f->2	h->2	i->2	k->2	l->2	m->3	n->1	o->19	p->4	r->1	s->5	t->1	v->3	
inna,	 ->1	
inna.	 ->1	
innan	 ->39	
innas	 ->46	!->1	,->1	.->2	
innat	 ->1	
inne 	a->2	f->1	h->1	n->1	o->1	p->2	s->1	
inne,	 ->5	
inne.	D->1	
inneb	a->1	o->1	ä->108	ö->6	
innef	a->6	
inneh	a->3	å->77	ö->4	
innel	a->1	
innen	 ->1	.->1	a->1	
inner	 ->59	,->3	.->3	l->2	s->2	
innes	 ->1	m->1	r->1	
innet	.->2	
innev	å->2	
innig	h->1	
innin	g->49	
innli	g->2	
innoc	k->24	
innop	r->2	
innor	 ->36	,->3	.->4	?->1	n->5	s->10	
innov	a->6	
inns 	2->1	G->1	S->1	a->15	b->5	c->1	d->57	e->51	f->24	g->4	h->5	i->43	j->2	k->3	l->1	m->19	n->19	o->9	p->8	r->10	s->15	t->14	u->1	v->4	y->2	ä->3	å->1	ö->2	
inns,	 ->3	
inns.	D->3	J->1	M->1	V->1	
ino i	 ->1	
ino k	o->1	
ino o	m->1	
ino, 	T->1	m->1	
ino.J	a->1	
ino.O	r->1	
inom 	5->1	E->33	F->1	G->1	I->1	L->1	S->1	V->1	a->6	b->3	d->43	e->16	f->7	g->8	h->3	i->4	j->3	k->23	l->3	m->7	n->2	o->9	p->2	r->55	s->11	t->5	u->16	v->12	å->1	ö->4	
inome	u->1	
inori	t->22	
inorm	e->2	
inorn	a->1	
inos 	h->1	i->1	o->1	
inos,	 ->2	
inott	i->1	
inprä	n->1	
inra 	k->1	o->10	
inrar	 ->1	
inras	 ->1	
inre 	a->2	e->2	g->1	m->68	v->9	
inres	a->4	
inrik	e->13	t->44	
inrym	s->1	
inrät	t->55	
inråd	e->1	
ins a	b->1	k->1	l->1	r->1	
ins d	ö->1	
ins f	y->1	
ins i	n->2	
ins j	u->1	
ins k	o->2	
ins l	i->1	
ins p	r->1	
ins r	a->1	
ins s	a->1	e->1	l->1	t->1	
ins t	e->1	
ins v	a->1	
ins å	t->1	
insam	l->8	
insat	s->41	
insbu	t->1	
inse 	a->7	d->2	h->1	v->3	
inse;	 ->1	
insee	n->1	
insem	e->3	
inser	 ->23	,->1	n->1	
insik	t->4	
insis	t->6	
insk 	b->1	s->1	
inska	 ->35	,->1	.->2	d->6	n->2	r->7	s->1	t->7	
inskn	i->16	
inskr	i->2	ä->11	
insla	g->6	
inspe	k->12	
inspi	r->3	
inst 	-->1	1->2	3->2	4->1	a->1	b->1	d->2	f->1	i->1	l->1	m->2	n->1	o->1	p->2	r->1	s->4	u->2	v->2	
inst,	 ->1	
insta	 ->5	l->1	n->31	
inste	r->8	
insti	n->3	t->135	
instm	a->1	
insto	n->27	
instr	e->8	u->53	
insts	v->1	
instä	l->25	m->23	
insyn	 ->7	,->1	.->3	e->2	
int b	a->1	
int-E	x->1	
inta 	d->1	e->3	
intag	a->1	i->4	
intar	 ->4	
inte 	-->3	1->1	B->1	E->3	a->138	b->140	c->1	d->56	e->55	f->119	g->74	h->163	i->47	j->1	k->102	l->65	m->60	n->49	o->32	p->45	r->35	s->103	t->72	u->49	v->50	ä->84	å->6	ö->12	
inte!	D->1	M->1	
inte,	 ->13	
inte.	A->1	B->1	D->3	H->2	J->2	S->1	V->2	Å->2	
inte:	 ->1	
inte?	F->1	H->1	
integ	r->42	
intel	l->8	s->5	
inten	s->12	t->1	
inter	i->16	n->82	p->1	v->10	
intet	 ->2	
intim	t->1	
intli	g->10	
intog	 ->2	
intol	e->4	
inton	s->1	
intre	s->120	
intro	d->6	
intry	c->15	
inträ	d->2	f->26	
intrå	n->1	
intyg	 ->1	a->3	
intäk	t->5	
inuc 	s->1	
inuer	l->2	
inus 	2->1	f->1	t->1	
inusg	r->2	
inut 	f->2	n->1	
inut.	(->1	)->1	J->1	
inute	r->10	
inval	d->1	
invan	d->18	
invec	k->2	
inven	t->1	
inver	k->7	
inves	t->15	
invit	 ->1	
invol	v->9	
invän	d->11	t->2	
invån	a->9	
inz F	l->2	
inär 	m->1	
inära	 ->8	
inäre	r->1	
inärf	r->1	
inärp	e->1	
inöva	d->1	
io Sá	n->1	
io Va	l->3	
io Vi	t->1	
io be	s->2	
io fa	t->1	
io fö	r->3	
io gr	a->1	
io gå	n->2	
io ha	r->1	
io lä	n->1	
io mi	l->6	n->1	
io må	n->2	
io pu	n->1	
io sa	f->1	
io si	n->1	
io sk	i->1	
io så	 ->1	
io ti	m->1	
io ut	t->1	
io än	d->1	
io år	 ->4	,->1	e->2	
io, a	n->1	
io, s	o->1	
io, t	i->1	
io-Pl	a->4	
io.Ja	g->1	
io.Nä	r->1	
io: v	i->1	
io; d	e->1	
iod a	v->2	
iod d	e->1	ä->1	
iod f	i->2	å->1	ö->1	
iod i	 ->3	n->1	
iod k	o->1	
iod o	m->1	
iod p	å->2	
iod r	e->1	ö->1	
iod s	o->2	
iod v	i->1	
iod ä	r->2	
iod, 	e->1	f->1	m->1	n->1	v->1	
iod.D	e->1	
iod.V	i->1	
iod?-	 ->1	
ioden	 ->31	,->2	.->4	s->2	
ioder	 ->1	n->1	
iodis	k->14	
ioeko	n->3	
ioelv	a->1	
iofem	 ->1	
ioför	k->1	
iogra	f->1	
iola 	v->1	
iolog	i->6	
ion (	A->5	
ion -	 ->3	
ion 1	2->5	
ion 5	2->1	
ion A	c->1	
ion H	a->1	
ion I	 ->1	
ion P	r->2	
ion a	l->1	n->1	p->1	t->4	v->18	
ion b	e->3	o->1	ö->1	
ion d	ä->8	
ion e	l->1	n->3	
ion f	r->5	u->1	å->1	ö->17	
ion g	e->3	r->1	å->1	
ion h	a->3	o->1	ä->3	ö->1	
ion i	 ->22	n->7	
ion j	a->1	
ion k	a->6	o->3	
ion m	e->12	o->2	y->1	
ion n	i->1	ä->2	
ion o	c->33	m->19	v->1	
ion p	å->9	
ion r	e->1	
ion s	a->1	k->8	o->49	p->1	t->2	ä->1	å->2	
ion t	a->2	i->17	y->1	
ion u	n->1	p->3	t->2	
ion v	e->1	i->5	å->1	
ion ä	n->1	r->5	
ion å	t->2	
ion" 	p->1	
ion) 	(->2	
ion, 	L->1	S->1	b->2	d->3	e->5	f->2	h->1	i->2	k->3	m->3	n->2	o->8	p->1	s->7	t->1	u->1	v->2	ä->3	
ion. 	I->1	O->1	R->1	
ion.1	4->1	
ion.B	r->1	
ion.D	E->1	e->14	ä->2	å->1	
ion.E	n->1	v->1	
ion.F	l->1	r->1	ö->3	
ion.G	ä->1	
ion.H	a->1	e->4	
ion.I	 ->6	
ion.J	a->10	
ion.K	o->2	
ion.M	i->2	ö->1	
ion.N	i->1	
ion.O	m->2	
ion.S	a->1	e->1	o->2	å->1	
ion.T	i->1	r->1	
ion.U	n->1	
ion.V	a->2	i->9	
ion.Å	 ->1	
ion: 	D->1	a->1	i->1	
ion; 	v->1	
ion? 	I->1	
ion?D	e->1	
ion?J	a->1	
ion?K	a->1	o->1	
ion?Ä	v->1	
ional	 ->8	-->2	.->1	a->44	e->4	f->2	i->28	l->1	p->37	r->1	s->6	t->1	
ionde	 ->1	n->1	
ionel	l->275	
ionen	 ->875	!->1	"->1	)->1	,->103	.->136	:->1	;->3	?->4	J->2	s->375	
ioner	 ->195	,->35	.->40	?->4	N->1	a->8	i->11	l->2	n->176	s->4	
ionis	m->3	t->2	
ionjä	r->1	
ions 	i->1	s->1	
ions-	 ->4	
ionsa	f->2	n->1	r->8	v->1	
ionsb	o->1	r->1	
ionsd	i->1	o->1	ö->1	
ionsf	o->1	r->2	u->1	ö->19	
ionsh	a->1	i->8	
ionsi	n->1	
ionsk	a->2	o->5	r->1	u->6	
ionsl	e->11	ä->1	
ionsm	e->4	o->1	ä->1	ö->1	
ionsn	i->2	
ionso	r->1	
ionsp	l->2	o->3	r->6	
ionsr	e->3	o->1	ä->12	
ionss	a->7	c->1	e->1	k->1	t->2	y->5	
ionst	e->2	j->1	
ionsu	n->3	p->1	t->3	
ionsv	i->1	
ionsä	m->1	
ionär	 ->65	!->32	,->74	.->11	e->65	s->1	
iopie	n->3	
iopla	s->1	
ior.D	e->1	
iorga	n->2	
iori 	o->1	s->1	v->1	
iorit	e->36	
ios i	n->1	
ios å	s->1	
iosfä	r->1	
iosju	 ->1	
iosäk	e->2	
iot i	 ->1	
iot s	o->1	
iotal	e->1	s->5	
iotek	e->2	
iotis	k->1	
iotus	e->1	
ioxid	 ->4	u->1	
ioxin	 ->1	k->1	
ip al	l->1	
ip at	t->2	
ip el	l->1	
ip en	 ->1	l->1	
ip fö	r->1	
ip i 	S->1	h->1	
ip in	o->1	t->4	
ip me	l->1	
ip oc	h->2	
ip om	 ->2	
ip rå	d->1	
ip so	m->4	
ip så	v->1	
ip är	 ->3	
ip äv	e->1	
ip, g	e->1	
ip, m	e->1	
ip, o	c->1	
ip.Ja	g->1	
ip.Sj	ä->1	
ip.Vi	 ->1	s->1	
ipa a	t->1	
ipa d	e->2	ä->1	
ipa e	k->1	n->1	
ipa i	 ->2	n->1	
ipa m	ä->1	
ipa o	c->1	r->1	
ipa p	å->1	
ipa r	ä->2	
ipa t	a->2	
ipa, 	t->1	
ipa.E	f->1	
ipa.K	o->1	
ipand	e->20	
ipara	g->1	
ipas 	o->1	
ipen 	"->1	a->3	b->4	f->2	g->1	h->6	i->8	k->1	m->3	n->2	o->24	p->2	s->4	t->2	v->1	ä->8	å->1	
ipen,	 ->11	
ipen.	.->1	D->5	E->1	J->4	P->1	S->2	T->1	V->1	Ä->1	
ipen:	 ->2	
ipenN	ä->1	
ipend	i->1	
iper 	a->1	d->2	e->3	f->5	i->3	l->1	m->2	o->7	p->2	s->11	t->1	u->2	ä->3	
iper,	 ->4	
iper.	F->2	O->1	V->2	
iper:	 ->1	
ipern	a->10	
ipes 	r->1	
ipet 	d->1	e->1	
ipet,	 ->1	
ipiel	l->8	
ipit 	o->1	s->1	
iplan	e->1	
iplig	 ->1	,->1	t->4	
iplin	 ->4	,->1	e->3	f->1	r->1	ä->4	
iplom	a->11	
ipna 	p->1	
ipnin	g->9	
ipoli	t->4	
ipote	n->1	
ippad	e->3	
ipper	 ->2	
iprod	u->3	
iprog	r->4	
ips a	v->1	
ipskä	l->1	
ique 	k->1	
iques	 ->1	"->1	
iquit	a->1	
ir Eu	r->2	
ir al	l->3	
ir an	s->1	t->1	
ir at	t->4	
ir av	 ->1	
ir bi	n->1	
ir br	e->1	
ir bä	t->1	
ir de	 ->1	n->3	s->1	t->7	
ir di	p->1	r->1	
ir en	 ->7	
ir et	t->3	
ir fo	r->1	
ir fr	a->1	i->1	
ir fö	r->3	
ir gr	u->1	
ir ha	l->1	
ir hj	ä->1	
ir ho	m->1	
ir i 	f->1	s->1	
ir in	d->1	g->1	o->1	
ir ja	g->1	
ir ju	 ->1	
ir ko	n->1	
ir la	g->1	
ir le	g->1	
ir lu	f->1	
ir lä	t->2	
ir me	n->1	r->3	
ir mi	n->1	
ir my	c->2	
ir må	n->1	
ir mö	j->3	
ir na	t->1	
ir ne	g->1	
ir nå	g->2	
ir nö	d->1	
ir of	u->1	
ir on	ö->1	
ir ot	å->1	
ir ou	t->1	
ir ra	t->1	
ir re	s->1	
ir rä	d->1	
ir sa	m->2	
ir se	k->1	n->1	
ir sk	y->1	
ir so	m->1	
ir st	u->1	ä->1	å->1	
ir sv	å->2	
ir sä	k->1	
ir så	 ->1	
ir ti	l->4	
ir tä	t->1	
ir ut	f->1	k->1	
ir va	l->1	
ir ve	r->2	
ir vi	 ->1	
ir än	d->1	
ir ås	k->1	
ir öv	e->1	
ir, g	e->1	
ir, i	n->1	
ir: O	m->1	
ira R	o->1	
ira m	e->1	
ira ä	r->1	
ira, 	i->1	o->1	
ira.J	a->1	
irake	l->1	
iraki	s->1	
irar 	o->1	
irare	 ->1	
irarn	a->1	
irate	r->1	
ire h	a->1	
ire, 	A->1	
ire-A	t->1	
ire.D	e->1	
irefo	r->4	
iregl	e->3	
irekt	 ->37	.->2	a->5	i->194	o->18	ö->1	
irer.	E->1	
irera	s->1	t->2	
irgiz	i->5	
irige	r->1	
irka 	1->1	e->1	h->1	t->1	
irkel	 ->1	
irkes	f->1	l->2	
irkla	r->2	
irkul	a->1	e->2	
irlän	d->11	
irman	 ->1	
irmou	t->1	
ironi	s->2	
irra 	s->1	
irrad	 ->1	e->1	
irran	d->1	
irrat	.->1	i->2	
irrep	a->1	
irrgå	n->1	
irrin	g->8	
irrit	a->1	e->3	
irrva	r->1	
irtan	d->1	
is (P	P->1	
is - 	m->1	n->1	s->1	
is Al	g->1	
is Ba	r->1	
is Go	l->1	
is Mi	t->1	
is Pa	c->1	
is Wu	r->1	
is al	l->3	
is an	a->1	i->1	p->1	v->2	
is at	t->13	
is av	 ->5	v->1	
is ba	r->1	s->1	
is be	h->3	k->1	
is br	a->1	y->1	
is bå	d->1	
is de	 ->2	f->1	l->1	n->3	t->5	
is dä	r->2	
is el	l->2	
is en	 ->4	
is et	t->2	
is ex	i->1	
is fi	n->2	
is fo	r->2	
is fr	a->1	å->3	
is fu	l->2	
is fy	l->1	
is få	r->2	
is fö	l->1	r->7	
is ge	n->2	
is go	d->3	
is gr	ä->1	
is gä	r->1	
is gå	 ->1	r->1	
is ha	 ->1	n->1	r->8	
is he	l->1	
is hj	ä->1	
is ho	p->1	
is hä	r->2	
is hö	g->1	
is i 	E->1	d->1	e->2	f->1	h->1	s->1	
is il	l->1	
is in	f->1	l->1	n->3	o->1	r->1	s->1	t->12	
is ju	s->2	
is ka	n->2	
is ke	m->1	
is ko	m->1	n->4	
is la	g->1	n->1	
is le	d->1	
is li	k->5	l->1	
is lo	v->1	
is me	d->2	n->1	r->1	
is mi	l->1	n->2	
is my	c->1	
is må	n->1	s->3	
is nä	m->1	r->2	
is oa	c->1	
is oc	h->4	k->14	
is om	 ->3	f->1	s->1	
is or	i->1	
is ot	r->1	
is pe	l->1	n->1	
is po	l->1	
is pr	i->1	o->1	
is på	 ->8	p->2	
is ra	s->1	
is re	d->1	
is ro	,->1	
is rä	k->1	
is sa	k->1	m->2	
is se	 ->1	
is si	d->1	
is sj	ä->1	
is sk	a->3	i->1	u->6	ö->1	
is sm	å->1	
is so	m->25	
is st	e->1	ä->2	ö->1	
is sv	å->1	
is sä	g->1	r->1	
is så	 ->3	
is ta	 ->1	
is te	k->1	
is ti	l->2	
is un	d->2	
is up	p->2	
is ut	i->1	m->1	v->2	
is va	d->1	r->1	
is vi	k->1	l->6	s->1	
is vä	c->1	g->2	l->1	
is än	n->2	
is är	 ->15	
is äv	e->4	
is ås	t->1	
is åt	 ->1	e->1	g->1	
is öv	e->3	
is! V	a->1	
is) f	ö->1	
is, E	v->1	
is, a	n->1	t->1	
is, d	e->2	i->1	v->1	
is, e	u->1	
is, i	 ->1	
is, k	o->2	
is, m	e->2	
is, n	ä->1	
is, o	c->3	
is, p	å->1	
is, s	o->1	å->1	
is, t	i->1	
is, v	a->1	
is-Jø	r->2	
is-fö	r->1	
is-no	t->1	
is-pr	o->1	
is. M	e->1	
is.Da	g->1	
is.De	s->1	t->1	
is.Då	 ->1	
is.Ef	t->1	
is.Fö	r->2	
is.Hu	r->1	
is.Ja	g->2	
is.Me	n->1	
is.Sa	m->1	
is.Se	d->1	
is.Vi	 ->1	
is.Än	d->1	
is: f	ö->1	
is; a	t->1	
is?Är	 ->1	
isa (	a->1	
isa R	y->1	
isa a	l->1	r->1	t->5	
isa b	e->1	ö->1	
isa d	e->4	
isa e	f->1	r->1	
isa f	ö->2	
isa g	r->1	
isa h	u->1	ö->1	
isa i	 ->5	n->3	
isa k	o->1	
isa l	i->1	
isa m	e->1	
isa o	c->1	m->1	s->1	
isa p	r->1	å->3	
isa s	i->7	o->1	t->1	
isa t	i->9	o->1	
isa u	t->1	
isa v	a->2	e->1	å->1	
isa ä	r->3	
isa, 	b->1	f->1	h->1	m->2	o->1	s->1	å->1	
isa..	.->1	
isa.B	a->1	
isa.D	e->3	ä->1	
isa.E	u->1	
isa.F	r->1	
isa.J	a->1	
isa.K	ä->1	
isa.R	å->1	
isa.S	a->1	
isa.U	p->1	
isa.Å	r->1	
isa?P	r->1	
isabe	t->1	
isade	 ->16	s->3	
isaka	d->1	
isan 	i->2	o->1	ä->1	
isan.	M->1	
isand	e->2	
isans	 ->1	
isar 	a->10	d->5	e->3	f->3	h->2	i->3	j->2	k->1	m->1	n->1	o->4	p->6	r->1	s->5	t->8	u->1	v->7	ä->3	
isar,	 ->2	
isar.	D->1	
isare	 ->2	
isas 	a->1	b->1	d->1	i->2	t->3	v->1	
isas,	 ->1	
isat 	a->9	d->2	e->4	h->1	i->1	m->1	o->1	p->4	s->8	v->1	
isat,	 ->1	
isat.	D->1	N->1	
isati	o->43	
isato	r->1	
isats	 ->3	
isavi	 ->1	
isbar	t->1	
isbes	t->9	
isbet	ä->1	
isbör	d->7	
iscay	a->6	
iscen	s->1	
isch!	 ->1	
ischl	e->4	
iscip	l->14	
isdag	 ->2	
isdik	t->5	
isdom	 ->1	
ise G	r->1	
iseen	d->1	
isekt	i->2	o->6	
isemi	t->3	
isen 	-->1	M->1	h->1	i->1	m->1	o->1	p->1	s->1	u->1	ä->2	
isen.	D->1	E->1	O->1	V->1	
isenb	e->3	
isens	 ->1	
iser 	f->1	i->1	o->3	u->1	
iser,	 ->1	
iser.	D->2	K->1	
isera	 ->39	.->1	d->26	n->2	r->12	s->12	t->10	
iseri	n->89	
isern	a->4	
ises 	i->1	p->1	
iset 	f->5	h->1	i->1	k->2	o->1	p->2	u->1	
iset.	D->1	F->1	
isfis	k->3	
isför	d->1	
ish P	e->1	
ishet	 ->1	,->1	.->1	
ision	 ->2	,->1	.->1	e->3	s->20	
isisk	,->1	a->65	e->2	t->2	
isiti	o->1	
isiär	a->1	
isk -	 ->1	
isk a	 ->1	g->1	l->7	n->4	r->3	s->1	t->2	
isk b	a->3	e->7	i->4	l->1	o->1	r->1	y->2	ö->1	
isk c	i->2	
isk d	e->7	i->7	
isk e	k->1	r->1	
isk f	e->1	i->2	l->2	o->2	r->4	y->1	ö->6	
isk g	e->4	l->1	r->3	
isk h	a->5	j->2	ä->1	
isk i	 ->1	d->1	m->1	n->10	
isk j	o->1	u->2	ä->2	
isk k	a->6	o->23	u->3	
isk l	a->4	e->5	i->5	ö->1	
isk m	a->6	e->3	i->3	o->1	y->2	
isk n	a->2	i->14	j->1	ä->1	
isk o	c->21	f->3	j->1	m->1	p->1	
isk p	a->1	e->2	l->2	o->16	r->4	u->1	
isk r	a->2	e->9	i->1	o->5	å->1	ö->1	
isk s	i->5	k->1	m->1	o->5	t->11	y->6	
isk t	i->6	r->2	y->1	
isk u	n->7	p->3	r->1	t->12	
isk v	e->1	i->1	ä->2	
isk ä	n->1	
isk å	k->13	
isk ö	v->3	
isk, 	e->2	f->1	k->1	m->2	s->1	
isk-i	s->1	
isk-s	k->1	
isk. 	J->1	
isk.D	e->1	
isk.H	e->2	
isk.I	 ->2	n->1	
isk.J	a->1	
isk.M	e->1	
isk.O	m->1	
isk.V	i->1	
iska 	E->2	F->1	K->1	P->1	T->1	a->31	b->50	c->3	d->19	e->17	f->85	g->43	h->19	i->81	j->3	k->130	l->31	m->69	n->11	o->124	p->71	r->91	s->110	t->22	u->271	v->29	ä->2	å->18	ö->5	
iska,	 ->12	
iska.	E->1	F->1	H->1	J->1	V->1	
iska:	 ->1	
iskab	e->1	
iskad	e->2	
iskan	 ->2	,->1	a->2	s->1	
iskar	e->2	n->1	t->1	
iskas	 ->1	
iskbe	d->4	s->4	
iske 	i->1	k->1	o->3	p->3	s->1	u->4	
iske)	 ->2	
iske,	 ->4	
iske.	-->1	D->1	
iskek	v->1	
iskem	ö->4	
isken	 ->16	,->1	
iskeo	m->2	
isker	 ->14	,->1	.->2	a->16	e->1	i->5	n->6	ä->1	
iskes	e->1	
isket	 ->3	,->1	r->3	s->1	
iskev	a->2	
iskfa	k->1	
iskfr	i->1	
iskfy	l->1	
iskfö	r->1	
iskha	n->6	
iskka	p->1	
iskko	m->2	
iskni	v->1	
iskof	ö->2	
iskoh	a->3	
iskol	i->3	
iskor	 ->40	,->3	.->1	n->24	s->14	
iskos	l->1	
iskre	t->1	
iskri	m->20	
iskt 	E->3	K->1	M->1	a->12	b->19	c->1	d->3	e->7	f->23	g->6	h->8	i->14	j->1	k->11	l->3	m->12	n->3	o->21	p->9	r->4	s->40	t->10	u->11	v->14	ä->5	å->1	ö->1	
iskt!	N->1	
iskt,	 ->7	
iskt.	A->1	B->1	D->4	G->1	J->1	S->1	Å->1	
iskup	p->1	
iskus	s->61	
iskut	a->3	e->78	
iskvo	t->2	
iskvä	r->3	
isläp	p->2	
ism -	 ->1	
ism e	l->2	t->1	
ism h	ä->1	
ism i	n->1	
ism m	å->1	
ism o	c->12	m->6	
ism p	å->1	
ism s	a->1	o->4	
ism u	n->1	
ism ä	n->1	r->1	
ism ö	v->1	
ism, 	a->1	f->1	i->1	m->1	n->2	o->2	s->1	v->1	ä->1	
ism.D	e->6	ä->1	
ism.F	r->1	
ism.H	e->1	
ism.I	 ->2	
ism.J	a->1	
ism.M	e->1	
ism.N	ä->1	
ism.O	c->2	
ism.V	a->1	i->3	
ism?V	i->1	
ismed	v->2	
ismen	 ->12	,->3	.->1	;->1	?->1	s->4	
ismer	 ->4	.->2	n->3	
ismis	k->2	
ismyn	d->2	
isnin	g->14	
isniv	å->1	
isnål	a->1	
isole	r->7	
isomr	å->1	
isont	a->2	e->1	
isor.	F->1	J->1	
isori	s->2	
isorn	a->1	
ispen	s->1	
ispli	t->1	
ispos	i->3	
israe	l->20	
iss b	a->1	r->1	
iss f	l->1	o->1	ö->3	
iss h	e->1	
iss i	 ->1	n->1	
iss m	a->1	e->1	i->1	ä->1	å->4	
iss o	e->1	m->1	r->2	s->1	
iss p	o->1	r->1	å->1	
iss r	e->1	
iss s	a->1	l->1	o->1	
iss t	i->2	v->1	y->2	
iss u	t->2	
iss v	i->1	å->1	
iss å	t->3	
iss ö	m->1	
iss, 	e->1	i->1	o->1	s->2	
iss.D	ä->1	
iss.E	n->1	
issa 	-->1	P->1	a->28	b->8	d->4	f->12	g->3	h->5	i->4	k->7	l->6	m->10	o->8	p->5	r->10	s->12	t->3	u->3	v->1	ä->8	å->1	ö->1	
issa.	M->1	
issab	o->8	
issad	 ->1	e->1	
issam	a->1	
issar	b->1	
issat	 ->1	
issbr	u->10	
issen	.->1	
isser	a->3	l->13	n->1	
issfa	l->1	
issfo	r->1	s->1	
issfö	r->4	
issgy	n->7	
isshe	t->4	
isshu	s->1	
issio	n->1151	
issit	u->1	
isskö	t->6	
issla	n->1	
issly	c->18	
isslö	s->1	
issnö	j->3	
isso 	e->1	i->1	o->1	ä->2	
isso,	 ->1	
issre	s->2	
isst 	b->1	d->1	f->1	j->1	k->2	n->1	
issta	 ->1	g->8	n->4	r->2	
isste	 ->4	x->1	
issto	l->1	
isstr	o->3	
issty	r->2	
isstä	n->4	
issup	p->2	
issys	 ->1	
issän	k->1	
ist E	u->3	
ist P	e->1	
ist a	n->1	t->3	v->2	
ist b	e->1	
ist f	a->1	r->1	ö->5	
ist k	o->1	r->1	
ist m	e->2	
ist n	ä->1	
ist o	c->3	
ist p	å->19	
ist s	a->1	o->1	t->1	v->1	
ist u	p->1	
ist v	i->2	
ist ä	r->2	
ist!T	v->1	
ist, 	k->1	m->2	o->2	
ist.G	i->1	
ista 	a->1	d->4	f->6	g->2	h->1	i->3	m->1	o->3	p->10	r->1	s->6	t->3	ä->6	ö->3	
ista,	 ->1	
ista.	.->1	D->1	E->1	S->1	V->2	
ista?	N->1	
istaN	ä->1	
istal	l->2	
istan	 ->48	,->4	.->13	d->12	s->3	
istas	 ->3	
istat	s->1	t->1	
istde	m->11	
iste 	o->1	p->1	u->1	
istef	r->1	
istel	s->1	
isten	 ->10	,->2	.->3	s->6	t->1	
ister	 ->54	!->1	,->6	.->13	a->19	m->2	n->45	p->3	r->14	
istfl	i->1	
istfä	l->8	
istgr	u->3	
istha	n->1	
istig	 ->1	t->2	
istik	 ->3	e->3	
istin	d->1	k->1	
istis	k->81	
istko	m->1	
istli	g->1	
istnä	m->2	
istor	i->36	
istpa	r->5	
istra	r->16	t->24	
istre	r->11	
istri	b->1	k->1	
ists 	p->1	
istse	k->2	
istyr	n->4	
istäl	l->2	
istå 	d->1	
iståe	n->1	
istån	d->22	
iståt	t->1	
isual	i->1	
isuel	l->1	
isum 	o->1	
isutv	e->1	
isväs	e->1	
isyst	e->1	
isäke	r->7	
isär 	d->2	s->1	
isäre	n->1	
it - 	j->1	m->1	
it FP	Ö->1	
it ak	t->2	
it al	l->3	
it an	f->1	g->1	
it ar	r->1	
it at	t->6	
it av	 ->2	
it be	t->1	v->1	
it bi	l->2	
it bo	r->2	
it bä	t->1	
it bå	d->1	
it de	 ->2	l->3	n->1	t->3	
it di	r->1	
it dä	r->3	
it ef	f->1	t->2	
it el	l->1	
it en	 ->21	g->1	
it er	t->1	
it et	a->1	t->11	
it fa	l->1	s->1	
it fe	l->2	
it fi	c->1	
it fl	e->1	
it fr	a->10	å->5	
it fö	r->8	
it ga	n->1	
it go	d->1	
it ha	l->1	r->1	
it hu	r->1	
it hä	n->7	r->1	
it hö	g->2	r->5	
it i 	a->1	d->2	e->1	f->2	g->1	v->1	
it ig	e->1	
it in	b->3	f->1	i->1	n->1	t->1	
it ko	m->1	n->1	r->1	
it kä	n->2	
it la	g->1	
it le	d->3	
it li	t->1	
it lo	v->1	
it lä	r->1	
it lå	n->1	
it me	d->7	r->1	
it mi	g->1	n->2	
it mo	t->2	
it my	c->4	
it mä	n->1	
it mö	j->3	
it ni	o->1	
it ny	t->1	
it nä	r->1	
it nå	g->4	
it nö	d->1	
it oc	h->4	
it oe	n->1	
it of	f->2	
it om	 ->1	k->1	
it pe	r->1	
it pl	a->1	
it po	s->1	
it pr	i->1	
it på	 ->6	,->1	s->1	
it ri	m->1	n->1	
it ru	l->1	
it se	n->1	
it si	g->10	n->1	t->1	
it sj	u->2	
it sk	u->1	
it sn	ö->1	
it so	m->1	
it sp	e->1	
it st	a->2	r->1	y->1	ä->3	ö->1	
it sv	å->1	
it sy	n->1	
it sä	r->1	
it så	 ->4	d->1	
it ta	g->1	
it ti	d->2	l->16	
it to	n->1	
it ty	c->1	d->1	
it un	d->6	
it up	p->15	
it ut	 ->1	l->1	s->1	t->1	
it va	d->1	n->1	r->2	
it vi	d->1	k->1	s->2	
it än	d->1	
it åt	g->1	
it öv	e->7	
it, b	ö->1	
it, e	n->1	t->1	
it, f	a->1	
it, m	e->1	
it, o	c->1	
it, v	i->1	
it, ä	v->1	
it-an	a->5	
it.Fr	u->2	
it.Fö	l->1	r->2	
it.I 	v->1	
it.Me	d->1	
it.Mo	t->1	
it.Nä	r->1	
it.Pa	r->1	
ita h	o->1	
ita i	 ->2	g->1	
ita o	c->2	s->1	
ita p	å->2	
ita s	i->1	
ita u	t->1	
ita v	a->1	
ita ä	r->1	
ita, 	u->1	
ita.D	ä->1	
ita.M	e->1	
ita.S	i->1	
itade	 ->1	
ital 	o->2	p->1	t->2	
ital,	 ->1	
ital.	S->1	
itale	t->5	
itali	e->18	s->2	
itals	k->3	
itame	n->8	
itan,	 ->1	
itann	i->14	
itano	 ->1	
itans	k->1	
itar 	o->1	p->5	s->2	v->1	
itari	s->4	
itas,	 ->1	
itat.	D->1	P->1	
itati	o->2	v->10	
itaue	n->1	
itbok	 ->12	,->1	.->5	e->35	
ite b	e->1	
ite e	x->1	
ite i	 ->1	
ite m	e->1	
ite s	k->1	
itel 	2->1	4->1	i->3	o->1	
iteln	 ->1	
iten 	-->2	b->1	d->2	e->1	f->1	g->1	k->1	m->4	n->1	o->1	p->2	t->1	u->1	ö->1	
iten.	D->1	J->1	
iter 	s->1	t->1	
iter,	 ->1	
iter-	b->1	
iter.	V->1	
itera	 ->5	.->2	d->4	r->10	s->5	t->1	
iteri	e->21	n->16	
iters	-->1	
itet 	-->2	a->10	b->3	d->1	e->3	f->6	g->4	h->4	i->18	k->3	l->3	m->11	o->32	p->3	s->12	t->4	v->2	ä->4	
itet!	H->1	
itet,	 ->35	
itet.	D->9	E->3	F->4	H->3	J->4	K->1	M->1	N->1	S->1	V->2	Ä->1	
itet:	 ->2	
itet?	H->2	N->1	
itete	n->55	r->20	
itets	-->1	a->2	b->3	f->2	g->1	h->2	k->3	n->1	o->1	p->19	r->3	s->2	
ithör	a->1	
itiat	i->80	
itica	l->1	
itie-	 ->1	
itied	e->2	
itiem	i->3	
itier	a->2	
itik 	-->2	J->1	a->5	e->2	f->19	h->4	i->7	k->3	m->11	n->1	o->25	p->1	r->2	s->26	t->1	u->2	v->3	ä->4	ö->1	
itik!	O->1	
itik"	 ->1	
itik,	 ->29	
itik.	.->1	D->8	E->2	F->2	H->3	I->1	J->1	M->1	R->2	T->1	V->2	Ä->1	
itik?	H->1	V->1	
itike	n->127	r->13	
itiko	m->6	
itiks	 ->1	
itima	 ->5	,->1	.->1	
itime	r->5	
itimi	t->6	
itimt	 ->2	,->1	
itin 	f->1	
itin.	A->1	
itio 	s->1	
ition	 ->20	,->4	.->2	;->1	a->2	e->42	s->8	
itise	r->10	
itish	 ->1	
itisk	 ->54	.->1	a->147	t->45	
itism	,->2	
itiv 	a->2	d->1	i->1	k->1	l->2	o->2	r->1	s->3	t->4	u->2	v->1	
itiv,	 ->1	
itiva	 ->26	
itivl	i->2	
itivt	 ->31	,->3	.->2	
itiös	 ->2	,->1	a->8	t->1	
itlan	d->2	
itlek	t->1	
itler	 ->3	,->1	-->1	s->1	
itlig	 ->3	h->2	
itlän	d->1	
itnin	g->1	
itori	e->9	n->8	u->8	
itrak	o->5	
itrea	 ->1	
itrov	i->1	
itrus	t->1	
itrut	t->1	
its a	n->1	v->7	
its b	e->1	
its d	e->1	
its e	t->1	
its f	r->3	ö->1	
its g	r->1	
its h	ä->1	
its i	 ->7	n->3	
its m	e->4	
its n	e->1	å->2	
its o	c->2	m->1	
its p	å->4	
its s	e->1	o->1	
its t	i->2	
its u	p->7	
its ä	n->1	r->1	
its, 	e->1	i->1	n->1	u->1	
its.B	e->1	
its.D	e->1	ä->1	
its.M	i->1	
its.S	o->1	
itt 2	3->1	
itt a	g->1	n->13	r->11	
itt b	e->10	i->2	
itt d	e->2	j->1	
itt e	g->12	r->2	
itt f	o->3	u->3	ö->10	
itt g	a->1	r->1	
itt h	e->4	u->1	
itt i	 ->5	b->1	n->2	
itt j	o->1	
itt k	a->1	o->2	
itt l	a->13	e->2	i->4	
itt m	a->1	e->6	o->2	
itt o	l->1	
itt p	a->6	e->1	r->1	å->2	
itt r	e->5	
itt s	a->2	e->1	l->1	o->1	p->1	t->8	v->1	y->1	
itt t	a->7	e->1	i->1	y->1	
itt u	n->1	p->2	t->3	
itt v	i->2	
itt y	t->5	
itt ä	m->2	n->2	
itt ö	d->1	p->1	
itt, 	f->2	r->1	
itt.M	i->1	
itta 	d->3	e->6	n->2	o->2	p->12	s->1	
ittad	e->1	
ittan	d->2	
ittar	 ->9	
ittat	 ->2	
itten	 ->3	.->1	
itter	 ->12	a->9	r->2	
ittet	 ->1	,->2	
ittil	l->44	
ittin	,->1	
ittis	k->16	
ittli	g->1	
ittna	 ->1	r->2	
ittne	 ->2	
ittni	n->2	
ittra	 ->1	d->1	f->1	s->1	
ittri	n->2	
ittsb	e->1	
ittsr	e->1	
itté 	-->2	e->1	f->3	h->1	m->1	s->2	
ittée	r->4	
ittéf	ö->2	
ittén	 ->23	,->4	.->2	?->1	s->11	
ittés	y->2	
itu m	e->20	
ituat	i->129	
itud 	7->1	
ituer	a->1	
itule	r->2	
itum.	D->1	
ituti	o->158	
ityd 	g->1	i->1	s->1	t->1	
ityd.	S->1	
itz i	 ->1	
itz. 	E->1	
itär 	o->1	v->1	
itära	 ->3	
itäre	r->1	
itärt	 ->1	
ium a	v->2	
ium b	l->1	
ium e	g->1	
ium i	n->2	
ium m	e->1	
ium o	c->3	
ium s	k->1	o->2	
ium!D	e->1	
ium, 	k->2	o->1	p->1	
ium.A	t->1	v->1	
ium.D	e->1	
ium.H	e->1	
ium.L	å->1	
ium.P	r->1	
ium.R	å->1	
ium.S	o->1	
ium.Ä	n->1	
iutsk	o->1	
iv (K	O->1	
iv - 	o->1	p->1	s->1	
iv 93	/->1	
iv 94	/->2	
iv 96	/->5	
iv En	l->1	
iv an	d->2	v->1	
iv at	t->2	
iv av	 ->1	v->1	
iv ba	s->1	
iv be	h->1	
iv bl	a->1	
iv de	 ->1	m->1	
iv di	s->2	
iv ef	t->1	
iv ek	o->2	
iv en	e->4	
iv fa	t->1	
iv fr	å->5	
iv få	r->2	
iv fö	r->10	
iv ge	n->1	
iv ha	 ->1	n->1	r->5	
iv hj	ä->1	
iv i 	d->3	s->2	v->1	
iv im	p->1	
iv in	o->1	r->2	t->3	v->1	
iv ka	n->1	r->1	t->1	
iv ko	m->2	n->5	s->1	
iv kv	a->1	
iv la	g->2	
iv le	d->1	
iv li	s->3	
iv lä	m->1	
iv lö	s->1	
iv me	d->1	n->1	
iv mi	l->1	n->1	
iv mo	t->1	
iv må	s->1	
iv oa	v->1	
iv oc	h->9	
iv om	 ->20	e->1	
iv op	i->1	
iv po	l->1	
iv på	 ->5	v->2	
iv re	f->1	
iv ri	k->1	
iv ro	l->2	
iv sa	k->1	
iv se	d->1	g->1	
iv si	d->1	
iv sk	a->1	u->1	
iv sn	a->1	
iv so	l->1	m->25	
iv st	a->5	i->1	r->2	å->1	
iv sy	f->1	s->2	
iv så	 ->2	d->1	s->1	
iv ta	l->1	
iv ti	l->15	
iv tr	ä->1	
iv ut	f->1	v->2	
iv ve	t->1	
iv vi	 ->1	d->1	l->2	
iv vä	n->1	
iv än	 ->1	
iv är	 ->5	
iv åt	g->2	
iv öv	e->1	
iv, 9	5->1	
iv, a	n->1	
iv, b	a->1	
iv, d	e->2	v->1	
iv, e	n->1	
iv, h	a->1	
iv, i	n->1	
iv, j	a->1	
iv, l	i->1	
iv, m	e->1	i->1	
iv, n	ä->1	
iv, o	c->4	m->1	
iv, s	o->2	t->1	ä->1	å->2	
iv, t	i->1	
iv, u	n->1	
iv. V	i->1	
iv.. 	(->1	
iv..H	e->1	
iv.At	t->1	
iv.Av	 ->1	
iv.Bl	a->1	
iv.De	 ->2	n->1	t->2	
iv.Då	 ->1	
iv.En	 ->1	
iv.Fö	r->4	
iv.I 	d->1	v->1	
iv.In	g->1	
iv.Lå	t->1	
iv.Me	n->2	
iv.Om	 ->1	
iv.Ri	k->1	
iv.Så	s->1	
iv.Vi	 ->1	s->1	
iv.Yt	t->1	
iv: F	ö->1	
iv: v	å->1	
iv; a	n->1	
iv?Fö	r->1	
iv?Ne	j->1	
iva a	n->2	r->1	v->2	
iva b	a->1	e->3	i->3	o->1	r->1	
iva c	e->1	
iva d	e->12	r->1	
iva e	f->4	n->8	t->1	x->1	
iva f	a->2	u->1	ö->6	
iva g	ä->1	
iva h	a->2	ö->1	
iva i	 ->2	d->1	g->1	n->3	
iva k	a->2	l->1	o->5	r->3	ä->1	
iva l	i->1	ö->1	
iva m	i->1	o->1	å->1	
iva n	i->1	å->1	
iva o	c->9	f->1	r->3	
iva p	a->1	o->4	r->2	u->1	å->2	
iva r	a->1	e->4	i->1	o->1	u->1	ä->1	
iva s	a->2	e->1	i->1	k->1	l->1	o->1	t->1	v->1	y->2	
iva t	e->1	i->9	r->1	
iva u	t->3	
iva v	e->2	ä->1	
iva å	s->1	t->3	
iva ö	v->1	
iva, 	f->1	s->1	u->1	ä->1	
iva.A	l->1	
iva.H	e->1	
iva.V	a->1	
ivade	s->1	
ivand	a->1	e->23	
ivare	 ->27	"->2	,->5	.->7	n->4	s->1	
ivark	o->1	
ivarl	ä->1	
ivarn	a->14	
ivarp	a->1	
ivas 	a->1	i->2	m->2	s->1	
ivas,	 ->1	
ivas.	I->1	M->1	
ivast	e->1	
ivat 	d->1	o->1	
ivat.	J->1	
ivata	 ->16	
ivate	k->1	
ivati	o->1	s->2	
ivats	 ->2	,->1	
ivavt	a->7	
ivbet	ä->1	
ivbor	d->1	
ive E	u->1	
ive a	l->1	n->1	
ive b	e->3	u->1	
ive d	e->4	
ive e	n->1	t->2	
ive f	o->1	
ive k	a->1	o->3	
ive l	a->2	
ive m	y->2	
ive p	a->3	
ive r	e->1	u->1	ä->1	
ive s	j->1	
ive t	i->1	r->1	
ivel 	a->7	g->3	l->1	n->1	o->6	p->1	t->2	u->1	v->1	ä->2	
ivel,	 ->2	
ivela	k->3	
ivels	e->5	u->3	
iven 	7->1	a->1	b->1	d->1	f->1	i->5	k->1	l->1	m->1	o->3	t->1	ö->1	
iven,	 ->2	
iven.	K->1	
ivenh	e->4	
ivens	 ->1	
iver 	O->1	a->3	e->5	f->1	h->1	k->1	m->1	n->2	r->1	s->1	t->2	u->2	v->1	
iver,	 ->1	
iver.	K->1	
ivera	 ->4	d->3	r->5	s->2	t->1	
iveri	 ->1	n->3	
ivers	a->1	e->5	i->2	
ives 	o->1	
ivet 	"->1	-->1	E->8	L->1	S->1	a->5	b->1	f->7	g->4	h->5	i->8	k->1	m->4	n->1	o->14	p->2	r->1	s->10	t->1	u->4	ä->8	
ivet"	 ->1	
ivet,	 ->13	
ivet.	 ->1	D->7	E->1	F->2	H->1	I->1	J->2	M->2	R->1	S->1	V->1	
ivets	 ->10	
ivetv	i->27	
ivför	m->1	s->3	
ivid 	h->1	s->1	
ivide	r->4	
ividu	a->1	e->7	
ivien	n->1	
ivier	 ->1	
ivil 	e->2	s->3	
ivil-	 ->1	
ivila	 ->3	
ivilb	e->2	
ivile	g->6	
ivilf	ö->2	
ivili	g->1	s->2	
ivill	i->12	
ivilr	ä->1	
ivils	k->2	
ivilt	 ->1	
ivise	r->3	
ivism	 ->1	
ivit 	a->2	b->2	d->1	e->8	f->1	g->1	h->1	i->1	l->3	m->1	o->1	s->7	t->2	u->6	v->1	
ivit.	F->1	
ivite	t->39	
ivits	 ->9	,->1	
ivkra	f->3	
ivla 	d->1	
ivla.	V->1	
ivlad	e->1	
ivlar	 ->5	
ivlat	 ->2	
ivlig	a->2	t->1	
ivlis	t->2	
ivna 	a->1	b->3	c->1	f->2	i->1	ä->1	
ivnin	g->11	
ivras	,->1	
ivrik	 ->1	
ivrät	t->4	
ivs a	v->2	
ivs e	f->1	n->1	
ivs g	e->1	
ivs i	 ->6	
ivs s	o->1	
ivs ö	v->1	
ivs, 	m->1	
ivs.D	e->1	
ivscy	k->3	
ivsdu	g->2	
ivskr	a->1	
ivskv	a->5	
ivsme	d->88	
ivsmi	l->3	
ivsup	p->1	
ivsvi	l->1	
ivt -	 ->1	
ivt a	n->1	r->3	t->7	
ivt b	e->3	l->1	
ivt d	e->2	
ivt e	l->1	
ivt f	r->1	u->1	ö->5	
ivt h	ö->1	
ivt i	 ->3	n->5	
ivt k	a->3	
ivt m	e->2	o->1	y->1	
ivt n	å->1	
ivt o	c->12	m->4	t->1	
ivt p	å->4	
ivt r	e->2	ä->2	
ivt s	a->2	e->2	k->1	n->1	o->1	p->1	t->4	v->2	ä->15	
ivt t	i->6	
ivt u	t->2	
ivt v	e->1	
ivt y	t->1	
ivt ä	r->1	
ivt å	l->2	
ivt ö	k->1	
ivt, 	d->2	i->1	m->1	o->1	p->1	r->1	
ivt. 	D->1	
ivt.D	e->2	
ivt.E	n->1	
ivt.I	n->1	
ivt.P	a->1	
ivt.Ä	v->1	
iväg 	o->1	s->1	
iväg,	 ->1	
ivå -	 ->1	
ivå a	v->3	
ivå d	ä->1	
ivå f	ö->5	
ivå g	e->2	
ivå h	a->1	
ivå i	 ->3	n->1	
ivå m	e->3	å->1	
ivå n	ä->1	
ivå o	c->5	f->1	m->1	
ivå p	å->2	
ivå s	o->8	å->1	
ivå u	p->1	t->2	
ivå v	i->1	
ivå ä	n->1	r->1	
ivå, 	a->1	b->2	d->1	f->2	g->1	m->1	o->2	r->2	v->1	
ivå.A	t->1	
ivå.B	i->1	
ivå.D	e->6	ä->1	
ivå.F	ö->1	
ivå.G	e->1	
ivå.H	e->2	
ivå.J	a->3	ä->1	
ivå.M	e->1	
ivå.N	ä->1	
ivå.P	å->1	
ivå.V	i->1	
ivå; 	d->1	
ivå?S	e->1	
ivåer	 ->6	,->2	.->4	:->1	n->1	
ivågr	u->3	
ivån 	-->1	f->1	i->2	m->1	p->3	
ivån.	D->3	H->1	
iwan 	i->1	
ix.De	 ->1	
ixas 	d->5	
ixen 	s->1	
ixtra	n->1	
iz el	l->1	
iz få	r->1	
iz fö	r->1	
iz so	m->1	
iz, G	i->1	
iz, t	a->1	
iz-ka	t->1	
izist	a->5	
iäker	h->1	
iär, 	i->1	
iära 	o->1	
iärer	 ->2	,->1	n->1	
iärmi	n->10	
iärpl	a->1	
iålde	r->1	
iåter	v->1	
ière 	k->1	
ié ut	a->1	
iös d	a->1	
iös o	c->1	
iös s	k->1	
iös u	t->1	
iös, 	k->1	
iösa 	a->1	m->3	o->1	p->2	s->2	
iösa,	 ->1	
iösa.	A->1	
iösar	e->2	
iöst 	a->2	l->1	o->1	s->2	
j 199	6->1	9->2	
j 200	2->1	
j Lib	e->1	
j ang	i->1	
j att	 ->1	
j avg	ö->1	
j ber	o->1	
j bes	v->1	
j bor	t->1	
j för	 ->2	r->1	
j i f	r->1	
j kom	m->1	
j lån	g->1	
j lös	t->1	
j mot	 ->1	
j när	 ->1	
j om 	n->1	
j til	l->1	
j är 	u->1	
j öve	r->1	
j, be	k->1	
j, bi	l->1	
j, de	t->1	
j, he	r->1	
j, ja	g->1	
j, ma	n->1	r->1	
j, na	t->1	
j, oc	h->1	
j, om	 ->1	
j, sk	a->1	
j, sä	g->1	
j, äv	e->1	
j-van	 ->1	
j.(Ap	p->1	
j.De 	t->1	
j.Exp	e->1	
j.I s	y->1	
j.Jag	 ->1	
j.Råd	e->1	
j.Ton	g->1	
j.Vi 	h->1	
ja - 	d->1	f->1	s->1	
ja Da	l->1	
ja FN	:->1	
ja Ha	i->1	n->1	
ja Jö	r->1	
ja Ma	l->1	
ja al	l->4	
ja an	s->9	v->4	
ja ar	b->3	t->1	
ja at	t->10	
ja av	 ->1	
ja be	 ->6	l->1	t->5	
ja bo	 ->1	
ja bö	r->5	
ja ch	a->1	
ja ci	t->1	
ja de	 ->14	m->2	n->13	s->6	t->12	
ja di	a->1	
ja ef	t->2	
ja ek	o->1	
ja el	l->2	
ja en	 ->15	
ja er	a->1	i->1	t->1	
ja et	t->4	
ja fo	r->2	
ja fr	a->7	å->6	
ja fu	n->2	
ja fä	s->1	
ja fö	r->21	
ja ge	 ->1	m->1	n->2	
ja gr	a->4	ä->1	
ja gö	r->10	
ja ha	 ->7	r->1	
ja hu	r->1	
ja hä	n->2	
ja hå	l->1	
ja hö	r->2	
ja i 	e->2	f->1	s->1	
ja in	i->1	v->1	
ja kl	.->1	
ja kn	y->1	
ja ko	m->3	n->2	
ja kr	i->2	
ja ku	l->2	
ja kv	i->3	
ja kö	p->1	
ja le	v->1	
ja li	k->2	
ja lo	k->1	
ja ly	f->1	
ja lä	g->2	
ja me	d->36	
ja mi	g->2	n->1	t->1	
ja my	c->1	
ja ny	a->1	
ja nä	m->2	s->1	
ja oc	h->7	
ja ol	i->1	
ja om	 ->1	
ja os	s->8	
ja pa	r->1	
ja pe	n->1	
ja pr	o->1	
ja på	 ->3	m->3	p->3	s->1	
ja re	g->1	s->2	
ja ri	k->1	
ja rä	d->1	k->2	
ja sa	m->3	
ja se	 ->2	
ja si	g->5	n->3	t->1	
ja sk	ä->1	
ja sl	å->1	
ja so	m->2	
ja st	r->4	ö->1	
ja sv	a->1	
ja sy	s->3	
ja sä	g->19	k->1	
ja t.	o->1	
ja ta	 ->9	c->9	
ja ti	l->14	
ja tv	å->1	
ja tä	n->1	
ja un	d->5	
ja up	p->11	
ja ur	s->1	
ja ut	 ->1	t->3	v->2	
ja va	r->4	
ja ve	t->4	
ja vi	s->1	
ja vå	r->2	
ja yr	k->1	
ja yt	t->1	
ja Ös	t->1	
ja åt	e->3	g->3	
ja öv	e->1	
ja, d	e->2	
ja, f	ö->1	
ja, g	a->1	
ja, h	e->1	
ja, l	e->1	
ja, m	e->1	
ja, p	r->1	
ja, t	i->1	ö->1	
ja, v	i->1	
ja...	L->1	
ja.He	r->1	
ja.Ja	g->2	
ja.Ko	m->1	
ja.Mi	n->1	
ja.Tr	o->1	
ja.Vi	 ->1	
jade 	a->2	d->2	e->1	f->2	g->1	h->1	i->3	m->1	u->1	Ö->1	
jades	 ->3	
jag -	 ->5	
jag 1	9->1	
jag G	a->1	
jag a	b->1	c->1	l->2	n->29	t->72	v->6	
jag b	a->8	e->26	l->2	
jag c	i->2	
jag d	e->7	o->3	ä->3	å->1	
jag e	m->5	n->6	r->12	t->1	
jag f	a->1	i->3	o->3	r->17	u->2	å->8	ö->41	
jag g	a->2	e->3	i->1	j->2	l->3	r->5	ä->7	ö->2	
jag h	a->38	e->7	o->16	ä->7	å->5	ö->5	
jag i	 ->16	n->57	
jag j	u->1	
jag k	a->22	l->2	o->25	r->1	u->2	ä->4	ö->1	
jag l	a->1	e->2	i->2	y->6	ä->3	å->1	
jag m	a->1	e->19	i->17	y->4	å->5	
jag n	a->5	i->1	o->2	u->5	y->2	ä->7	ö->1	
jag o	c->23	f->1	m->3	r->2	
jag p	e->4	o->4	r->1	å->9	
jag r	e->15	i->2	ä->1	å->1	ö->4	
jag s	a->8	e->9	j->14	k->39	o->1	p->1	t->7	v->2	y->2	ä->34	å->2	
jag t	a->28	i->8	r->41	v->3	y->17	ä->5	
jag u	n->4	p->16	t->10	
jag v	a->6	e->12	i->90	ä->7	å->1	
jag ä	l->1	n->3	r->34	v->2	
jag å	 ->2	t->2	
jag ö	n->1	
jag, 	a->1	e->2	f->2	g->1	h->1	i->1	m->1	o->1	s->1	u->1	ä->3	
jag. 	D->1	
jag.S	k->1	
jagar	 ->1	,->1	
jakt 	e->1	p->3	
jakti	g->6	
jaktl	i->14	
jala 	k->2	
jalis	t->4	
jalit	e->1	
jamo,	 ->1	
jan a	t->4	v->7	
jan d	e->1	
jan e	n->1	t->1	
jan f	i->1	r->4	
jan g	e->1	
jan h	a->1	ä->1	
jan i	 ->3	
jan o	c->1	m->1	
jan p	å->2	
jan t	i->1	
jan u	t->2	
jan, 	m->1	o->1	p->1	
janal	y->1	
jande	 ->51	.->2	:->8	n->3	t->13	
janua	r->16	
japan	s->1	
jar a	l->1	n->2	
jar b	l->2	y->1	
jar d	e->2	i->1	ä->1	
jar e	n->3	u->1	
jar f	i->1	
jar g	e->1	
jar k	u->1	
jar m	a->1	e->2	i->1	
jar n	u->1	
jar o	c->3	m->1	
jar p	a->1	r->1	å->1	
jar r	ö->2	
jar s	e->1	i->1	å->1	
jar t	i->2	r->1	
jar u	n->1	
jar å	 ->1	
jar.D	e->1	
jar.M	a->1	
jarba	s->1	
jard 	e->1	
jarde	r->14	
jare 	f->1	i->1	k->1	s->1	
jare.	 ->1	I->1	
jaren	 ->1	.->1	
jarna	 ->5	s->1	
jas a	v->8	
jas f	r->2	u->2	ö->4	
jas g	e->1	
jas i	 ->1	n->1	
jas m	e->1	
jas o	c->2	
jas s	o->1	
jas u	n->1	
jas å	t->1	
jas, 	f->3	m->1	
jas.H	e->2	
jas.M	e->2	
jas.N	ä->1	
jas.V	i->1	
jat -	 ->1	
jat a	n->2	
jat f	ö->1	
jat h	ö->1	
jat j	u->1	
jat l	a->1	
jat m	ä->1	
jat o	s->1	
jat s	a->1	i->2	t->2	
jat t	i->1	
jat v	i->1	
jat.I	 ->1	
jat.J	a->1	
jata 	o->1	
jats 	d->1	f->1	
jats,	 ->2	
jd - 	u->1	
jd at	t->1	
jd av	 ->18	
jd ga	r->1	
jd me	d->1	
jd på	 ->1	
jd sä	k->1	
jd ut	b->1	
jd.Ja	g->1	
jda m	e->6	ö->1	
jda, 	d->1	f->1	o->1	
jdas 	g->1	
jdat 	f->1	
jde a	t->1	
jde b	e->1	
jde d	e->1	
jde p	å->1	
jde s	å->1	
jde u	p->1	
jden 	e->1	
jder 	b->1	d->2	f->7	
jdern	a->9	
jdes 	a->1	i->1	
jdosk	o->1	
jdpun	k->2	
jdrik	t->1	
jdska	d->2	
jdåtg	ä->1	
je (B	e->1	
je - 	h->1	
je 10	0->1	
je Ba	r->1	
je EU	-->1	
je Eu	r->1	
je an	a->1	s->1	
je as	p->1	
je at	t->1	
je av	t->1	
je be	h->2	r->1	
je bi	l->1	
je bo	k->1	
je da	g->7	
je de	l->2	m->1	
je di	s->1	
je en	s->5	
je eu	r->2	
je fa	l->6	
je fi	n->1	
je fo	l->2	r->4	
je fr	a->1	ä->1	
je fö	r->4	
je ga	r->1	
je ge	o->1	
je gr	u->1	
je gä	l->1	
je gå	n->4	
je ha	l->2	
je in	d->1	g->1	s->1	
je ko	m->2	
je ku	l->1	
je la	n->31	
je lä	n->2	
je me	d->14	
je mi	l->2	
je må	n->2	s->2	
je no	t->1	
je oa	v->1	
je oc	h->4	
je pe	l->1	
je pr	o->1	
je pu	n->4	
je re	g->2	
je ri	k->2	
je rä	t->1	
je sa	k->1	m->1	
je so	m->4	r->1	
je st	a->3	
je su	v->1	
je vi	l->2	
je vä	r->2	
je är	 ->1	
je år	 ->6	.->3	t->1	
je åt	g->1	
je öv	e->3	
je, a	n->1	t->2	
je, v	i->1	
je- o	c->1	
je.Ge	n->1	
je.Ja	g->1	
je: u	t->1	
jebef	r->1	
jebol	a->4	
jebäl	t->10	
jedel	 ->4	a->2	
jedom	a->1	
jefad	e->1	
jeför	f->1	o->1	
jeind	r->2	u->1	
jejor	d->3	
jekok	a->1	
jekon	c->1	
jekt 	f->7	h->1	i->1	l->1	m->2	o->2	p->1	s->11	v->2	ä->1	
jekt"	,->1	
jekt,	 ->6	
jekt.	D->1	S->1	
jekt?	T->1	U->1	
jekta	d->2	
jekte	n->9	t->14	
jekti	v->3	
jelan	d->6	
jelin	j->1	
jelse	 ->1	r->3	
jemäs	s->1	
jen b	ö->1	
jen h	a->1	
jen i	 ->1	
jen.D	ä->1	
jer 9	7->1	
jer a	t->2	
jer b	l->1	
jer d	e->4	
jer e	l->1	x->1	
jer f	ö->10	
jer g	ä->1	ö->1	
jer h	a->1	ö->1	
jer i	 ->5	n->2	
jer j	a->1	
jer k	a->1	o->1	
jer l	e->1	
jer m	a->1	e->3	i->1	å->1	
jer n	i->1	ä->2	
jer o	c->6	m->3	
jer p	r->1	å->1	
jer r	e->1	
jer s	i->10	o->8	
jer u	t->2	
jer v	i->4	
jer ä	r->1	
jer å	t->1	
jer".	D->1	
jer, 	d->1	e->1	i->1	m->2	p->1	r->1	s->2	u->1	
jer.D	e->1	
jer.H	e->1	
jer.M	e->1	
jer.V	i->1	
jer: 	a->1	
jerad	 ->4	e->7	
jerat	 ->3	,->2	
jerna	 ->28	,->3	.->2	s->2	
jeska	d->1	
jesta	r->1	
jet a	t->2	
jetan	k->9	
jetra	n->1	
jetru	s->1	
jetti	d->1	
jetto	n->1	
jeuts	l->2	
jeväc	k->3	
jeåte	r->1	
jflöd	e->1	
jikis	t->5	
jkan 	k->1	
jkont	r->2	
jkott	.->1	
jlig 	a->2	e->1	i->1	m->1	o->1	r->1	s->1	
jlig.	 ->1	J->1	
jliga	 ->30	.->1	
jlige	n->6	
jligg	j->3	ö->9	
jligh	e->131	
jligt	 ->88	!->1	,->8	.->22	
jning	 ->11	.->3	e->2	s->3	
jobb 	e->1	o->1	
jobb,	 ->2	
jock 	o->1	
jocka	 ->1	
jol o	c->2	
jol, 	o->1	
jol.K	ä->1	
jon i	n->1	
joner	 ->59	,->2	.->1	n->1	
jonis	e->1	
jonta	l->1	
jor o	c->1	
jor.F	r->1	
jord 	-->1	
jord.	E->1	V->1	
jorda	 ->2	,->1	
jordb	r->54	ä->10	
jorde	 ->31	,->1	.->1	n->3	s->5	
jordm	å->1	
jords	k->1	
jorit	e->42	
jorna	.->1	
jort 	a->2	b->1	d->10	e->13	g->1	h->2	i->1	k->2	m->2	n->4	o->4	p->1	r->1	s->8	u->3	v->2	å->1	
jort,	 ->8	
jort.	D->1	I->1	J->1	L->1	R->1	S->1	
jorto	n->9	
jorts	 ->18	,->3	.->2	
jos a	n->1	
journ	a->2	e->1	
jovis	 ->1	)->1	b->9	e->1	f->3	k->2	
js av	 ->1	
js ka	n->1	
js oc	h->1	
js ti	l->1	
js up	p->2	
js, f	ö->1	
js.(E	N->1	
jsmål	 ->1	.->1	
jt i 	E->1	
jt os	s->1	
jt si	g->1	
jt ut	 ->1	
jt vi	s->1	
jts t	i->2	
jts u	p->1	
jts, 	o->1	
ju Eg	y->1	
ju Mo	r->1	
ju ab	s->1	
ju al	l->5	
ju an	v->1	
ju at	t->3	
ju av	 ->1	
ju ba	r->2	
ju de	 ->1	t->1	
ju di	r->1	
ju dä	r->1	
ju då	 ->1	
ju em	e->1	
ju en	 ->1	
ju fö	g->1	r->1	
ju gå	n->1	
ju hä	r->1	
ju in	b->1	d->1	g->2	o->1	s->1	t->5	
ju is	o->1	
ju lä	n->1	
ju me	d->1	r->4	
ju mo	r->1	
ju må	s->1	
ju oc	k->7	
ju of	t->1	
ju pa	r->1	
ju po	r->1	
ju pu	n->1	
ju på	 ->1	
ju re	d->2	s->1	
ju sa	m->2	
ju si	n->1	
ju so	m->1	
ju st	ä->2	ö->1	
ju ti	l->1	
ju ut	t->1	
ju vi	l->1	
ju än	d->2	
ju är	 ->5	
ju, o	c->1	
ju, p	r->1	
ju, å	t->1	
juade	s->1	
jubla	n->1	
juda 	a->1	b->3	d->1	e->3	i->1	k->1	m->1	n->1	o->1	p->1	u->1	
judan	 ->1	d->4	
judar	s->1	
judas	,->1	.->1	
judda	 ->1	
juden	 ->1	
juder	 ->11	,->1	
judet	 ->3	.->1	
judeu	t->1	
judic	e->1	
judik	a->3	
judis	k->1	
judit	 ->1	
judli	g->1	
judna	 ->2	
judni	n->1	
juger	 ->1	
jugo 	g->1	å->1	
jugof	e->1	
jugon	d->1	
juk.J	a->1	
juka 	P->1	
juka,	 ->1	
jukdo	m->1	
jukfö	r->1	
jukhu	s->7	
jukni	n->2	
jukvå	r->3	
jul o	c->1	
julfe	r->1	
juli 	1->4	2->2	f->1	u->1	
juli,	 ->2	
julkl	a->1	
junde	 ->4	
junge	l->2	
jungf	r->1	
juni 	1->6	2->2	f->2	i->1	v->1	
junka	 ->3	.->1	
junke	r->2	
junki	t->2	
junkn	a->1	
junkt	u->1	
jup ö	n->1	
jupa 	f->1	m->1	o->1	s->1	u->1	
jupa,	 ->1	
jupad	 ->1	
jupar	e->1	
jupas	 ->1	t->2	
jupat	 ->2	
jupet	 ->3	,->2	
jupgå	e->7	
jupni	n->5	
jupsi	n->1	
jupt 	b->2	d->1	o->1	s->1	v->1	ö->1	
jur o	c->1	
jur ä	r->1	
jur, 	a->1	f->1	
jur- 	o->2	
jur.D	ä->1	
jur.H	e->1	
jurar	t->1	
juren	s->1	
juret	 ->1	
jurfo	d->4	
jurid	i->30	
juris	 ->4	.->1	d->5	t->7	
jurli	v->2	
jus p	å->1	
jus.I	n->1	
juset	 ->7	.->1	
just 	a->2	b->3	d->17	e->1	f->12	g->3	h->14	i->4	l->2	m->3	n->12	o->1	p->5	r->1	s->7	v->3	ö->1	
just,	 ->1	
just.	D->1	K->1	
just:	 ->1	
juste	r->6	
justi	c->4	t->6	
juta 	i->1	m->1	r->1	u->5	v->1	
jutan	d->1	
jutas	 ->3	
juten	 ->2	
juter	 ->6	
jutit	s->5	
jutni	n->1	
juts 	s->1	u->4	
jutto	n->2	
jutva	p->1	
juvel	e->2	
jäl d	e->1	
jäl, 	i->1	
jäl.F	r->1	ö->1	
jälen	"->1	.->1	
jälp 	a->27	d->1	f->6	n->1	o->2	p->1	s->2	t->5	v->2	ö->1	
jälp,	 ->2	
jälp.	D->1	H->1	I->1	J->1	V->1	
jälpa	 ->37	n->3	r->1	
jälpe	n->4	r->1	
jälpl	i->1	
jälps	.->1	
jälpt	 ->1	a->1	e->1	
jälpv	i->1	
jält 	a->1	e->1	p->1	
jälv 	a->5	b->2	f->5	g->1	h->3	i->3	k->1	m->1	o->3	s->7	t->1	u->2	v->2	ä->3	
jälv,	 ->5	
jälv.	D->1	J->1	K->1	V->1	
jälva	 ->61	,->3	.->5	
jälvb	e->3	i->1	ä->1	
jälvf	a->2	ö->1	
jälvh	j->1	
jälvk	l->20	o->1	
jälvp	l->1	
jälvs	t->15	ä->1	
jälvt	 ->5	
jälvä	n->1	
jämfö	r->16	
jämka	 ->1	r->1	
jämli	k->13	
jämn 	s->1	
jämn,	 ->1	
jämn.	D->1	
jämna	 ->4	d->1	
jämni	n->2	
jämnv	i->1	
jämsi	d->1	
jämst	ä->23	
jämt 	e->1	ö->1	
jämt.	D->1	
jämvi	k->2	
jäna 	a->1	n->1	s->2	
jänad	e->1	
jänar	 ->14	.->2	
jänst	 ->6	,->1	.->2	e->110	f->1	g->3	
jänt 	a->1	p->1	
jänta	 ->27	
jära.	N->1	
järde	 ->8	-->1	d->2	
järer	n->1	
järn-	 ->2	
järna	.->1	n->1	
järnv	ä->15	
järta	 ->3	d->1	n->2	t->14	
järtl	i->7	
järv 	o->1	
järva	 ->2	r->1	
järvh	e->1	
järvt	 ->2	
jätte	 ->19	,->1	d->1	
jävul	e->1	s->1	
jö fö	r->2	
jö i 	d->1	
jö ka	n->1	
jö mo	t->1	
jö sa	k->1	
jö so	m->1	
jö vi	n->1	
jö!De	t->1	
jö, f	o->7	
jö, h	ä->1	
jö, l	i->1	
jö, s	m->1	
jö, u	p->1	
jö- o	c->2	
jö.De	t->2	
jö.Då	 ->1	
jö.Me	n->1	
jö.Un	d->1	
jö.Vi	l->1	
jöanp	a->1	
jöans	v->2	
jöavt	a->1	
jöbel	a->1	
jöbes	k->1	t->1	
jöbro	t->1	
jöd f	ö->1	
jödep	a->1	
jödir	e->1	
jöds 	t->1	
jöer 	f->1	i->1	s->1	
jöern	a->1	
jöfak	t->1	
jöfar	l->1	t->8	
jöfrå	g->4	
jöför	b->1	h->1	s->2	
jöinf	o->1	
jökas	t->1	
jökat	a->10	
jökon	f->1	s->5	
jökra	v->8	
jökva	l->1	
jölag	s->1	
jömin	i->1	
jömän	 ->2	
jömäs	s->11	
jömål	 ->2	s->1	
jön e	l->1	n->1	
jön f	ö->1	
jön h	å->1	
jön i	 ->1	
jön o	c->6	
jön p	å->1	
jön s	o->1	
jön t	i->1	
jön ä	r->1	
jön!D	e->1	
jön, 	a->1	d->1	h->1	m->1	o->3	s->1	u->1	
jön.D	e->2	ä->1	
jön.E	n->1	
jön.F	r->1	
jön.J	a->1	
jön.L	å->1	
jön.M	a->1	
jön.U	n->1	
jön.V	i->1	å->1	
jönk 	h->1	r->1	u->1	
jönk.	D->1	
jönor	m->2	
jöns 	f->1	s->1	
jöomr	å->4	
jöovä	n->1	
jöper	s->1	
jöpol	i->8	
jöpro	b->3	g->1	
jöpåv	e->1	
jör -	 ->2	
jöråd	e->1	
jörör	e->2	
jösek	t->1	
jösid	a->1	
jöska	d->2	
jösky	d->11	
jöskä	l->2	
jöss 	o->1	p->1	ä->1	
jöss)	 ->1	
jöste	d->4	
jöstö	d->1	
jösyn	p->6	
jötra	n->1	
jöuts	k->1	
jövän	l->7	
jövär	d->3	
k - d	e->2	ä->1	
k - n	ä->1	
k - o	c->1	
k - v	i->1	
k Det	t->1	
k Jör	g->1	
k Kir	g->1	
k TV 	a->1	
k a p	r->1	
k agi	t->1	
k al-	S->1	
k all	d->1	m->7	
k ana	l->1	
k and	r->1	
k ang	e->2	
k ant	a->1	i->1	
k anv	ä->1	
k art	.->2	i->1	
k asp	e->1	
k att	 ->24	
k av 	D->1	a->5	d->3	k->2	s->1	v->1	
k bak	å->1	
k bal	a->2	
k bar	a->2	
k bas	a->1	t->1	
k bel	y->1	
k ber	o->1	ä->1	
k bes	i->1	k->1	l->1	t->1	
k bet	r->1	y->4	
k bil	i->4	
k bli	r->1	
k blo	c->1	
k boj	k->1	
k bor	d->1	
k bro	t->1	
k byg	g->1	
k byr	å->2	
k böj	e->1	
k civ	i->2	
k dag	 ->1	s->1	
k de 	g->1	
k deb	a->4	
k dem	o->2	
k den	n->1	
k det	 ->3	,->1	a->1	t->1	
k dia	l->2	
k dim	e->1	
k dis	k->4	
k eft	e->3	
k ege	n->1	
k ej 	b->1	
k eko	n->1	
k ell	e->4	
k eme	l->1	
k en 	f->1	g->1	m->1	s->1	ö->1	
k ene	r->1	
k eni	g->1	
k ers	ä->1	
k eta	p->1	
k ett	 ->1	
k fed	e->1	
k fie	n->1	
k fil	o->1	
k fin	n->2	
k fla	g->2	
k fon	d->1	
k for	c->1	s->1	
k fra	m->2	
k fru	 ->2	
k frä	m->1	
k frå	g->4	n->3	
k fys	i->1	
k få 	p->1	
k får	 ->2	
k för	 ->44	,->1	.->1	d->1	e->2	n->1	
k gav	 ->1	
k gem	e->1	
k gen	o->3	
k ges	t->1	
k gjo	r->1	
k glu	p->1	
k gra	n->1	
k gru	p->1	
k grö	n->2	
k gäl	l->3	
k går	 ->2	
k ham	n->1	
k han	d->4	
k har	 ->12	
k hel	t->1	
k hjä	l->2	
k hon	 ->1	o->1	
k hop	p->1	
k hur	 ->1	
k huv	u->1	
k hän	d->2	
k hör	 ->1	a->2	
k i A	f->1	k->1	
k i E	u->2	
k i K	i->1	
k i L	u->1	
k i T	a->1	u->1	
k i W	i->1	
k i a	l->1	
k i d	e->1	
k i e	t->1	
k i f	.->1	o->1	r->2	
k i g	e->1	
k i h	i->1	
k i k	a->2	
k i m	i->1	
k i n	å->1	
k i o	c->1	
k i r	e->1	
k i s	a->1	t->2	y->1	
k i u	p->1	
k i v	å->2	
k ide	n->1	
k imm	i->1	
k in 	b->1	
k ind	u->1	
k ing	e->1	
k inl	e->1	
k ino	m->2	
k inr	e->1	i->2	
k ins	p->1	t->4	
k int	e->14	r->1	
k jag	 ->4	
k jor	d->1	
k ju 	i->1	s->1	
k jur	i->1	
k jus	t->1	
k jäm	s->1	
k jät	t->1	
k kam	p->1	
k kan	 ->5	a->3	d->1	s->1	
k kar	t->1	
k kat	a->3	
k kla	r->1	
k klo	a->1	
k kom	m->6	
k kon	f->3	k->4	s->2	t->14	
k kos	t->1	
k kul	t->3	
k kun	n->1	
k kur	s->1	
k kvi	n->1	
k kän	n->1	s->1	
k lag	 ->1	,->1	.->1	s->2	
k led	a->2	
k leg	i->3	
k liv	s->5	
k lov	a->1	
k lyc	k->1	
k läg	g->1	
k läk	a->1	
k län	g->1	
k lös	n->1	
k mak	t->3	
k mar	k->2	
k mat	e->1	
k med	 ->11	b->1	v->1	
k mel	l->2	
k men	 ->1	
k mer	 ->1	
k mig	,->1	
k mil	i->1	j->1	
k min	o->1	
k mis	s->1	
k mod	e->2	
k mot	 ->5	
k myc	k->2	
k myn	d->3	
k mås	t->6	
k möj	l->2	
k nat	i->2	u->1	
k ned	 ->1	
k niv	å->14	
k nju	t->1	
k nu 	s->1	
k nya	 ->1	
k när	 ->5	
k någ	o->2	r->1	
k och	 ->72	
k ock	s->2	
k off	e->4	
k ojä	m->1	
k om 	T->1	e->1	f->1	k->1	l->2	m->3	r->1	
k oms	t->1	
k ope	r->1	
k ori	e->1	
k oss	 ->3	
k par	l->3	
k per	s->2	
k pla	n->2	
k pol	i->19	
k poä	n->1	
k pro	c->2	d->2	f->1	
k pun	k->1	
k på 	1->1	E->1	V->1	a->3	d->3	g->1	n->1	o->2	
k rak	t->1	
k ram	,->1	
k ras	i->1	
k rea	g->1	
k ref	o->3	
k reg	e->2	i->1	
k rek	o->1	
k ren	s->2	
k ret	r->1	
k ris	k->1	
k rol	l->5	
k rät	t->1	
k råd	g->1	
k rör	a->2	
k sad	e->2	
k sam	t->1	
k se 	s->1	
k seg	l->1	
k sen	a->1	
k sig	n->2	
k sit	u->3	
k sjä	l->1	
k ska	d->1	l->3	p->1	
k sku	l->1	
k sky	l->1	
k skö	t->1	
k smi	t->1	
k sna	b->1	
k sol	i->2	
k som	 ->58	
k sta	b->1	d->2	r->1	t->4	
k str	a->4	i->1	u->3	
k svå	r->1	
k syn	p->3	v->3	
k säg	a->1	
k säk	e->1	
k sär	s->1	
k så 	a->1	m->15	
k såd	a->1	
k ter	r->1	
k tig	e->1	
k til	l->29	
k tra	d->1	s->1	
k tro	t->1	
k tvi	v->1	
k tvu	n->1	
k typ	,->1	
k tän	k->1	
k und	e->3	
k uni	o->5	
k upp	f->3	g->1	l->1	s->1	
k urs	p->1	
k ut 	p->1	
k uta	n->1	
k utb	i->2	
k utg	ö->1	
k utm	a->2	
k utt	r->1	
k utv	e->7	i->1	ä->1	
k vad	 ->1	
k var	 ->2	e->7	i->1	
k ver	k->1	
k vi 	b->1	i->1	l->1	r->1	
k vid	 ->3	a->1	
k vik	t->1	
k vil	j->4	k->1	l->3	
k vin	d->1	
k vit	t->1	
k väg	 ->1	,->1	r->1	
k vär	t->1	
k än 	r->1	
k änn	u->1	
k är 	W->1	b->1	d->3	f->2	g->1	n->2	v->2	
k åkl	a->13	
k åte	r->1	
k åtm	i->2	
k öve	r->4	
k övn	i->1	
k!And	r->1	
k!Om 	v->1	
k" - 	e->1	
k" fö	r->1	
k" oc	h->1	
k, 15	 ->1	
k, Re	a->1	
k, at	t->1	
k, be	n->1	
k, de	c->1	n->2	s->3	t->3	
k, dv	s->2	
k, då	 ->2	
k, ef	t->2	
k, en	 ->2	
k, ex	e->1	
k, fi	n->1	
k, fr	a->1	u->4	å->1	
k, fö	r->3	
k, go	d->1	
k, gå	r->1	
k, ha	r->1	
k, he	r->6	
k, hä	r->1	
k, i 	b->1	h->1	
k, in	n->1	t->3	
k, ko	m->5	
k, kä	r->1	
k, me	n->8	
k, mo	d->1	
k, ne	d->1	
k, nä	r->2	
k, nå	g->1	
k, oc	h->2	k->1	
k, sa	m->2	
k, sk	a->1	
k, so	m->6	
k, så	 ->2	
k, ti	l->1	
k, tr	a->11	o->1	
k, ut	a->1	
k, va	r->2	
k, vi	l->2	
k, vä	g->1	
k, är	l->1	
k- el	l->1	
k- oc	h->2	
k-bri	t->1	
k-dam	m->1	
k-fra	n->1	
k-isr	a->1	
k-pos	i->1	
k-ska	n->1	
k. De	t->1	
k. Ja	g->1	
k. Me	n->1	
k. an	s->1	
k. in	t->1	
k. sk	o->1	
k. so	f->1	
k..(F	R->1	
k.Att	 ->2	
k.Avg	å->1	
k.Bet	ä->1	
k.Byg	g->1	
k.De 	f->1	h->1	u->1	
k.Den	n->1	
k.Det	 ->11	t->5	
k.Där	f->1	
k.Då 	k->1	o->1	
k.En 	a->1	
k.Ett	 ->1	
k.Eur	o->1	
k.Fak	t->1	
k.Fru	 ->1	
k.Frå	g->3	
k.För	s->1	
k.Gen	o->1	
k.Han	 ->2	
k.Her	r->7	
k.Hit	 ->1	
k.Hur	 ->1	
k.Här	 ->1	
k.I b	e->1	
k.I d	e->1	
k.I g	å->1	
k.Inf	ö->1	
k.Jag	 ->7	
k.Kin	n->1	
k.Kom	m->1	
k.Men	 ->3	
k.Ni 	h->1	
k.Och	 ->1	
k.Om 	m->1	
k.Ref	o->1	
k.Rik	t->1	
k.Syr	i->1	
k.Tac	k->1	
k.Trä	d->1	
k.Tvä	r->1	
k.Tyv	ä->1	
k.Van	 ->1	
k.Vi 	d->1	m->1	r->1	s->3	t->1	v->1	
k.Vil	k->1	
k.Äve	n->2	
k: ge	m->1	
k: vi	 ->1	
k?Her	r->1	
k?Nej	,->1	
k?Reg	e->1	
k?Vad	 ->1	
ka "s	h->1	
ka - 	b->1	d->1	f->1	o->1	
ka 17	0->1	
ka 25	0->1	
ka Ah	e->1	
ka Ba	r->1	
ka EU	-->1	
ka Eu	r->5	
ka FP	Ö->1	
ka Fl	é->1	
ka Gr	a->1	o->1	
ka Ka	r->1	
ka Ko	c->1	
ka Ku	n->1	
ka La	n->1	
ka PV	C->1	
ka Pa	l->2	
ka Po	e->2	
ka Sc	h->1	
ka TV	-->1	
ka ab	s->1	
ka ak	t->3	
ka al	d->1	l->14	
ka am	b->1	
ka an	a->1	d->3	k->1	l->1	m->1	s->3	t->3	v->6	
ka ar	b->11	g->3	m->2	r->1	v->1	
ka as	p->2	
ka at	l->1	o->2	t->34	
ka au	k->1	
ka av	 ->4	a->1	s->3	
ka ba	l->1	n->1	s->2	
ka be	d->4	f->7	g->4	h->5	k->2	m->1	r->1	s->17	t->8	v->1	
ka bi	d->2	l->14	
ka bl	.->1	i->1	
ka bo	r->1	
ka br	a->1	å->1	
ka bu	d->6	
ka by	g->3	r->1	
ka bå	t->1	
ka bö	r->2	
ka ce	n->3	
ka da	g->1	
ka de	 ->14	b->3	f->1	l->7	m->9	n->21	p->1	r->1	s->5	t->16	
ka di	k->1	m->2	r->1	s->2	
ka dj	u->2	
ka do	m->4	
ka du	m->1	
ka dy	r->2	
ka dä	r->1	
ka ef	f->4	t->2	
ka ek	o->8	v->1	
ka el	l->2	
ka em	e->1	
ka en	 ->11	a->2	h->1	
ka er	 ->6	,->1	f->1	s->1	
ka et	a->1	c->1	n->1	t->5	
ka eu	r->2	
ka ex	e->1	i->1	t->3	
ka fa	k->2	l->1	r->5	s->4	t->1	
ka fi	n->1	s->4	
ka fl	a->1	y->2	
ka fo	l->27	n->1	r->8	
ka fr	a->6	i->1	u->3	å->18	
ka fu	s->2	
ka fy	r->1	
ka få	 ->2	n->1	
ka fö	d->1	l->5	r->101	
ka ga	m->1	r->2	
ka ge	 ->1	m->15	n->8	o->1	
ka gi	c->1	l->1	v->1	
ka gr	u->31	y->1	ä->1	
ka gä	r->2	
ka ha	 ->1	l->1	m->3	n->5	r->1	v->3	
ka he	l->2	n->4	r->4	
ka hi	n->2	s->1	t->1	
ka hj	ä->1	
ka ho	n->2	
ka hu	n->1	r->2	v->1	
ka hä	l->1	n->4	
ka hå	l->3	r->3	
ka hö	g->2	
ka i 	G->1	a->2	d->6	f->2	l->1	m->1	p->2	s->3	t->1	u->2	
ka id	e->1	
ka ih	o->1	
ka im	m->1	
ka in	b->1	c->1	d->4	f->1	i->3	k->1	l->1	n->4	s->38	t->41	v->1	
ka is	o->1	
ka ja	g->1	
ka jo	r->2	
ka jä	m->2	r->1	
ka ka	l->1	m->2	n->4	r->5	t->4	
ka ki	n->1	
ka kl	a->1	o->1	y->1	
ka ko	l->6	m->77	n->50	s->1	
ka kr	a->7	e->2	i->11	å->1	
ka ku	l->6	n->1	s->11	
ka kv	i->2	o->1	ä->1	
ka ky	l->1	
ka kä	n->3	r->1	
ka la	g->4	n->1	
ka le	d->13	
ka li	b->8	g->1	k->1	t->2	v->4	
ka lo	b->1	k->2	
ka lä	g->2	m->1	n->14	
ka lö	n->1	s->1	
ka ma	j->1	n->1	r->6	s->3	
ka me	d->45	r->1	t->3	
ka mi	g->1	k->1	l->6	n->15	s->1	t->4	
ka mo	b->1	d->4	t->3	
ka my	c->4	n->15	
ka mä	n->1	
ka må	l->13	n->5	s->1	t->1	
ka mö	j->7	
ka na	t->11	
ka ne	d->1	
ka ni	 ->1	v->2	
ka no	r->2	
ka nu	n->1	
ka ny	a->2	
ka nä	m->1	r->3	s->1	t->2	
ka nå	g->2	
ka nö	d->2	
ka ob	a->1	
ka oc	h->68	
ka oe	g->1	
ka of	f->4	t->2	
ka oi	n->1	
ka ok	l->1	
ka ol	y->1	
ka om	 ->4	b->2	r->10	s->4	
ka on	ö->1	
ka op	e->1	p->1	
ka or	d->75	g->2	o->2	s->1	
ka os	s->1	
ka pa	r->22	
ka pe	n->4	r->3	
ka pl	a->8	
ka po	l->20	p->1	
ka pr	e->4	i->7	o->26	
ka pu	n->7	
ka på	 ->26	,->1	
ka ra	d->3	m->1	p->16	
ka re	a->2	f->1	g->54	n->3	p->3	s->7	v->2	
ka ri	k->6	s->5	
ka ru	t->1	
ka rä	t->8	
ka rå	d->22	
ka rö	s->4	
ka sa	k->2	m->12	n->1	
ka sc	e->2	
ka se	 ->1	d->1	g->1	k->3	
ka si	g->7	n->9	t->16	
ka sj	ä->1	ö->3	
ka sk	a->3	e->2	i->4	o->2	r->1	u->1	y->1	ä->7	
ka sl	a->2	u->3	
ka so	c->27	l->1	m->4	
ka sp	e->2	r->1	ä->1	
ka st	a->16	e->3	i->1	o->4	r->10	u->1	y->2	ä->1	å->3	ö->11	
ka sv	a->1	å->6	
ka sy	f->1	n->1	s->12	
ka sä	k->3	t->4	
ka så	 ->1	d->2	
ka ta	k->1	l->2	n->1	x->1	
ka te	k->1	n->4	r->6	x->1	
ka ti	d->1	g->1	l->29	
ka tj	ä->2	
ka to	l->1	
ka tr	a->2	e->2	u->1	ä->3	ö->1	
ka tv	i->1	
ka ty	d->1	p->3	s->1	
ka tä	c->1	
ka um	g->1	
ka un	d->9	i->242	
ka up	p->7	
ka ut	 ->3	a->1	b->1	f->2	g->2	m->1	s->4	t->5	v->20	
ka va	d->4	l->7	n->3	p->2	r->8	
ka ve	r->15	
ka vi	 ->2	c->1	k->7	l->9	s->2	
ka vo	n->1	t->2	
ka vä	g->1	l->3	n->3	r->6	x->2	
ka vå	r->7	
ka äg	e->1	
ka äm	b->1	
ka än	d->8	
ka är	 ->10	
ka äv	e->2	
ka åk	l->4	
ka åt	a->6	e->2	g->20	
ka öa	r->1	
ka ög	o->1	
ka öp	p->1	
ka ös	t->1	
ka öv	e->7	r->1	
ka", 	v->1	
ka, a	t->1	
ka, b	i->1	
ka, d	e->1	ä->1	
ka, e	l->1	t->1	u->1	
ka, f	r->2	å->1	ö->2	
ka, h	a->2	e->1	
ka, j	o->1	
ka, k	a->1	
ka, m	e->3	å->1	
ka, n	u->1	ä->1	
ka, o	c->4	
ka, r	ä->1	
ka, s	e->1	n->1	o->5	t->1	v->1	
ka, t	i->1	r->1	
ka, v	a->1	i->2	
ka, ä	v->1	
ka, ö	p->1	
ka-ol	y->1	
ka.(I	h->1	
ka.Bo	r->1	
ka.De	 ->1	n->1	t->2	
ka.Ef	t->1	
ka.Em	e->1	
ka.En	 ->2	
ka.Fö	r->1	
ka.He	r->1	
ka.Hu	r->1	
ka.I 	a->1	f->1	l->1	
ka.Ja	g->5	
ka.Lå	t->1	
ka.Me	d->1	
ka.Mi	n->1	
ka.Oc	h->1	
ka.På	 ->2	
ka.Rå	d->1	
ka.Ta	c->1	
ka.Va	r->1	
ka.Ve	m->1	
ka.Vi	 ->3	
ka.Å 	a->1	
ka: "	i->1	
ka: a	t->1	
ka?"J	a->1	
ka?I 	d->1	
kabar	é->1	
kabeh	a->1	
kabek	ä->1	
kabel	.->1	
kabin	e->3	
kad a	n->4	v->3	
kad d	e->1	
kad e	n->1	
kad f	l->1	ö->1	
kad i	n->2	
kad j	ä->1	
kad k	o->6	
kad m	i->1	
kad p	a->1	o->1	r->1	
kad r	ä->1	
kad s	a->1	n->1	y->5	ä->2	
kad t	i->1	r->1	
kad u	p->1	
kad ö	p->1	
kad.D	e->1	
kada 	E->1	d->4	e->1	f->1	k->1	s->1	
kada!	D->1	
kada,	 ->1	
kada.	M->1	
kadad	e->2	
kadan	.->1	a->2	
kadar	 ->6	
kadat	.->1	s->3	
kade 	I->1	a->7	d->2	e->1	f->1	k->4	m->2	o->2	p->4	r->3	s->3	u->1	v->3	ö->1	
kade,	 ->1	
kade.	D->1	H->1	S->1	V->1	
kadee	r->2	
kadef	o->1	
kadem	i->2	
kades	 ->13	,->1	t->1	
kadin	s->1	
kadli	g->10	
kadmi	u->3	
kador	 ->12	,->4	.->2	n->8	
kadra	g->3	
kaffa	 ->19	d->3	n->1	r->1	t->1	
kaffe	n->1	
kafrå	g->1	
kagån	g->4	
kakad	e->1	
kakat	 ->1	
kal a	r->1	
kal b	i->1	
kal f	ö->1	
kal n	i->2	
kal o	m->1	
kal p	o->1	
kal s	i->1	j->1	o->1	
kal: 	p->1	
kala 	a->2	b->1	d->2	e->3	g->2	h->2	i->1	l->2	m->9	o->7	p->4	r->2	s->2	
kala.	K->1	S->1	
kalan	 ->1	.->1	
kaldj	u->1	
kaler	n->1	
kalie	r->4	s->1	
kalig	 ->1	a->2	
kalis	e->4	
kall 	7->1	E->1	a->30	b->73	c->3	d->27	e->3	f->55	g->48	h->41	i->46	j->12	k->71	l->22	m->12	n->7	o->15	p->8	r->5	s->46	t->33	u->28	v->61	ä->6	å->10	ö->10	
kalla	 ->10	d->10	n->6	r->7	t->5	
kalle	l->2	
kallt	,->1	.->1	
kalpa	t->1	
kalt 	b->1	f->1	i->2	t->1	
kalt,	 ->1	
kalt.	J->1	
kalv 	m->1	
kalyd	a->1	
kam f	ö->1	
kam o	m->1	
kam!D	e->1	
kam, 	o->1	
kamli	g->2	
kamma	 ->1	r->59	
kamme	n->1	
kamp 	f->2	i->1	m->5	
kampa	n->6	
kampe	n->16	
kampå	l->1	
kamra	t->1	
kan -	 ->3	
kan A	l->1	
kan E	u->3	
kan I	s->1	
kan a	c->10	g->2	l->1	n->11	r->1	t->5	v->9	
kan b	a->7	e->19	i->9	l->7	y->2	ö->2	
kan d	e->24	o->1	r->4	y->1	ä->4	å->4	ö->1	
kan e	l->1	m->5	n->8	r->4	t->1	x->2	
kan f	a->6	i->6	o->4	r->7	u->2	y->1	å->17	ö->37	
kan g	a->7	e->18	l->1	o->6	å->6	ö->23	
kan h	a->5	e->4	i->4	j->4	o->1	u->3	ä->6	
kan i	 ->8	d->1	f->1	g->1	n->67	s->1	
kan j	a->32	u->1	
kan k	a->2	l->1	o->25	r->2	u->1	ö->1	
kan l	e->10	i->2	o->1	y->4	ä->7	ö->4	
kan m	a->27	e->9	i->1	y->1	ä->1	å->1	ö->1	
kan n	a->2	i->4	o->1	ä->3	å->3	
kan o	c->20	m->9	p->2	r->1	
kan p	l->1	o->1	r->2	å->15	
kan r	e->6	i->2	ä->4	ö->3	
kan s	a->5	e->4	k->11	l->3	o->3	p->5	t->14	ä->13	å->2	
kan t	a->22	i->18	j->1	r->1	y->2	ä->1	
kan u	n->7	p->17	t->18	
kan v	a->29	i->42	ä->4	å->1	
kan ä	g->2	n->2	r->4	v->1	
kan å	s->3	t->9	
kan ö	v->5	
kan, 	g->1	i->1	k->1	o->3	
kan.(	L->1	
kan.D	e->2	ä->1	
kan.O	c->1	
kan.V	å->2	
kanad	e->2	
kanal	,->1	.->2	e->4	y->2	
kanda	l->9	
kande	 ->183	(->1	,->25	.->43	:->3	?->1	n->19	t->85	
kandi	d->14	n->1	
kanen	 ->4	,->1	.->1	
kaner	 ->1	"->1	n->9	
kanik	 ->1	
kanin	e->1	
kanis	m->9	
kanon	e->1	
kans 	a->1	l->1	
kansk	a->10	e->56	t->1	
kansl	e->1	i->1	
kant 	d->1	f->1	o->1	
kant,	 ->2	
kant.	H->1	
kante	n->1	
kaos 	n->1	o->1	
kap -	 ->1	
kap a	t->2	v->20	
kap b	ö->2	
kap d	e->1	ä->2	
kap e	l->1	
kap f	r->1	ö->2	
kap g	r->1	
kap h	a->1	
kap i	 ->5	n->2	
kap k	o->1	
kap m	e->1	å->1	
kap n	ä->1	
kap o	c->12	m->3	
kap s	k->2	o->9	
kap t	i->1	
kap u	n->1	p->1	
kap v	a->1	
kap" 	f->1	
kap"!	I->1	
kap",	 ->1	
kap, 	d->2	e->3	f->2	h->1	i->1	o->3	u->1	v->2	ä->1	
kap. 	S->1	
kap.D	a->1	e->6	
kap.E	u->1	
kap.I	 ->2	
kap.J	a->2	
kap.S	l->1	
kap.T	i->1	
kap.V	i->2	
kap: 	K->1	
kapa 	O->1	a->2	b->3	d->4	e->39	f->8	g->1	h->3	i->3	j->1	k->5	l->1	n->8	o->2	r->1	s->9	t->6	v->1	y->1	ä->1	
kapac	i->5	
kapad	e->5	
kapan	d->24	
kapar	 ->25	.->2	e->2	
kapas	 ->13	
kapat	 ->7	.->1	s->2	
kapen	 ->40	,->7	.->7	s->71	
kaper	 ->4	,->1	.->1	n->16	
kapet	 ->61	)->1	,->13	.->6	?->1	s->15	
kapit	a->17	e->6	u->2	
kapli	g->37	
kapp 	u->1	
kapp,	 ->1	
kapp.	V->1	
kappa	d->3	
kapro	b->1	
kaps 	f->1	
kaps-	 ->1	
kapsa	v->2	
kapsb	e->3	
kapsd	i->1	
kapsf	r->1	
kapsi	n->14	
kapsk	o->3	
kapsl	a->3	
kapsm	a->2	e->1	ä->16	å->1	
kapsn	i->11	
kapso	r->1	
kapsp	e->2	o->2	r->3	
kapsr	a->1	e->9	ä->8	
kapss	t->3	y->1	
kapså	t->2	
kapte	n->2	
kar 1	0->1	
kar F	ö->1	
kar L	a->1	
kar T	h->1	
kar a	l->1	n->3	t->8	v->1	
kar b	e->2	i->1	r->1	
kar d	e->17	r->1	
kar e	l->2	n->1	r->4	u->1	
kar f	a->1	i->2	l->1	r->2	ö->8	
kar g	e->1	
kar h	a->4	e->2	
kar i	 ->7	n->8	
kar j	a->1	
kar k	o->9	r->2	
kar l	a->1	ä->1	
kar m	e->5	i->4	o->1	ä->2	
kar n	ä->1	ö->1	
kar o	c->7	m->2	r->1	
kar p	a->1	å->2	
kar r	e->2	i->1	ä->2	å->3	
kar s	a->1	e->1	i->1	k->1	o->5	t->4	u->2	ä->2	å->1	
kar t	a->1	i->1	
kar u	n->1	p->1	t->2	
kar v	a->7	e->1	i->5	ä->2	å->1	
kar ä	r->1	
kar ö	n->1	v->3	
kar, 	T->1	f->2	k->2	m->1	o->1	s->1	
kar.D	e->1	
kar.E	u->1	
kar.J	a->1	
kar.M	i->1	
kar.O	c->1	
kar.V	i->3	
kar: 	v->1	
kara?	D->1	
karak	t->11	
karan	 ->1	s->5	
kare 	a->2	b->2	f->4	h->1	i->1	j->1	k->1	o->5	s->7	v->2	ä->4	
kare,	 ->9	
kare.	J->1	M->1	
karen	 ->10	.->3	
kares	 ->2	,->1	
kareu	r->1	
karga	 ->1	
karko	n->2	
karla	n->1	
karlä	n->5	
karna	 ->39	!->1	,->1	.->2	s->9	
karpt	 ->2	
karri	ä->2	
kars 	p->1	
karta	 ->1	d->2	
karte	l->13	r->1	
kartl	ä->1	
kas a	t->2	v->8	
kas b	e->1	
kas d	e->1	
kas e	f->2	l->1	n->1	
kas f	r->2	å->1	ö->3	
kas h	a->3	
kas i	 ->3	n->2	
kas k	a->1	l->1	o->1	
kas l	ä->1	
kas m	a->1	e->15	y->1	ä->1	å->1	
kas n	ä->1	å->1	
kas o	c->5	f->1	l->1	r->1	
kas p	o->1	å->1	
kas r	u->1	
kas s	k->1	o->1	
kas t	i->3	
kas u	p->2	t->1	
kas v	a->1	e->1	
kas ä	g->2	r->2	
kas å	s->1	
kas ö	m->1	v->2	
kas!H	e->1	
kas, 	a->1	e->2	i->1	m->2	o->3	p->1	
kas.D	e->1	ä->1	
kas.F	l->1	
kas.H	e->1	i->2	
kas.I	 ->1	n->1	
kas.J	a->1	
kas.M	e->1	
kaska	d->1	
kasmu	g->1	
kasse	r->1	
kasso	r->2	
kast 	a->1	k->1	s->1	t->8	
kast,	 ->1	
kasta	 ->7	n->1	r->3	s->2	t->4	
kaste	 ->9	n->1	t->4	
kastn	i->1	
kasus	 ->3	
kaså 	e->1	h->1	s->1	v->1	
kat -	 ->2	
kat 9	0->1	
kat a	d->1	n->1	t->3	v->2	
kat d	e->2	r->1	
kat e	n->1	t->1	
kat f	r->1	å->1	ö->2	
kat h	o->1	ä->2	
kat i	 ->2	n->1	
kat k	o->1	r->1	
kat m	a->1	e->3	i->1	
kat o	c->4	l->1	m->1	
kat p	å->5	
kat r	e->1	
kat s	i->1	k->1	o->2	t->1	å->1	
kat t	i->1	
kat u	n->1	p->1	t->1	
kat y	t->1	
kat ä	n->1	
kat, 	m->1	n->1	o->1	s->2	u->2	ä->1	
kat.D	e->3	
kat.H	u->2	ä->1	
kat.Ö	v->1	
katal	o->2	y->2	
katas	t->88	
kateg	o->8	
kater	 ->1	.->1	
katio	n->18	
katol	i->4	s->3	
kator	e->4	n->1	
kats 	a->4	f->8	g->4	h->1	i->2	m->2	p->1	s->2	t->1	u->1	å->1	
kats,	 ->1	
kats.	D->1	E->2	
kats?	K->1	
katt 	-->1	f->1	p->1	
katt,	 ->2	
katt.	D->1	P->1	
katta	 ->4	d->4	r->9	
katte	-->1	b->15	f->3	i->2	l->1	n->1	p->1	r->6	s->2	
kattn	i->10	
kavis	a->4	
kay f	ö->2	
kay h	a->1	
kay, 	J->1	a->1	s->1	
kay.V	i->1	
kayDe	 ->1	
kaybe	t->1	
kays 	b->2	
kbar 	s->1	
kbara	 ->3	
kbarh	e->5	
kbart	 ->3	
kbedö	m->4	
kbest	å->4	
kbild	n->1	
kborr	e->1	
kbära	n->1	
kdamm	a->1	
kdel 	f->5	
kdel,	 ->1	
kdel.	E->1	
kdele	n->1	
kdom 	o->1	
kdörr	e->1	
ke (f	i->1	
ke - 	a->1	n->1	s->1	v->1	
ke It	a->1	
ke ag	e->1	
ke an	s->1	
ke at	t->4	
ke ba	k->1	r->1	
ke be	h->2	
ke bi	n->1	
ke bl	a->1	i->1	
ke de	t->4	
ke dy	k->1	
ke då	 ->1	
ke el	l->3	
ke en	 ->2	h->1	l->1	t->1	
ke et	t->1	
ke fi	n->2	
ke fr	a->1	
ke fö	r->6	
ke ge	n->4	
ke gö	r->1	
ke ha	 ->1	r->3	
ke i 	S->1	d->1	f->3	h->1	k->1	n->1	s->1	v->2	
ke in	b->1	o->1	t->8	
ke ka	n->1	
ke ko	m->7	n->1	
ke ku	l->2	
ke kä	n->1	
ke la	g->1	
ke le	d->2	
ke li	b->1	v->1	
ke lä	g->1	t->1	
ke lå	n->1	
ke ma	n->1	
ke me	d->2	n->1	s->1	
ke mi	n->1	
ke må	s->2	
ke na	t->1	
ke ni	 ->1	o->2	
ke oc	h->11	k->3	
ke of	f->1	
ke om	 ->2	b->2	r->1	
ke pr	e->3	
ke på	 ->45	
ke re	g->1	n->1	
ke rö	r->1	
ke se	d->1	
ke sk	u->1	
ke sn	a->1	
ke so	m->8	
ke sp	r->1	
ke sä	g->2	
ke ta	l->1	
ke te	k->1	
ke ti	l->11	
ke ty	c->1	
ke un	d->1	
ke ut	a->2	m->1	r->3	
ke va	r->2	
ke vi	l->3	s->1	
ke vo	r->2	
ke är	 ->10	
ke äv	e->1	
ke ön	s->1	
ke!Äv	e->1	
ke) f	ö->1	
ke) o	c->1	
ke, B	e->1	
ke, S	p->1	
ke, b	å->1	
ke, d	e->3	
ke, f	ö->1	
ke, g	e->1	
ke, h	a->2	e->1	
ke, i	n->1	
ke, k	r->1	
ke, m	e->1	
ke, n	y->1	ö->1	
ke, o	c->3	
ke, s	o->1	
ke, u	n->1	
ke, v	i->2	
ke, å	t->1	
ke-al	b->1	
ke-av	v->1	
ke-da	n->1	
ke-di	s->2	
ke-fo	s->1	
ke-me	t->1	
ke-sp	r->3	
ke-st	a->9	
ke. D	e->1	
ke.- 	(->1	
ke.. 	V->1	
ke..(	E->1	
ke.De	t->5	
ke.Dä	r->1	
ke.Fr	u->2	
ke.Fö	r->2	
ke.He	r->1	
ke.I 	E->1	
ke.Ja	g->2	
ke.Me	n->2	
ke.Ni	 ->1	
ke.Om	 ->1	
ke.Vi	 ->3	d->1	
ke.Ös	t->1	
ke: i	 ->1	
keEn 	v->1	
keFru	 ->1	
keNäs	t->1	
keban	o->1	
ked l	ä->1	
ked o	m->1	
ked t	i->1	
ked.D	e->1	
keda 	f->1	o->1	
kedan	d->1	
kedat	 ->1	
kede 	g->1	o->1	ä->1	
kede.	R->1	
kedet	 ->3	
kedja	 ->1	n->2	
kedjo	r->1	
kedom	 ->2	,->2	a->3	e->3	
kefri	h->1	
keför	h->1	
kegån	g->1	
kekvo	t->1	
kel -	 ->1	
kel 1	 ->2	0->1	1->1	2->2	3->5	4->1	5->3	6->1	
kel 2	.->1	2->1	5->4	8->5	9->2	
kel 3	.->2	0->1	3->2	7->2	9->1	
kel 4	 ->4	.->1	2->1	8->2	
kel 5	 ->1	.->1	0->2	2->1	6->1	
kel 6	 ->9	.->1	2->1	7->1	
kel 7	 ->7	,->1	
kel 8	1->10	2->2	7->2	8->2	
kel 9	.->1	4->1	5->1	
kel a	l->1	n->2	
kel b	ö->1	
kel f	a->1	ö->1	
kel k	a->1	o->1	
kel n	ä->1	
kel o	c->2	m->1	
kel s	o->3	
kel ä	r->3	
kel, 	i->1	o->1	s->1	u->1	
kel.E	u->1	
kel.T	v->1	
kel.V	i->1	
kel.Ä	n->1	
kel: 	U->1	V->1	
kelfr	å->2	
kelfu	n->1	
kelma	j->1	
keln 	f->1	t->5	ä->1	
keln,	 ->1	
kelpr	o->1	
kelri	k->1	
kelro	l->1	
kelse	 ->5	.->1	n->3	r->1	
kelsk	i->1	
kelt 	a->5	d->2	e->3	f->5	g->1	i->2	n->2	o->1	p->1	s->3	t->1	u->2	
kelti	s->1	
kelvä	g->2	
kemed	e->1	
kemik	a->5	
kemis	k->1	t->1	
kemål	 ->3	
kemöj	l->4	
ken (	e->1	
ken -	 ->3	
ken 1	9->2	
ken G	r->1	
ken J	u->1	
ken K	i->2	o->1	
ken S	y->1	ã->1	
ken T	y->3	
ken a	n->1	t->12	v->4	
ken b	e->4	i->1	å->1	ö->1	
ken d	e->2	o->1	
ken e	l->1	n->1	t->2	
ken f	i->1	l->2	o->1	r->5	u->1	å->1	ö->25	
ken g	o->1	r->2	ä->1	
ken h	a->4	j->1	o->1	ä->1	ö->1	
ken i	 ->16	n->14	
ken j	a->2	u->3	
ken k	a->4	n->1	o->3	r->1	
ken l	a->1	i->3	
ken m	a->1	e->12	i->1	o->3	å->7	
ken n	a->1	ä->2	
ken o	c->16	m->7	
ken p	å->17	
ken r	o->1	å->3	
ken s	a->1	k->9	o->10	t->1	u->1	v->1	y->1	ä->2	
ken t	i->10	v->2	
ken u	n->3	p->2	t->5	
ken v	a->2	i->2	ä->1	
ken y	t->1	
ken Ö	s->1	
ken ä	r->4	
ken å	 ->2	s->1	t->2	
ken ö	v->1	
ken, 	L->1	d->2	e->2	f->2	g->3	h->1	i->1	k->1	m->3	n->1	o->4	s->4	t->1	u->1	v->1	y->1	ä->1	
ken. 	O->1	
ken.A	l->1	
ken.B	e->1	
ken.D	e->13	
ken.E	n->1	r->1	t->1	
ken.F	i->1	y->1	ö->1	
ken.H	e->2	ä->1	
ken.I	 ->1	
ken.J	a->5	o->1	
ken.K	o->1	
ken.M	e->2	
ken.P	a->1	
ken.S	o->1	
ken.V	i->1	
ken: 	"->1	J->1	R->1	
ken?F	ö->1	
ken?J	a->1	
ken?V	i->1	
kenHe	r->1	
kens 	b->1	e->1	f->5	g->1	h->1	i->4	k->1	m->1	n->3	o->3	p->1	r->2	s->3	å->1	ö->2	
kensk	a->9	
keomr	å->2	
kepol	i->1	
kepos	i->1	
kepp 	i->1	o->1	
kepps	b->2	r->2	v->2	
kepsi	s->1	
kepti	k->3	s->5	
ker -	 ->1	
ker C	o->1	
ker E	u->1	
ker a	l->5	s->1	t->33	v->2	
ker b	e->4	i->1	o->1	y->2	ö->2	
ker d	e->17	o->2	ä->4	
ker e	n->3	t->2	
ker f	a->1	i->1	l->1	o->1	r->3	ö->4	
ker g	a->1	i->1	r->1	ö->1	
ker h	a->3	e->3	ö->1	
ker i	 ->12	n->16	
ker j	a->15	u->1	
ker k	a->1	o->4	
ker m	a->3	e->7	i->4	y->1	å->3	ö->1	
ker n	e->1	i->3	ä->2	å->1	
ker o	c->13	f->1	m->4	s->2	
ker p	r->2	å->32	
ker r	e->2	ä->2	å->2	
ker s	a->1	i->1	k->3	l->1	o->17	ä->4	å->1	
ker t	i->6	r->1	
ker u	n->1	p->5	t->1	
ker v	a->1	e->2	i->5	å->1	
ker ä	n->2	r->4	
ker ö	v->1	
ker, 	a->1	e->1	h->2	i->2	m->3	n->1	o->1	s->1	t->1	
ker.-	 ->1	
ker.B	e->1	
ker.D	e->4	
ker.G	e->1	
ker.H	ä->2	
ker.M	i->1	
ker.N	ä->1	
ker.P	l->1	
ker.V	i->2	
ker: 	e->1	i->1	
kera 	a->1	s->1	
kerad	 ->2	e->1	
keran	d->1	
kerar	 ->18	
keras	 ->1	
kerat	 ->2	s->1	
keres	u->1	
kerhe	t->235	
kerik	o->1	
kerin	g->5	
kerip	o->1	
keris	e->2	
keriu	t->1	
kerli	g->15	
kern 	E->2	
kerna	 ->21	,->3	.->4	s->2	
kerns	 ->1	
kers 	b->1	u->1	
kerst	ä->24	
kert 	a->1	g->2	h->1	i->4	k->4	l->1	m->1	o->2	p->1	s->5	t->1	v->2	ö->1	
kert!	J->1	
kert,	 ->2	
kerth	e->1	
keräg	a->1	
kerät	t->1	
kes a	n->1	
kes b	e->1	
kes d	e->2	
kes f	i->1	o->2	r->6	
kes i	n->2	
kes k	v->1	
kes n	y->1	
kes o	b->1	c->1	m->1	
kes p	r->1	
kes r	e->2	
kes s	i->1	l->1	
kes v	ä->1	
kes- 	o->4	
kesar	b->1	
kesek	t->1	
keset	i->1	
kesfr	å->4	
kesfö	r->1	
kesha	n->4	
kesis	k->1	
keska	r->1	
keskv	a->1	
kesla	g->2	
kesli	v->2	
kesmi	n->9	
kesmä	s->1	
kespo	l->3	
keste	i->1	
kesut	b->7	
kesva	l->1	
ket (	E->2	I->1	
ket -	 ->2	
ket B	e->1	
ket E	u->2	
ket G	r->1	
ket P	o->1	
ket V	a->1	
ket a	k->2	l->7	m->1	n->8	r->4	t->20	v->9	
ket b	a->2	e->9	l->3	o->1	r->6	ä->1	
ket d	e->8	r->1	y->1	å->1	
ket e	g->2	n->7	r->1	t->1	u->2	x->3	
ket f	a->13	i->2	l->1	o->2	r->2	u->1	å->2	ö->21	
ket g	a->1	e->3	j->1	l->5	o->6	r->4	ä->2	ö->4	
ket h	a->7	e->3	i->2	å->1	ö->6	
ket i	 ->6	l->1	m->1	n->26	r->1	
ket j	a->6	u->2	ä->2	
ket k	a->2	l->5	o->21	r->5	u->1	v->2	ä->6	
ket l	a->2	e->1	i->9	ä->13	å->4	
ket m	a->4	e->18	i->1	o->1	å->2	ö->1	
ket n	a->1	e->1	i->1	o->7	u->1	y->2	ä->1	å->2	ö->1	
ket o	c->12	f->1	g->1	m->11	n->2	p->2	r->6	s->1	t->2	
ket p	a->3	e->2	l->1	o->11	å->8	
ket r	a->1	e->7	i->6	å->1	ö->1	
ket s	a->2	e->4	i->1	j->2	k->15	m->1	n->5	o->8	p->2	t->42	v->6	y->6	ä->9	å->1	
ket t	i->7	r->4	u->3	y->9	
ket u	n->1	p->7	r->1	t->6	
ket v	a->6	e->1	i->60	o->1	ä->22	å->2	
ket ä	g->1	n->1	r->21	
ket å	t->2	
ket ö	v->1	
ket!(	P->1	
ket, 	D->1	I->1	J->1	W->1	e->1	f->6	g->1	h->6	i->1	k->1	m->4	o->5	s->2	t->1	u->2	ä->1	
ket.D	e->1	ä->1	
ket.E	t->1	u->1	
ket.I	 ->1	
ket.J	u->1	
ket.M	e->2	
ket.N	ä->1	
ket.O	c->1	
ket.S	k->1	
ket.V	i->1	
ket: 	v->1	
ket; 	D->1	a->1	u->1	
ket?O	c->1	
ketet	 ->2	.->1	
ketin	g->2	
ketma	t->1	
ketry	c->3	
kets 	d->1	f->1	k->1	o->1	r->6	s->3	u->1	
kett 	e->4	g->1	i->3	o->1	s->2	u->2	
kett,	 ->1	
kett.	 ->1	
kevat	t->2	
kfakt	o->1	
kfart	y->7	
kford	o->1	
kfrit	t->2	
kfron	t->1	
kfyll	t->1	
kföre	b->1	n->7	
kförh	å->1	
kförs	ä->1	
kförv	a->1	
kgilt	i->2	
kgrun	d->31	
kgrup	p->2	
kh ha	r->1	
kh-av	t->1	
kh.De	t->1	
kh.Fö	r->1	
khant	e->6	
kheer	 ->3	,->4	J->1	b->3	s->3	
khet 	a->1	b->1	e->3	i->2	m->20	o->1	s->2	
khet,	 ->1	
khet.	 ->1	F->1	
khete	n->3	r->5	
kholm	 ->1	,->1	.->1	
khus 	1->1	
khus,	 ->2	
khus.	G->1	
khuse	t->2	
khusl	ä->1	
khäls	a->9	
ki Li	i->2	
ki.De	t->1	
kick 	d->1	o->2	
kick.	D->1	
kicka	 ->4	d->2	r->3	s->1	t->2	
kickl	i->1	
kidna	p->1	
kien 	o->1	s->1	
kien,	 ->1	
kiet 	D->1	I->1	a->1	e->1	f->1	h->7	i->2	n->2	o->3	p->1	s->3	t->1	v->1	ä->2	
kiet,	 ->2	
kiet.	D->1	O->1	
kiets	 ->4	
kifte	 ->1	,->1	.->1	t->3	
kig s	a->1	
kigt 	E->1	n->3	
kild 	b->2	f->2	i->1	k->3	m->1	o->1	p->1	r->2	t->2	u->2	
kild.	F->1	
kilda	 ->35	s->2	
kilde	 ->2	,->1	.->1	
kildr	a->3	
kilja	 ->4	k->4	s->2	
kilje	d->1	f->1	l->1	r->7	
kiljt	 ->1	
killi	g->2	
killn	a->44	i->1	
kilo 	g->1	m->1	o->1	
kilo,	 ->1	
kilom	e->1	
kilt 	E->2	S->2	a->3	b->9	d->7	e->3	f->14	g->4	h->3	i->11	j->1	k->3	l->1	m->11	n->5	o->2	p->8	s->5	t->12	u->4	v->17	ä->2	å->1	
kin o	c->2	
kin s	o->2	
kin.D	e->1	
kinen	 ->1	s->1	
kiner	i->1	
kines	e->2	i->7	
king 	o->1	
kingr	a->2	i->1	
kinli	g->1	
kipa 	r->2	
kipan	d->1	
kipni	n->9	
kirer	.->1	
kis f	r->1	
kis i	 ->1	
kis p	å->1	
kis! 	V->1	
kisbe	t->1	
kisk 	a->1	b->1	l->1	n->1	o->1	p->2	
kiska	 ->57	
kiske	 ->3	
kiss 	f->1	
kisse	r->3	
kista	n->12	
kit a	t->1	v->1	
kit f	r->1	
kit t	i->1	
kitin	 ->1	.->1	
kits 	f->1	
kiv l	ä->1	
kiver	a->1	
kjuta	 ->9	n->1	s->3	
kjute	n->2	r->5	
kjuti	t->5	
kjuts	 ->5	
kjutv	a->1	
kkapi	t->1	
kki L	i->2	
kkomm	u->2	
kkunn	i->1	
kkuns	k->1	
kkuyu	 ->2	
kköy 	-->1	
kl. 1	1->6	2->6	3->1	5->2	7->1	9->1	
kl. 2	0->1	1->2	
kl.12	.->1	
kla a	r->1	v->1	
kla d	e->2	
kla e	k->1	n->7	t->2	
kla f	r->1	ö->2	
kla h	e->1	
kla i	n->1	
kla k	o->1	
kla l	i->1	
kla n	a->1	y->2	ä->1	
kla o	c->5	
kla r	e->1	
kla s	i->2	k->2	o->1	t->1	
kla t	j->1	
kla u	t->1	
kla v	i->1	
kla ö	s->1	
kla.M	e->1	
klad 	h->1	m->1	
klade	 ->9	s->1	
klaga	 ->7	!->1	.->1	d->2	n->8	r->59	t->1	
klage	l->3	
klagl	i->8	
klago	m->3	s->1	
klam 	f->2	
klame	r->1	
kland	 ->16	)->1	,->11	.->5	e->7	s->3	
klang	,->1	
klapp	j->1	s->1	
klar 	-->1	a->4	b->2	d->1	e->2	i->2	m->3	o->1	p->1	r->3	t->2	u->2	ä->1	
klar,	 ->4	
klar.	J->1	M->1	
klara	 ->36	,->1	.->2	d->5	r->29	s->5	t->5	
klare	 ->3	
klarg	ö->17	
klarh	e->12	
klari	n->24	
klarl	a->3	ä->2	
klarn	a->12	
klart	 ->86	,->2	.->1	:->1	e->7	
klas 	a->1	e->1	i->4	m->1	o->3	p->3	s->3	v->1	y->2	
klas.	D->3	
klas:	 ->1	
klass	 ->2	a->1	e->3	i->15	p->1	
klast	 ->1	e->1	
klat 	a->2	
klat,	 ->1	
klats	 ->3	.->1	
klaus	u->6	
klave	r->1	
kled 	m->1	
kleri	 ->3	e->1	
klern	a->1	
klet 	g->1	
klibb	i->1	
klien	t->1	
klig 	a->2	e->1	f->3	h->3	j->1	k->5	l->2	m->5	o->1	r->1	s->4	t->2	u->7	v->1	
klig,	 ->2	
klig.	 ->1	D->1	
kliga	 ->84	.->2	d->1	n->4	s->4	t->2	
klige	n->147	
kligh	e->29	
kligt	 ->54	,->4	.->7	v->5	
klima	t->14	
kling	 ->60	,->17	.->11	a->1	e->53	s->35	
kloak	l->1	
klock	a->2	
kloka	 ->1	s->1	
klokt	 ->5	
klude	r->4	
klukt	 ->1	
klusi	v->20	
klyft	a->2	o->3	
klyve	r->1	
klägg	a->1	
klöst	 ->1	
km lå	n->1	
km mi	n->1	
km, t	i->1	
km.Tr	o->1	
kmeni	s->2	
kmete	r->2	
kmode	l->1	
kna d	e->2	
kna i	n->1	
kna m	e->4	
kna s	a->1	
kna t	a->1	
kna u	p->3	
kna v	å->1	
kna, 	s->1	
kna.V	i->1	
knad 	a->2	f->1	h->1	i->2	k->1	s->2	
knad,	 ->6	
knad.	D->1	E->1	
knade	 ->3	n->133	r->17	s->5	
knads	a->4	d->1	e->14	i->1	k->1	l->1	m->2	o->1	p->3	v->1	
knand	e->20	
knapp	 ->1	a->11	t->4	
knar 	E->1	R->1	a->1	b->2	d->2	e->3	j->2	k->1	m->15	o->3	t->1	u->1	v->3	å->1	
knas 	a->5	b->1	e->2	f->1	g->1	i->4	j->1	l->1	o->1	p->1	s->5	t->2	
knas,	 ->3	
knas.	E->1	V->1	
knat 	e->1	i->3	k->1	m->1	o->3	s->1	u->1	
knat,	 ->1	
knats	 ->6	,->1	
kneex	e->1	
kneli	g->1	
knes 	e->1	
knik 	D->1	s->4	u->1	
knike	n->4	r->3	
kning	 ->127	"->2	,->14	.->17	a->41	e->73	s->75	
knipa	.->1	
knipp	a->3	
knisk	 ->14	a->18	t->4	
knivå	 ->1	
knolo	g->3	
know-	h->1	
knuss	l->1	
knute	n->3	t->1	
knutn	a->2	
knutp	u->1	
knyta	 ->5	
knyte	r->2	
knytn	i->1	
knyts	 ->1	
knäck	a->2	
ko Ca	d->5	
ko, A	s->1	
ko.Ty	 ->1	
koali	t->14	
kod f	ö->5	
kod h	a->1	
kod k	o->1	
koden	 ->1	.->2	
koder	 ->2	,->1	
kodif	i->2	
koeff	i->1	
koffe	r->1	
kofin	-->2	
koför	a->1	f->1	
kog e	v->1	
kog f	r->1	
kog i	n->1	
kogar	 ->1	,->1	.->1	n->7	
kogen	 ->1	,->2	.->2	
kogri	k->1	
kogsa	r->1	v->1	
kogsb	r->6	
kogsf	a->1	
kogsk	o->1	
kogso	m->1	
kogsp	o->1	
kogss	e->4	
kogsu	t->1	
kogsv	å->1	
kogsä	g->2	
kogår	d->1	
kohan	d->3	
koher	e->1	
kohol	,->1	
koka 	s->1	
kokor	 ->1	
kol- 	o->1	
kola 	f->1	ä->1	
kolan	 ->2	,->1	.->1	
koldi	o->5	
kolen	.->1	
kolib	a->1	
koliv	 ->2	.->1	
koll 	f->1	i->2	o->1	s->2	
koll.	D->1	J->1	V->1	
kolle	g->195	k->10	n->1	t->16	
kolli	s->3	
kolog	i->16	
kolon	i->1	
kolor	 ->2	,->1	
kolos	s->1	
kom -	 ->1	
kom a	t->1	
kom d	e->10	å->2	
kom e	r->1	
kom f	l->1	r->4	ö->2	
kom h	i->1	
kom i	 ->1	n->2	
kom l	j->1	
kom m	a->1	e->1	i->1	o->1	
kom n	u->1	
kom o	s->3	
kom p	r->2	
kom r	e->1	y->1	å->1	
kom s	a->1	
kom t	i->2	
kom u	t->1	
kom v	i->1	
kom ö	v->3	
kom, 	n->1	
kom.D	e->1	
koman	e->1	
kombi	n->1	
komli	g->9	
komma	 ->101	,->1	.->2	n->55	s->1	
komme	l->15	n->84	r->718	t->5	
kommi	s->1044	t->102	
kommu	n->32	
komna	 ->13	,->1	.->1	n->1	r->28	s->1	
kompe	n->10	t->11	
kompl	e->28	i->16	
kompo	n->4	
kompr	o->21	
kområ	d->10	
komrö	s->6	
komst	 ->7	e->8	f->1	h->1	k->1	
kon a	v->1	
konad	e->1	
konar	 ->1	
konce	n->31	p->7	r->2	
konci	s->2	
konfe	d->1	r->170	s->1	
konfi	d->2	s->2	
konfl	i->16	
konfr	o->1	
kongr	e->1	
konju	n->1	
konkr	e->57	
konku	r->272	
konom	e->4	i->282	
konse	k->60	r->7	
konso	l->3	
konst	 ->1	,->1	a->40	i->25	r->36	
konsu	l->5	m->60	
konta	k->17	m->2	n->1	
konte	x->1	
konti	n->7	
konto	r->7	
kontr	a->7	o->182	
konve	n->22	r->5	
koope	r->1	
kop b	e->1	
kop, 	A->3	
kopia	 ->1	
kopie	r->1	
kopou	l->5	
koppl	a->4	i->2	
kor -	 ->1	
kor a	t->1	v->1	
kor d	e->1	ä->2	ö->1	
kor e	f->1	
kor f	a->1	i->1	o->1	r->3	ö->15	
kor h	a->2	i->1	
kor i	 ->10	n->3	
kor l	e->1	i->1	
kor m	e->2	å->1	
kor n	ä->1	
kor o	c->6	
kor p	å->1	
kor s	e->3	k->2	o->20	
kor t	i->5	
kor u	t->2	
kor v	a->2	i->1	
kor ä	n->1	r->2	
kor, 	e->1	f->1	k->2	m->2	o->1	r->1	s->3	v->1	
kor.B	r->1	
kor.D	e->4	
kor.E	t->1	
kor.G	e->1	
kor.J	a->1	
kor.T	i->1	
kor.Ö	V->1	
koran	d->1	
kord 	b->1	
kordt	i->1	
korea	 ->1	
koren	 ->16	,->1	.->4	
korli	g->2	
korna	 ->24	,->2	.->5	s->3	
korre	k->27	s->1	
korri	d->2	
korru	m->2	p->7	
kors 	a->1	d->1	f->2	h->3	i->1	l->1	o->1	r->1	s->2	t->1	y->1	
kort 	E->1	a->1	b->1	d->3	f->10	g->3	i->2	k->2	l->1	n->1	o->4	p->4	r->2	s->11	t->5	u->2	v->2	
kort,	 ->3	
kort.	D->2	E->1	J->2	
kort:	 ->1	
kort?	J->1	
korta	 ->4	d->1	s->1	
korte	n->1	t->19	
kortf	a->2	
kortn	i->1	
korts	i->4	
kosam	t->1	
koslä	k->1	
kosta	 ->2	d->2	r->4	t->1	
kosth	å->1	
kostn	a->104	
kosts	a->2	
kosys	t->4	
kotik	a->7	
kott 	a->2	b->1	d->1	e->2	f->5	i->2	o->1	s->5	u->1	
kott,	 ->2	
kott.	D->1	L->1	M->1	O->2	
kotte	n->3	t->132	
kottl	a->5	
kotts	 ->2	b->2	d->1	
kouri	.->1	
kov n	y->1	
kov o	c->1	
kovet	 ->1	
kpart	i->10	
kprob	l->1	
kprov	s->3	
kra a	t->1	
kra d	i->1	
kra e	n->1	r->11	
kra f	ö->1	
kra g	r->1	
kra h	u->1	
kra i	 ->1	
kra k	o->1	
kra m	e->1	
kra o	c->1	r->2	s->3	
kra p	l->1	å->4	
kra s	i->1	o->1	t->1	ä->1	
kra v	i->1	
kra ö	p->1	
krad 	i->1	
krade	 ->2	
kraft	 ->38	,->9	.->5	?->2	e->26	f->12	i->34	s->10	t->5	v->8	
krans	.->1	
krar 	a->1	e->1	f->1	s->1	
krar.	J->1	
krare	 ->2	
krarn	a->3	
kras.	J->1	
krasc	h->3	
krass	t->1	
krast	e->5	
krat 	h->1	s->1	
krate	r->23	s->1	
krati	 ->14	"->1	,->3	.->9	e->3	f->1	n->20	r->1	s->91	
kratt	a->1	r->1	
krav 	-->1	b->1	f->4	g->1	i->1	l->1	n->1	o->3	p->16	s->8	t->1	u->1	
krav,	 ->4	
krav.	(->1	.->1	D->2	E->1	R->1	
krav?	V->1	
krava	l->1	
krave	n->25	t->15	
kreat	i->2	ö->1	
kredi	t->2	
krege	r->1	
kreng	ö->2	
krepu	b->3	
krera	 ->1	
kret 	b->1	e->1	f->3	h->1	i->2	k->1	o->2	p->1	s->2	t->3	u->2	
kret:	 ->1	
kreta	 ->36	r->3	
krete	r->2	s->12	
kreti	s->2	
krets	 ->2	,->1	a->3	e->2	l->2	
krev 	d->1	i->1	n->1	o->1	t->1	u->1	
krevs	 ->2	
krida	n->12	
kride	r->7	
krids	 ->2	
krift	 ->2	e->12	l->8	
krig 	m->1	o->1	p->1	s->2	v->1	
krig"	.->1	
krig,	 ->1	
krig.	J->1	
krige	t->12	
krigs	h->1	s->1	
krik.	G->1	
krike	 ->24	,->8	.->1	:->1	s->5	
krikt	a->2	n->2	
krimi	n->27	
kring	 ->30	a->7	g->2	s->16	
kris 	h->1	i->1	m->1	s->1	u->1	v->1	ä->1	
kris?	Ä->1	
krise	n->6	r->3	
krism	e->2	
kriso	m->1	
kriss	i->1	t->1	
krist	a->2	d->11	
krita	n->1	
krite	r->21	
kriti	k->16	s->32	
kriva	 ->8	n->2	s->1	
krivb	o->1	
krive	l->5	n->4	r->14	t->2	
krivi	t->8	
krivn	a->3	i->5	
krivs	 ->8	
kroat	e->1	
kroek	o->5	
krofi	n->1	
krofö	r->1	
krokr	e->2	
krom 	g->1	
krom,	 ->1	
kroma	d->1	
kronj	u->1	
kropp	e->1	
kross	a->1	
krost	a->1	
krot.	J->1	
krota	 ->1	d->2	r->2	s->5	
krotf	ä->1	
krotn	i->15	
krov 	f->3	o->2	s->1	
krov"	,->1	
krov,	 ->1	
krov.	 ->1	D->1	
krove	t->3	
krovk	o->1	
krovs	i->1	
kry.D	e->1	
krygg	a->1	
kryph	å->3	
krypt	o->2	
kryss	a->1	
kryte	r->1	
kräck	 ->1	a->2	e->1	l->2	n->1	s->1	t->1	
krädd	a->1	
kräft	a->29	e->1	
kräkt	a->1	
krämd	 ->1	
kräml	i->1	
krämm	a->1	e->2	
kränk	a->2	b->1	e->5	n->13	s->3	t->5	
kräpn	i->1	
krätt	e->1	
kräva	 ->27	n->2	s->5	
krävd	e->4	
kräve	r->44	
krävs	 ->52	,->3	
krävt	 ->1	s->1	
krång	e->1	l->1	
kröna	s->1	
ks an	s->1	
ks av	 ->3	
ks be	s->1	t->1	
ks de	 ->1	s->1	
ks do	k->1	
ks ef	t->1	
ks fr	i->1	
ks ge	n->1	
ks in	t->1	
ks mi	g->1	n->1	
ks må	l->1	
ks na	t->1	
ks oc	h->4	k->1	
ks om	 ->1	
ks pa	p->1	
ks pe	r->1	
ks re	f->1	
ks sa	m->1	
ks so	c->1	
ks st	r->1	
ks su	v->1	
ks ti	d->1	l->1	
ks ty	d->1	
ks up	p->1	
ks ut	t->1	
ks va	r->1	
ks ve	r->1	
ks vi	s->1	
ks öv	e->1	
ks, d	å->1	
ks.Dä	r->1	
ks.OL	A->1	
ks.På	 ->1	
ks.Ut	m->1	
ks.Vi	 ->1	
ks; d	e->1	
ksake	r->1	
ksam 	d->1	f->2	n->1	o->3	p->4	u->1	ö->1	
ksam.	I->1	
ksamh	e->88	
ksamm	a->20	
ksamt	 ->6	,->1	
ksanl	ä->1	
ksbor	d->1	
ksbåd	a->1	
kscen	a->1	
ksche	f->1	
ksdra	b->3	
kseko	n->1	
ksekr	e->1	
ksfal	l->2	
ksfon	d->1	
ksfrå	g->1	
ksilv	e->3	
kskör	t->1	
kslob	b->1	
kslut	 ->1	
ksodl	i->1	
ksom 	A->1	B->1	F->1	a->9	b->2	c->1	d->8	e->5	f->6	h->1	i->2	j->1	m->4	n->2	o->3	p->2	s->3	v->2	ä->1	
ksomr	å->2	
kson 	f->1	i->1	
kspol	i->6	
kspri	n->1	
kspro	d->2	
ksref	o->1	
ksreg	i->1	
ksris	k->2	
kssek	t->5	
kssyn	p->1	
kstan	,->1	
kstav	l->1	
kstyr	e->1	
kstäd	e->1	
kstäl	l->21	
ksvat	t->1	
kswag	e->1	
ksägn	e->1	
kså "	m->1	
kså -	 ->2	
kså 1	9->1	
kså E	u->3	
kså F	l->1	
kså M	o->1	
kså a	b->1	k->1	l->4	n->9	r->1	t->49	v->8	
kså b	a->3	e->13	i->1	l->1	o->2	r->1	y->1	ä->2	ö->4	
kså d	e->21	i->1	o->1	ä->2	
kså e	k->1	n->21	r->1	t->9	
kså f	a->2	i->3	o->1	r->7	u->2	å->5	ö->23	
kså g	a->1	e->4	l->1	o->2	ä->3	å->3	ö->4	
kså h	a->10	e->7	o->2	u->3	ä->3	å->1	
kså i	 ->22	a->1	n->14	
kså j	a->1	
kså k	a->8	l->3	o->18	r->2	u->1	ö->1	
kså l	i->1	y->1	
kså m	e->17	i->3	o->1	y->4	å->11	ö->2	
kså n	o->2	y->1	ä->3	å->5	ö->2	
kså o	a->2	c->1	m->7	r->1	
kså p	a->2	e->1	l->1	å->14	
kså r	a->1	e->2	å->1	ö->2	
kså s	a->4	e->5	k->13	l->1	n->1	o->3	p->1	t->7	v->1	ä->11	å->1	
kså t	a->16	i->11	o->1	r->1	y->1	ä->1	
kså u	n->4	p->9	t->5	
kså v	a->13	e->2	i->16	ä->1	å->3	
kså z	i->1	
kså ä	g->1	n->2	r->17	
kså å	t->3	
kså ö	v->3	
kså, 	e->1	f->1	h->1	i->1	m->1	o->4	s->1	
kså.D	e->1	
kså.I	n->1	
kså.J	a->1	
kså.N	i->1	
kså.P	å->1	
ksöde	 ->1	
kt (8	0->2	
kt - 	e->1	n->1	o->1	v->1	
kt -,	 ->1	
kt 1 	u->1	
kt 1,	 ->1	
kt 11	 ->1	
kt 2 	i->2	
kt 26	 ->1	
kt 4 	i->1	l->1	
kt 5,	 ->1	
kt 6 	o->1	
kt 7 	i->1	
kt D 	k->1	
kt EU	 ->1	.->1	
kt Eu	r->4	
kt Fl	o->1	
kt Fr	a->1	
kt Ko	s->1	
kt Mü	n->1	
kt ab	s->1	
kt al	l->1	
kt an	a->2	s->5	
kt ar	b->3	
kt at	t->46	
kt av	 ->6	
kt ba	k->1	x->1	
kt be	d->2	g->2	k->1	r->3	s->2	t->6	v->1	
kt bi	d->3	n->3	s->6	
kt bl	i->3	
kt br	y->1	
kt bu	d->1	
kt by	g->2	
kt bä	t->1	
kt ch	a->1	
kt ci	v->1	
kt d)	 ->1	
kt da	t->1	
kt de	 ->1	c->1	f->2	m->1	n->2	p->1	t->4	
kt do	k->1	
kt dr	a->1	
kt dä	r->4	
kt e)	 ->1	
kt ef	t->1	
kt eg	e->2	
kt ek	o->1	
kt el	l->2	
kt en	 ->3	g->1	
kt er	 ->1	f->1	k->1	s->1	t->1	
kt et	t->3	
kt ex	e->2	
kt fa	k->2	l->1	s->1	
kt fe	l->1	m->1	n->1	
kt fi	n->3	
kt fl	y->1	
kt fr	a->1	e->1	i->1	å->3	
kt fu	l->1	
kt fy	r->1	
kt fä	n->1	
kt få	 ->4	t->1	
kt fö	r->56	
kt ge	n->2	
kt gr	a->2	ö->1	
kt gä	l->3	
kt gå	 ->2	
kt gö	r->3	
kt ha	d->1	n->3	r->13	
kt he	l->1	
kt hi	n->1	
kt hu	n->1	r->3	
kt hä	n->1	r->1	
kt hå	l->2	
kt i 	M->1	b->1	d->3	e->1	f->2	h->2	j->1	m->1	r->1	s->1	
kt in	b->1	f->3	g->1	i->2	n->3	o->2	s->2	t->12	
kt is	o->2	
kt ju	s->1	
kt ka	l->1	n->6	s->1	
kt kl	a->3	
kt ko	m->7	n->4	r->2	
kt ku	l->1	n->2	
kt kv	a->1	
kt kä	n->1	
kt la	b->1	g->1	n->2	
kt le	d->1	v->1	
kt ly	c->1	
kt lä	g->2	n->1	t->1	
kt ma	n->1	r->2	t->1	
kt me	d->17	l->1	n->3	
kt mi	l->1	n->2	s->4	
kt mo	d->1	t->5	
kt my	c->3	
kt må	n->1	
kt mö	j->1	
kt ny	l->1	
kt nä	r->5	
kt nö	d->1	t->1	
kt oc	h->42	
kt om	 ->12	.->1	d->1	o->1	
kt op	e->1	
kt or	g->1	
kt pa	r->4	
kt pe	r->3	
kt po	l->3	
kt på	 ->41	d->1	
kt ra	t->1	
kt re	l->1	p->1	s->1	
kt ri	s->1	
kt rä	t->2	
kt rö	s->1	
kt sa	m->6	
kt se	 ->1	t->9	
kt si	g->1	n->2	
kt sk	a->5	e->1	r->1	u->3	y->1	
kt sm	i->1	
kt so	m->42	
kt sp	e->1	
kt st	a->3	o->1	ä->2	å->1	ö->9	
kt sv	a->2	å->1	
kt sy	f->1	s->1	
kt sä	t->18	
kt så	 ->1	
kt ta	g->5	l->1	
kt te	r->1	
kt ti	l->9	
kt to	m->1	
kt tr	e->1	
kt tv	å->2	
kt un	d->1	
kt up	p->5	
kt ur	s->3	
kt ut	,->2	a->2	b->1	k->1	m->1	n->1	o->1	t->1	v->1	
kt va	d->2	l->6	r->3	t->2	
kt ve	r->2	
kt vi	d->9	k->1	l->5	n->1	s->3	
kt vä	r->3	
kt vå	r->1	
kt äm	n->1	
kt än	 ->4	n->1	
kt är	 ->15	,->1	.->1	
kt äv	e->2	
kt åt	a->1	
kt ög	o->1	
kt öl	 ->1	
kt öv	e->4	
kt!Nä	r->1	
kt", 	e->1	
kt, "	e->1	
kt, a	r->1	
kt, b	o->1	
kt, d	e->2	
kt, e	f->1	l->1	n->2	t->1	
kt, f	o->1	ö->2	
kt, g	l->1	
kt, i	 ->1	
kt, l	å->1	
kt, m	e->6	o->1	å->1	
kt, n	ä->2	
kt, o	b->1	c->4	m->1	
kt, r	a->1	
kt, s	o->3	ä->1	
kt, t	.->1	r->1	
kt, u	t->2	
kt, v	a->1	i->3	
kt, ä	r->1	v->1	
kt. D	e->1	
kt.(P	r->1	
kt.Al	l->1	
kt.Av	s->1	
kt.Be	t->1	
kt.Bo	r->1	
kt.Bå	d->2	
kt.De	 ->3	n->5	s->2	t->7	
kt.Di	r->1	
kt.Dä	r->1	
kt.Då	 ->1	
kt.Fe	l->1	
kt.Fö	r->1	
kt.Ge	n->1	
kt.He	r->1	
kt.I 	d->1	f->1	v->1	
kt.Ja	g->6	
kt.Ko	m->1	
kt.Ma	n->3	r->1	
kt.Me	n->1	
kt.Mi	n->1	
kt.Må	n->1	
kt.Nu	 ->1	
kt.Nå	g->1	
kt.Oc	h->1	
kt.Om	 ->3	
kt.Pr	e->1	
kt.Re	g->1	
kt.Sl	u->2	
kt.Ta	c->1	
kt.Ti	l->1	
kt.Un	g->1	
kt.Va	d->1	r->2	
kt.Vi	 ->2	
kt.Vå	r->1	
kt.Å 	a->1	
kt: J	a->1	
kt: V	i->1	
kt: d	e->1	
kt: u	t->1	
kt; e	n->1	
kt; å	 ->1	
kt?Eu	r->1	
kt?Tä	n->1	
kt?Ut	g->1	
kta a	l->1	n->3	r->2	t->2	
kta b	e->10	i->2	
kta d	e->5	ö->1	
kta e	f->1	l->1	r->2	t->3	
kta f	å->2	ö->2	
kta g	i->1	o->1	
kta h	o->1	
kta i	 ->1	d->1	n->1	
kta k	o->4	r->1	
kta m	e->1	i->1	y->1	
kta o	c->2	s->2	
kta p	o->1	r->1	å->2	
kta r	a->2	e->4	ö->1	
kta s	a->1	i->4	j->1	k->1	l->2	o->3	t->1	ä->1	
kta t	o->1	
kta u	n->1	p->4	r->1	t->1	
kta v	a->1	i->1	
kta, 	j->1	s->1	
kta.F	ö->1	
kta.J	a->3	
ktabe	l->2	
ktabi	l->1	
ktad 	a->1	f->2	m->1	p->2	
ktad.	H->1	J->1	
ktade	 ->12	,->1	s->1	
ktadm	i->2	
ktaga	n->1	
ktain	s->2	
ktake	l->2	
ktaku	l->1	
ktala	n->1	
ktan 	a->1	p->4	
ktand	e->6	
ktans	v->7	
ktar 	a->2	b->1	d->4	f->1	i->1	m->1	o->1	s->5	u->4	v->1	ö->1	
ktar,	 ->1	
ktar.	F->1	M->1	
ktare	 ->6	,->1	n->6	
ktarn	a->6	
ktas 	a->1	d->2	i->4	m->2	p->1	s->5	u->1	v->2	
ktas.	B->1	
ktat 	d->2	k->1	m->1	o->2	p->2	s->4	ä->1	
ktat,	 ->2	
ktat.	D->1	
ktato	r->1	
ktats	 ->4	,->1	.->1	
ktatu	r->2	
ktbal	a->2	
ktbar	h->1	t->2	
ktbef	o->2	
ktdel	n->1	
ktdik	t->1	
kte E	u->1	
kte J	o->1	
kte a	t->4	v->1	
kte d	e->2	
kte e	n->1	
kte i	 ->1	n->1	
kte j	a->1	
kte k	r->1	
kte m	i->2	
kte o	c->1	m->1	
kte p	å->1	
kte s	e->1	i->2	o->4	v->1	
kte t	i->2	
kte u	t->1	
kte v	ä->1	
kte, 	e->1	f->1	k->1	
kte.F	ö->1	
kte.M	a->1	
ktels	e->13	
kten 	-->3	a->29	b->3	d->3	e->1	f->16	g->9	h->5	i->10	k->2	l->1	m->2	n->3	o->10	p->4	s->17	t->1	u->2	v->8	ä->11	ö->6	
kten,	 ->16	
kten.	 ->2	A->1	D->9	F->1	H->2	I->1	J->2	M->2	O->2	P->1	S->1	U->1	V->2	Ä->1	Ö->1	
ktens	 ->3	k->1	
kter 	-->1	a->11	b->3	d->2	e->1	f->8	g->1	i->12	j->1	k->1	m->8	n->3	o->11	p->9	s->23	t->2	u->1	v->5	ä->6	
kter,	 ->20	
kter.	 ->1	)->1	D->3	E->1	F->8	H->1	J->2	M->1	P->1	T->1	V->1	
kter:	 ->2	
kter?	H->1	T->1	
ktera	 ->12	,->1	.->1	d->2	r->15	s->9	
kteri	e->1	s->2	
ktern	a->31	
ktert	 ->2	
ktes 	a->3	e->1	m->1	
ktet 	K->1	a->2	c->1	e->1	f->2	h->1	k->1	m->2	p->1	u->1	ä->1	
ktet,	 ->1	
ktets	 ->1	
ktfar	t->1	
ktför	e->1	l->1	
kthav	a->1	
kthet	.->1	
kthål	l->1	
ktieb	ö->1	
ktieä	g->2	
ktig 	-->2	b->3	d->7	f->18	g->2	h->3	i->2	j->1	k->5	l->2	m->4	o->6	p->9	r->10	s->3	t->5	u->3	å->1	
ktig,	 ->7	
ktig.	D->4	I->1	J->3	M->2	N->1	
ktig?	J->1	
ktiga	 ->91	,->4	.->2	d->1	r->10	s->43	t->2	
ktigh	e->65	
ktigt	 ->144	,->14	.->10	
ktik 	e->1	
ktik,	 ->1	
ktike	n->10	
kting	a->12	e->1	f->1	
ktinn	o->1	
ktinv	e->1	
ktion	 ->34	"->1	,->5	.->10	a->2	e->39	i->4	s->29	
ktisk	 ->2	,->1	a->19	t->52	
ktiv 	(->1	-->1	9->8	a->2	b->2	d->2	e->7	f->6	h->7	i->6	k->7	l->3	m->3	o->24	p->5	r->1	s->22	t->2	u->1	v->4	ä->4	å->2	ö->1	
ktiv,	 ->15	
ktiv.	A->1	D->4	F->4	I->2	L->1	O->1	V->1	
ktiv:	 ->2	
ktiv?	F->1	N->1	
ktiva	 ->33	,->2	.->2	r->11	s->1	v->7	
ktive	 ->15	n->8	r->1	t->86	
ktivf	ö->3	
ktivi	s->3	t->37	
ktivt	 ->47	,->2	.->3	
ktkon	c->1	
ktlig	 ->2	a->2	e->14	
ktlin	j->74	
ktlös	.->1	h->2	
ktmed	e->1	l->1	
ktmis	s->1	
ktnin	g->55	
ktobe	r->8	
ktor 	a->2	d->1	f->1	i->2	o->1	s->6	ä->1	
ktor,	 ->5	
ktor.	D->1	J->3	T->1	
ktora	t->18	
ktore	r->33	
ktorh	a->1	
ktori	e->1	s->2	t->4	
ktorn	 ->21	)->1	,->12	.->10	?->1	s->4	
ktorp	o->1	
ktors	 ->1	a->1	i->1	ö->1	
ktpun	k->2	
ktra 	ö->1	
ktric	i->1	
ktron	i->9	
ktrum	 ->1	e->1	
kts a	v->1	
kts e	f->1	l->1	
kts i	 ->1	
kts l	i->1	
kts o	c->1	l->1	
kts u	n->2	p->1	
kts ö	v->1	
kts!F	ö->1	
ktsan	a->3	
ktsba	s->1	
ktsfo	r->1	
ktsfö	r->3	
ktsme	t->1	
ktspl	a->1	
ktspr	o->1	
ktta 	E->1	d->2	
kttag	e->1	
kttar	 ->1	
kttas	 ->3	
ktual	i->1	
ktuel	l->34	
ktum 	a->56	i->1	m->1	o->1	s->1	ä->4	
ktum,	 ->1	
ktum.	V->2	
ktume	t->1	
ktur 	-->1	f->5	g->1	o->2	s->4	u->1	ä->1	
ktur,	 ->4	
ktur.	D->1	F->1	V->1	
kturb	e->1	
kture	l->12	n->10	r->30	
kturf	o->58	
kturm	ä->1	
kturn	ä->1	
kturp	o->11	r->1	
kturr	e->1	
kturs	t->3	
kturu	t->2	
kturå	t->1	
ktyg 	f->3	n->1	o->1	s->1	
ktyg?	D->1	
ktygs	s->1	
ktyr.	E->1	
ktär 	a->2	f->1	o->1	
ktär,	 ->1	
ktär.	R->1	
ktäre	n->2	r->1	
ktör 	i->1	
ktör,	 ->1	
ktöre	n->1	r->19	
ktörs	k->1	
kubik	m->2	
kugga	 ->1	n->1	
kuggb	o->1	
kula 	o->1	
kula.	J->1	
kulat	i->5	
kulda	n->1	
kuldb	e->1	
kulde	n->1	
kuler	a->2	
kulis	s->1	
kull 	b->3	f->2	g->1	h->1	i->2	s->2	v->1	ä->1	
kull,	 ->2	
kull.	D->1	K->1	V->1	
kulle	 ->484	,->2	
kullk	a->1	
kulor	 ->1	
kultu	r->121	
kulär	a->1	
kumen	t->46	
kumul	a->1	e->1	
kund,	 ->1	
kunde	 ->27	r->3	
kundv	a->1	
kundä	r->1	
kunga	r->15	
kunna	 ->208	n->2	r->2	t->43	
kunni	g->6	
kunsk	a->17	
kupan	t->1	
kupat	i->1	
kuper	a->3	
kuppg	i->1	
kur f	ö->1	
kurar	n->1	
kurre	n->280	r->5	
kurs 	i->1	m->2	o->1	
kurs,	 ->1	
kurs.	D->1	
kurse	n->3	r->7	
kursä	n->1	
kus f	ö->1	
kus s	t->1	
kus.D	e->1	
kuser	a->3	
kussi	o->61	
kust 	e->1	
kustb	e->1	
kuste	n->15	r->5	
kustl	i->2	
kustm	y->3	
kusto	m->2	
kustr	e->1	
kustv	a->1	
kuta 	l->1	s->1	
kutab	e->2	l->1	
kutan	,->1	.->1	
kuter	a->78	
kuum 	o->1	
kuumt	a->1	
kuyu 	i->1	s->1	
kva, 	s->1	
kvald	a->2	
kvali	f->15	t->36	
kvant	i->7	
kvar 	d->1	e->4	f->2	i->4	m->1	p->5	r->1	s->1	
kvar,	 ->2	
kvar.	D->1	J->1	
kvar;	 ->1	
kvarh	ä->1	å->2	
kvars	t->8	
kvat 	b->1	f->1	r->1	
kvata	 ->2	
kvati	o->1	
kvens	 ->4	.->1	e->41	
kvent	 ->9	,->2	a->4	e->1	
kvest	o->3	
kvick	s->3	
kvidd	 ->2	.->1	
kvinn	a->1	l->2	o->56	
kvist	 ->1	
kvot 	p->1	s->1	v->1	ä->1	
kvot!	D->1	
kvot,	 ->1	
kvote	n->3	r->7	
kväl 	h->1	i->1	m->1	u->1	
kväll	 ->2	,->2	.->2	?->1	a->1	e->2	
kväml	i->15	
kvämt	 ->1	
kvärd	 ->1	a->2	e->3	i->5	
kvärt	 ->6	,->1	
kväva	 ->2	
kvård	 ->1	)->1	s->1	
ky fö	r->1	
kydd 	a->4	b->1	e->1	f->13	i->2	m->3	o->3	s->4	v->2	ö->1	
kydd)	,->1	
kydd,	 ->3	
kydd.	D->2	J->1	N->1	R->1	V->1	
kydda	 ->24	d->2	n->1	r->2	s->2	
kydde	t->18	
kydds	m->4	n->6	o->2	p->1	s->2	t->1	
kyfal	l->1	
kyhög	a->1	
kyla.	H->1	
kylan	 ->1	
kyldi	g->29	
kylig	a->1	
kylla	 ->2	s->1	
kylle	r->1	
kylls	 ->1	
kymme	r->6	
kymra	d->7	r->2	t->1	
kymts	 ->1	
kynda	 ->5	n->1	r->2	s->3	
kynds	a->4	
kyrko	g->1	
kyvär	d->1	
käl -	 ->2	
käl 6	,->1	
käl a	t->2	
käl b	i->1	
käl d	å->1	
käl e	f->1	
käl f	ö->4	
käl h	a->2	ä->1	
käl i	n->4	
käl n	i->1	
käl o	c->2	
käl s	k->1	o->5	
käl t	i->5	
käl ä	r->2	
käl, 	k->1	
käl.A	l->1	
käl.D	e->1	
käl.F	ö->1	
käl.J	a->1	
kälen	 ->3	
kälet	 ->8	,->1	
kälig	 ->1	
källa	 ->6	.->1	r->1	
källo	r->39	
kämda	 ->1	
kämma	s->2	
kämne	n->1	
kämpa	 ->27	n->1	r->4	t->2	
kämpn	i->12	
kämts	a->1	
känd 	(->1	m->4	
känd,	 ->2	
känd.	K->1	
kända	 ->9	.->3	
kände	 ->14	,->1	s->5	
känka	 ->2	
känna	 ->27	,->1	.->2	g->9	n->23	s->7	
känne	d->1	l->1	r->70	t->6	
känns	 ->3	.->1	
känsl	a->15	i->21	o->7	
känt 	-->1	a->3	d->2	e->3	f->1	m->1	o->1	s->4	t->1	u->2	
känt,	 ->2	
känts	 ->8	
kär n	e->1	
kär p	o->1	
kära 	b->1	k->47	l->2	o->2	p->1	
käre 	k->1	
kärl 	o->1	
kärle	k->2	
kärna	n->4	
kärne	n->8	
kärnf	r->2	
kärni	n->3	
kärnk	a->1	r->20	
kärnp	r->2	u->2	
kärns	t->1	ä->3	
kärnt	e->2	
kärnv	a->8	
kärpa	 ->6	s->2	
kärpn	i->1	
kärpt	a->2	
kärs 	n->1	
kådad	 ->1	e->1	
kådar	e->1	
kådli	g->6	
kådni	n->1	
kålen	 ->1	
kår, 	s->1	
kåt i	 ->2	
kåtst	r->1	
köksb	o->1	
köl n	ä->1	
köl, 	s->1	
kölar	.->1	
köldb	e->1	
köldg	r->1	
könen	 ->3	
könhe	t->1	
könsg	r->1	
könsk	a->5	
köp a	v->2	
köpar	e->3	n->1	
köper	 ->1	
köpkr	a->1	
köpsb	e->1	
köpsl	a->1	
köpt 	i->1	
kör ö	v->1	
kör.K	o->1	
köra 	d->1	f->1	m->1	
köras	 ->1	
körd 	a->1	
körda	t->1	
körde	n->1	
körni	n->2	
körs 	i->2	
körsp	o->1	
kört 	e->1	f->1	i->1	
köt 9	3->1	
köt l	o->1	
köta 	E->1	d->1	m->1	s->3	
kötas	 ->1	
köter	 ->1	
köts 	b->1	i->1	
köts.	V->1	
kötse	l->5	
kött 	o->1	s->2	t->1	v->1	
kötte	 ->2	
köttk	r->1	
kötts	 ->1	-->1	p->1	
kövla	d->1	
köy -	 ->1	
l "Mi	s->1	
l (Br	y->1	
l (ko	d->2	
l - d	e->2	å->1	
l - f	ö->1	
l - n	a->1	å->1	
l - o	m->1	
l - r	i->1	
l - s	o->1	ö->1	
l - u	t->2	
l - ö	v->1	
l -, 	d->1	
l 1 i	 ->1	
l 1 o	c->2	
l 1 u	r->1	
l 1, 	2->1	a->1	
l 1-o	m->4	
l 1-r	e->5	
l 1-s	t->2	
l 1.J	a->1	
l 10 	0->1	
l 105	 ->1	
l 110	 ->1	
l 12 	o->1	
l 12,	 ->1	
l 13 	(->1	A->1	i->2	
l 13.	F->1	
l 143	 ->1	
l 15 	p->1	
l 158	 ->1	)->1	.->1	
l 16)	 ->1	
l 193	 ->1	
l 195	 ->1	
l 199	9->2	
l 2 -	 ->1	
l 2 0	0->1	
l 2 b	l->1	
l 2 e	l->1	
l 2 o	c->1	
l 2 s	o->1	
l 2, 	i->1	
l 2,4	8->1	
l 2,6	 ->1	
l 2-o	m->2	
l 2-s	t->1	
l 2.1	 ->1	
l 2.2	 ->1	
l 2.M	e->1	
l 226	 ->1	
l 25 	t->1	
l 255	 ->4	
l 280	 ->4	.->1	
l 299	.->2	
l 3 0	0->1	
l 3.1	)->1	
l 3.8	 ->1	
l 30 	i->1	m->1	
l 33 	f->1	i->1	
l 37 	i->1	
l 37.	2->1	
l 39 	i->1	
l 4 c	 ->1	
l 4 i	 ->4	
l 4 p	r->1	
l 4.2	)->1	
l 42 	i->1	
l 48 	i->2	
l 5 g	ä->1	
l 5.4	 ->1	
l 50 	i->1	m->1	
l 50,	 ->1	
l 52 	i->1	
l 56,	 ->1	
l 5b 	k->1	
l 5b.	D->1	
l 6 i	 ->6	
l 6 o	c->3	
l 6, 	t->1	
l 6.S	å->1	
l 62 	i->1	
l 67 	i->1	
l 7 i	 ->6	
l 7 n	ä->1	
l 7, 	s->1	
l 7,4	2->1	
l 700	 ->1	
l 75 	-->1	
l 77 	m->1	
l 81 	o->1	
l 81.	1->4	3->5	
l 82,	 ->1	
l 82.	I->1	
l 83 	p->1	
l 85 	p->1	
l 87.	1->1	2->1	
l 88 	i->1	ä->1	
l 9 m	i->1	
l 9.1	 ->1	
l 91 	p->1	
l 94 	n->1	p->1	
l 94,	 ->1	
l 95 	i->1	
l Alb	r->1	
l Bar	n->1	
l Bas	k->1	
l Bou	r->2	
l Bry	s->2	
l Chi	q->1	
l Con	a->1	
l Cou	n->1	
l Den	 ->1	
l Dim	i->1	
l EG 	t->1	
l EG-	k->1	r->1	
l EU 	"->1	o->1	
l EU-	k->1	
l EU.	N->1	
l EU:	s->2	
l Eft	a->1	
l Eur	o->25	
l Fra	n->3	
l För	e->4	
l Gen	e->1	
l Gre	k->1	
l Hei	n->1	
l Hil	t->1	
l Int	e->2	
l Irl	a->1	
l Kan	 ->1	
l Kar	a->1	
l Kau	f->1	
l Kin	a->1	
l Kir	g->2	
l Kos	o->9	
l Kou	c->1	
l Kul	t->1	
l Lor	d->2	
l McN	a->1	
l Mic	h->1	
l Mor	a->1	g->1	
l Nie	l->2	
l Nya	 ->1	
l OLF	A->1	
l PPE	-->1	
l Pal	e->1	
l Pat	t->2	
l Pea	k->1	
l Pol	l->1	
l Pur	v->1	
l Rap	k->1	
l Rio	f->1	
l Sch	ü->1	
l She	l->1	
l Sol	a->2	b->1	
l St.	V->1	
l Str	a->1	
l Syr	i->1	
l The	a->1	
l Tib	e->1	
l Tre	d->1	
l Tys	k->2	
l Uls	t->1	
l Ver	h->1	
l Wal	l->1	
l Was	h->1	
l Wil	h->1	
l Wur	t->1	
l abs	o->1	
l acc	e->1	
l age	r->1	
l ald	r->2	
l all	a->20	e->1	m->6	s->1	t->7	
l and	e->1	r->4	
l anf	ö->1	
l ang	å->1	
l anl	e->1	
l anm	ä->2	
l ann	a->1	
l anp	a->1	
l ans	e->1	j->1	l->1	v->7	ö->2	
l ant	a->3	
l anv	ä->11	
l app	e->1	
l arb	e->8	
l arm	o->1	
l art	 ->1	i->4	
l att	 ->300	
l av 	E->7	F->2	I->1	J->1	K->1	O->1	a->9	b->4	d->44	e->7	f->6	g->3	h->1	i->2	k->7	l->3	m->5	n->1	o->2	p->4	r->3	s->5	t->4	u->2	v->4	ä->1	å->1	ö->1	
l av,	 ->1	
l avg	ö->2	
l avk	r->1	
l avl	ä->1	
l avm	a->1	
l avs	e->1	k->1	l->7	
l avt	a->2	
l avv	e->1	i->1	ä->1	
l bac	k->1	
l bag	a->1	
l bal	a->1	
l ban	k->1	t->1	
l bar	a->11	
l bas	e->1	
l be 	P->1	e->1	h->1	k->2	s->1	
l bed	r->1	ö->4	
l bef	i->1	o->2	ä->1	
l beg	r->6	ä->1	
l beh	a->3	o->2	å->2	ö->3	
l bek	ä->1	
l bem	ö->1	
l ber	 ->1	e->2	ä->1	ö->1	
l bes	l->9	t->4	
l bet	a->17	e->1	o->5	r->4	y->6	ä->4	
l bev	a->2	i->3	
l bib	e->3	
l bid	r->5	
l bil	 ->1	a->1	d->1	l->1	p->1	
l bla	n->1	
l bli	 ->21	r->2	
l blo	m->2	
l bor	d->2	t->1	
l bot	t->3	
l bra	 ->1	
l bri	s->2	
l bro	t->1	
l brä	n->1	
l brö	s->1	
l bud	g->1	
l byg	g->2	
l bär	a->3	
l bäs	t->1	
l bät	t->2	
l båd	a->2	
l böd	e->1	
l bör	 ->3	j->10	
l ca 	3->1	
l cen	t->1	
l cit	e->2	
l cor	r->1	
l dag	s->1	
l de 	a->3	b->4	d->1	e->3	f->9	g->3	h->3	i->2	k->3	l->1	m->7	n->6	o->5	p->5	r->1	s->9	t->2	u->1	v->2	ä->1	
l deb	a->4	
l dec	e->1	
l def	i->1	
l del	 ->6	.->3	a->3	e->1	t->2	
l dem	 ->6	,->2	.->1	o->2	
l den	 ->68	,->1	.->1	n->20	
l der	a->5	
l des	 ->1	s->12	
l det	 ->45	,->5	.->6	?->1	t->31	
l dia	l->3	
l dir	e->17	
l dis	c->2	k->6	
l doc	k->2	
l dom	s->2	
l dra	 ->1	r->1	
l dri	v->1	
l dry	f->1	
l dum	h->1	p->2	
l där	 ->3	e->1	f->13	
l då 	a->1	d->1	u->1	
l då?	I->1	
l eff	e->2	
l eft	e->4	
l ege	n->3	
l eko	n->3	
l ell	e->7	
l eme	l->2	
l emi	g->1	
l en 	"->2	a->9	b->7	c->3	d->3	e->8	f->4	g->7	h->5	i->5	k->5	l->2	m->2	n->1	o->5	p->4	r->4	s->18	t->2	u->1	v->5	ä->1	ö->5	
l enb	a->1	
l end	a->3	
l ene	r->2	
l enk	e->1	
l enl	i->1	
l ent	r->1	
l er 	a->1	b->1	s->1	
l er,	 ->4	
l er:	 ->1	
l erb	j->1	
l erf	o->1	
l erh	å->1	
l eri	n->2	
l ers	ä->1	
l ert	 ->1	
l ett	 ->32	
l eur	o->3	
l exe	m->45	
l exi	s->1	
l fal	l->3	
l fam	i->1	
l far	t->1	
l fas	c->1	t->1	
l fat	t->7	
l feb	r->1	
l fel	a->2	
l fic	k->1	
l fin	a->2	n->4	
l fis	k->1	
l fle	r->1	
l fly	k->1	t->1	
l fon	d->3	
l for	d->1	m->2	t->7	
l fra	m->10	
l fre	d->2	
l fri	 ->2	g->1	h->1	
l fru	 ->1	
l frä	m->8	
l frå	g->16	n->15	
l ful	l->5	
l fun	g->9	
l fyl	l->2	
l fär	g->1	
l fäs	t->1	
l få 	d->1	e->3	f->1	g->1	k->1	u->1	v->1	ö->1	
l fån	g->1	
l får	 ->2	
l föl	j->24	
l för	 ->76	a->2	b->7	d->8	e->25	f->6	h->4	i->1	k->4	l->7	m->11	o->8	s->26	t->5	v->3	ä->5	
l gag	n->3	
l gam	l->1	m->1	
l gan	s->1	
l gar	a->2	
l ge 	a->1	d->1	e->2	i->1	k->1	m->1	n->1	r->1	u->1	
l gem	e->8	
l gen	e->1	o->16	
l ges	 ->1	t->1	
l get	t->1	
l gis	s->1	
l glä	d->1	
l god	 ->2	a->1	k->4	o->3	
l gra	n->1	t->7	
l gru	n->12	p->1	
l gäl	l->8	
l gär	n->7	
l gå 	a->1	f->1	i->1	s->1	t->3	u->1	v->1	å->1	
l gå.	V->1	
l gån	g->2	
l gör	 ->2	a->22	s->1	
l ha 	a->2	d->1	e->20	g->2	h->1	i->1	k->3	m->3	n->1	s->1	t->4	
l ha.	A->1	
l ham	n->1	
l han	d->10	s->6	t->6	
l har	 ->16	m->1	
l hav	e->1	s->13	
l hed	e->1	
l hel	a->2	t->2	
l hem	l->2	
l hen	n->1	
l her	r->4	
l hin	d->4	n->1	
l hjä	l->6	
l hon	o->1	
l hop	p->1	
l hum	a->1	
l hur	 ->5	
l hyc	k->1	
l häl	s->1	
l hän	d->1	s->2	
l här	 ->4	m->1	
l hål	l->2	
l hög	e->1	r->1	s->2	
l hör	a->3	
l i 1	5->1	
l i A	m->1	
l i D	a->1	
l i E	u->4	
l i F	r->1	
l i M	o->1	
l i V	e->1	
l i a	l->2	n->2	r->2	
l i d	a->2	e->14	
l i e	f->1	n->1	
l i f	o->1	r->5	ö->2	
l i g	e->3	
l i i	n->1	
l i k	e->1	
l i l	a->1	i->1	
l i m	e->1	i->2	o->1	å->1	
l i n	a->1	
l i o	k->1	r->1	
l i p	a->1	
l i s	i->6	t->1	y->1	ä->1	
l i t	a->1	
l i u	t->2	
l i v	a->1	i->3	ä->1	å->2	
l i ä	n->1	
l ick	e->1	
l idé	n->1	
l in 	i->1	
l inb	e->1	l->1	
l ind	i->2	u->3	
l inf	o->3	ö->4	
l ing	e->1	å->3	
l inl	e->5	
l inn	e->3	
l ino	m->9	
l inr	i->1	ä->4	
l ins	e->1	i->1	k->1	t->3	y->1	
l int	a->2	e->56	r->2	
l inv	a->1	
l inö	v->1	
l isr	a->1	
l jag	 ->106	,->2	
l jan	u->1	
l jor	d->1	
l ju 	a->1	d->1	i->1	s->1	
l jul	i->1	
l jus	t->1	
l jäm	s->2	
l kal	l->1	
l kam	m->2	p->1	
l kan	 ->13	
l kas	t->1	
l kat	a->1	
l kla	r->4	
l kny	t->1	
l kod	e->1	
l kol	l->5	
l kom	m->55	p->1	
l kon	c->2	f->1	k->7	s->3	t->7	v->2	
l kor	r->1	t->2	
l kos	t->1	
l kra	v->1	
l kri	m->1	s->1	t->1	
l krä	v->2	
l kul	t->1	
l kun	n->57	
l kve	s->1	
l kvi	n->4	
l kvä	l->1	
l kän	n->1	
l kär	n->2	
l kök	s->1	
l lag	f->1	
l lan	d->2	
l led	a->5	
l let	t->1	
l lig	g->7	
l lik	a->2	
l liv	 ->1	.->1	e->1	s->2	
l luc	k->1	
l lyc	k->3	
l lyd	a->1	
l lyf	t->1	
l lys	s->2	
l läg	g->4	
l läm	n->5	p->1	
l län	d->2	
l lär	a->1	
l läs	b->1	
l lät	t->2	
l låt	a->3	
l löp	t->1	
l lös	a->1	n->1	
l maj	o->2	
l mak	t->5	
l man	 ->11	
l mar	k->5	
l med	 ->25	b->3	d->2	e->1	l->11	v->4	
l mel	l->10	
l men	 ->2	
l mer	 ->4	
l met	a->1	
l mid	d->1	
l mig	 ->2	,->1	
l mil	j->1	
l min	 ->5	a->2	d->3	i->5	n->1	s->1	u->1	
l mis	s->1	
l mit	t->2	
l mob	i->1	
l mot	 ->2	i->2	s->1	v->1	
l mus	i->1	
l myc	k->5	
l myn	d->3	
l män	 ->1	
l mär	k->1	
l mål	 ->3	
l mån	a->2	g->4	
l mås	t->7	
l möj	l->4	
l möt	e->2	
l nac	k->4	
l nat	i->4	u->6	
l ni 	f->1	g->1	n->2	v->1	
l niv	å->11	
l nog	g->1	
l nor	m->1	
l nu 	g->1	h->1	l->1	t->1	
l ny 	g->1	l->1	
l nya	 ->4	
l nyl	i->1	
l nyt	t->6	
l näm	n->4	
l när	 ->9	m->1	
l näs	t->4	
l nå 	h->1	
l någ	o->10	r->1	
l nöd	v->2	
l oac	c->1	
l och	 ->127	
l ock	s->27	
l oen	i->1	
l off	e->2	
l ofö	r->1	
l oig	e->1	
l ojä	m->1	
l oli	k->3	
l oly	c->2	m->1	
l om 	J->1	a->11	b->1	d->8	f->1	g->1	h->2	k->1	m->1	t->1	u->1	v->1	
l om,	 ->1	
l omf	a->9	
l oml	o->1	
l omr	å->2	ö->2	
l oms	t->1	ä->1	
l omv	a->1	ä->1	
l opt	i->1	
l ord	f->3	
l org	a->2	
l oro	 ->1	,->1	.->1	
l orä	t->1	
l oss	 ->2	,->2	
l oän	d->2	
l par	l->10	
l pas	s->1	
l pel	a->1	
l pen	g->1	s->3	
l per	i->1	s->5	
l pil	o->1	
l pla	n->3	s->1	t->1	
l pol	i->6	
l pos	i->2	
l pra	k->1	
l pre	c->1	m->1	s->5	
l pri	n->1	s->1	v->5	
l pro	b->1	c->2	d->1	g->2	j->2	t->1	
l pun	k->2	
l på 	-->1	a->6	b->1	d->10	e->3	f->2	g->1	h->2	i->1	k->1	m->1	n->1	s->1	v->2	å->1	ö->1	
l på,	 ->1	
l på.	B->1	
l pål	ä->1	
l påm	i->1	
l påp	e->3	
l pås	k->1	t->1	
l påt	v->1	
l påv	e->1	
l rad	 ->1	
l ram	.->1	a->1	
l rat	i->1	
l red	a->3	l->1	o->2	
l ref	o->1	
l reg	e->7	i->5	l->2	
l rek	o->4	
l rep	a->1	
l res	o->2	p->5	u->4	
l ret	r->1	
l rev	i->1	o->1	
l rik	e->1	t->4	
l ris	k->2	
l rol	l->4	
l rym	m->1	
l räc	k->4	
l räk	e->1	
l rät	t->18	
l råd	e->20	
l rör	a->2	l->1	
l rös	t->1	
l sak	e->3	n->1	
l sam	a->1	e->1	m->13	t->3	v->1	
l san	n->1	
l sat	s->1	
l se 	d->2	e->1	f->1	i->1	k->1	p->1	t->5	u->2	v->1	
l ser	v->1	
l ses	 ->2	
l set	t->1	
l sig	 ->3	n->1	
l sim	u->1	
l sin	 ->7	a->7	
l sis	t->12	
l sit	t->6	u->3	
l sjä	l->3	
l sjö	s->4	
l ska	f->1	l->6	p->9	t->1	
l ske	 ->3	p->1	
l ski	l->5	
l skj	u->2	
l sko	g->3	
l skr	o->1	
l sku	l->6	
l sky	d->6	l->1	
l skö	t->2	
l slu	t->15	
l slå	 ->2	
l små	 ->2	
l sna	b->1	
l soc	i->4	
l sol	i->3	
l som	 ->105	
l spe	c->1	l->2	
l spä	n->1	
l sta	d->2	n->2	r->2	t->3	
l ste	e->1	
l sti	m->1	
l sto	r->13	
l str	a->1	u->4	y->1	
l sty	r->1	
l stä	l->3	r->2	
l stå	 ->6	l->19	n->17	
l stö	d->2	t->1	
l sub	s->3	v->1	
l sus	p->1	
l suv	e->1	
l sva	g->1	r->2	
l svå	r->1	
l syn	e->1	v->1	
l sys	s->5	
l säg	a->38	s->1	
l säk	e->9	r->1	
l sän	d->1	k->1	
l sär	s->4	
l sät	t->2	
l så 	a->2	l->1	s->1	
l såd	a->2	
l sör	j->1	
l ta 	d->2	h->5	i->2	s->1	u->6	ö->1	
l tac	k->21	
l tal	a->8	e->2	m->1	s->1	
l tas	 ->3	
l ten	d->1	
l ter	r->1	
l tex	t->1	
l tid	e->1	i->2	
l til	l->40	
l tit	t->2	
l tol	k->2	
l tot	a->1	
l tra	n->2	
l tre	 ->2	d->2	
l tro	 ->2	t->1	v->2	
l try	g->3	
l trä	d->3	f->1	
l tur	i->1	
l tvi	n->1	
l tvä	r->1	
l två	 ->5	n->1	
l tyc	k->2	
l tyd	l->1	
l täc	k->1	
l tän	k->1	
l u-l	ä->1	
l und	a->2	e->13	v->1	
l uni	o->3	
l upp	d->1	e->1	f->3	h->2	m->4	n->7	r->4	s->2	
l ur 	j->1	k->1	p->1	s->1	
l urs	p->1	
l urv	a->1	
l uta	n->8	r->1	
l utb	r->1	y->1	
l utf	o->5	ö->2	
l utg	ö->3	
l utn	y->1	
l uto	m->1	
l utr	o->2	
l uts	k->3	l->8	ä->1	
l utt	a->4	r->4	
l utv	e->6	i->4	
l utö	v->2	
l vad	 ->10	
l val	.->1	
l van	 ->1	
l vap	e->1	
l var	 ->2	a->33	f->7	j->3	k->1	m->1	
l ver	k->15	
l vet	 ->2	,->1	a->5	e->1	
l vi 	a->6	b->2	d->1	f->3	g->1	h->3	i->7	l->1	m->2	n->3	o->2	r->2	s->4	v->2	ä->1	
l via	 ->1	
l vic	e->1	
l vid	 ->4	a->3	t->3	
l vik	t->1	
l vil	k->6	l->1	
l vis	a->4	s->7	
l vol	y->1	
l von	 ->3	
l vor	e->2	
l väg	s->1	
l väl	d->1	k->1	
l vän	d->1	s->1	
l vär	n->1	
l väs	e->1	
l vår	 ->6	a->5	t->5	
l yrk	e->2	
l ytt	r->3	
l Öst	e->1	
l ägn	a->1	
l än 	a->1	e->6	k->1	
l änd	a->1	r->9	å->5	
l är 	"->1	a->8	d->3	e->5	f->3	g->1	i->3	j->2	k->1	l->1	o->2	r->1	s->1	u->2	v->5	ö->1	
l är?	H->1	
l äve	n->6	
l åkl	a->2	
l år 	2->1	o->1	
l åsi	k->1	
l åst	a->2	
l åt 	a->1	
l åta	l->2	
l åte	r->14	
l åtg	ä->3	
l åts	t->1	
l ått	a->1	
l öka	 ->3	.->1	s->1	
l ökn	i->1	
l öns	k->1	
l öpp	e->3	
l öst	e->1	
l öve	r->20	
l! In	g->1	
l! Ja	g->1	
l!Her	r->1	
l!Här	 ->1	
l!Jag	 ->1	
l!Men	 ->1	
l!Til	l->1	
l" me	d->1	
l" oc	h->1	
l", s	o->1	
l", v	i->1	
l".I 	n->1	
l'eau	 ->1	
l, An	v->1	
l, Re	d->1	
l, Ty	s->1	
l, an	g->1	
l, at	t->5	
l, av	 ->1	s->1	
l, be	v->1	
l, de	 ->2	n->1	t->1	
l, di	s->1	
l, dv	s->1	
l, dä	r->2	
l, då	 ->1	
l, ef	t->3	
l, el	l->2	
l, er	k->1	
l, et	t->2	
l, eu	r->1	
l, fo	r->1	
l, fr	a->2	
l, fö	r->5	
l, ge	n->1	
l, gr	u->1	
l, ha	n->1	r->3	
l, hu	r->1	
l, hä	v->1	
l, i 	a->1	h->1	k->1	l->1	s->2	v->1	
l, in	t->1	
l, ja	g->1	
l, ju	 ->1	s->1	
l, ka	n->1	
l, ko	m->1	n->2	
l, ku	n->1	
l, la	n->1	
l, li	k->1	
l, lä	k->1	
l, me	d->4	n->15	
l, mo	t->1	
l, na	t->1	
l, ni	 ->1	
l, nä	m->2	r->3	
l, nå	g->2	
l, oc	h->30	
l, om	 ->2	
l, po	l->1	
l, pr	o->1	
l, på	 ->1	
l, re	s->1	
l, rä	k->1	
l, rö	r->1	
l, si	n->1	
l, so	m->15	
l, så	 ->5	v->1	
l, sö	n->1	
l, ti	l->1	
l, to	b->1	n->1	
l, tå	g->1	
l, un	i->1	
l, ut	a->4	
l, va	r->3	t->1	
l, vi	 ->2	d->2	l->2	s->1	
l, än	 ->1	
l, äv	e->3	
l, ån	y->1	
l, åt	e->2	
l, öv	e->1	
l- oc	h->18	
l-2-o	m->1	
l-Del	g->1	
l-Fin	a->3	
l-Hei	n->1	
l-I);	 ->1	
l-II)	 ->1	
l-Rob	l->1	
l-Sha	r->1	
l-She	i->5	
l-Syr	i->1	
l-för	d->1	
l-pro	g->1	
l-soc	i->2	
l. 11	.->6	
l. 12	.->6	
l. 13	.->1	
l. 15	.->2	
l. 17	.->1	
l. 19	.->1	
l. 20	.->1	
l. 21	.->2	
l. De	t->1	
l. En	 ->1	
l. Ja	g->1	
l. oc	h->1	
l.12.	0->1	
l.All	m->1	
l.Ang	å->1	
l.Avs	l->1	
l.Bet	ä->1	
l.Bil	t->1	
l.Bäs	t->1	
l.De 	n->1	s->1	
l.Den	 ->7	
l.Des	s->1	
l.Det	 ->23	t->11	
l.Där	 ->1	f->2	
l.EU-	k->1	
l.Eft	e->1	
l.Enl	i->3	
l.Ett	 ->3	
l.Eur	o->2	
l.Fin	a->2	
l.Fra	n->1	
l.Fru	 ->3	
l.Frå	g->1	
l.För	 ->8	
l.Gen	o->1	
l.Har	 ->1	
l.Her	r->8	
l.Hur	 ->1	
l.Här	 ->1	
l.I A	m->1	
l.I d	e->1	
l.I e	n->1	
l.I f	l->1	ö->1	
l.I o	c->1	
l.I s	j->1	
l.I u	p->1	
l.Ing	e->1	
l.Int	e->1	
l.Ja 	e->1	
l.Jag	 ->21	
l.Kan	 ->1	
l.Kom	m->3	
l.Kos	t->1	
l.Kul	t->1	
l.Kär	a->1	
l.Lyn	n->1	
l.Mar	k->1	
l.Med	 ->1	
l.Men	 ->8	
l.Min	 ->1	
l.Mål	e->1	
l.När	 ->4	
l.Om 	v->1	
l.Ork	a->1	
l.Per	s->1	
l.Pro	d->1	
l.På 	d->1	
l.Res	u->1	
l.Sam	m->2	t->1	
l.San	n->1	
l.Sch	ü->1	
l.Sjä	l->1	
l.Små	 ->1	
l.Som	 ->1	
l.Str	ä->1	
l.Så 	e->1	t->1	v->1	
l.Sås	o->1	
l.Tan	k->1	
l.Tro	r->1	
l.Två	 ->1	
l.Tän	k->1	
l.Utm	a->1	
l.Vi 	a->1	d->1	h->3	k->3	m->4	s->4	t->1	v->3	ä->3	
l.Von	 ->1	
l.Vår	a->1	
l.a. 	a->2	b->1	d->1	e->2	f->5	g->2	i->2	m->1	n->3	o->2	p->1	s->3	u->1	v->1	
l.Än 	e->1	
l.Änd	r->1	
l.Är 	d->1	
l.Äve	n->1	
l: "h	e->1	
l: Eu	r->1	
l: Fi	r->1	
l: Os	l->1	
l: Un	d->1	
l: Ve	m->1	
l: Vi	 ->1	
l: at	t->1	
l: de	t->1	
l: en	 ->1	
l: ja	g->1	
l: pr	o->1	
l; at	t->1	
l; fö	r->1	
l; i 	e->1	
l?. (	E->1	
l?Dag	e->1	
l?Ell	e->1	
l?Hur	 ->1	
l?Jag	 ->2	
l?Kol	l->1	
lFina	 ->1	
la - 	i->1	s->1	
la 90	-->1	
la Al	e->1	
la Ba	l->1	
la EU	-->2	:->2	
la Eu	r->20	
la Fö	r->1	
la Hi	c->1	
la Ko	s->1	u->1	
la Lo	i->1	
la Me	l->1	
la Pa	k->1	
la Su	a->1	
la UC	K->1	
la ag	e->1	
la ak	t->3	
la al	l->5	
la an	d->7	f->1	o->1	s->7	
la ar	b->4	v->1	
la as	p->8	y->1	
la at	o->2	t->30	
la av	 ->6	,->1	d->1	s->4	t->3	v->1	
la ba	k->2	r->1	
la be	f->1	g->1	h->3	k->2	l->2	r->1	s->16	t->4	
la bi	d->4	l->10	
la bl	a->1	i->1	
la bo	l->3	r->1	
la br	o->1	ä->2	
la bu	d->2	
la bö	r->3	
la de	 ->51	l->2	m->22	n->25	s->19	t->14	
la di	a->5	g->1	m->5	p->1	r->3	s->2	
la do	k->1	m->5	
la dr	a->1	
la dö	d->1	
la ef	t->2	
la eg	n->1	o->1	
la ek	o->7	
la el	e->2	l->8	
la em	o->2	
la en	 ->30	d->1	e->4	h->1	s->1	
la er	 ->1	,->1	a->4	f->2	k->1	
la et	t->8	
la eu	r->7	
la ev	e->2	
la ex	e->1	
la fa	k->1	l->8	m->1	r->11	s->5	
la fi	l->1	n->3	
la fl	e->1	o->1	
la fo	l->2	n->2	r->13	
la fr	a->3	i->3	o->1	å->26	
la fu	n->1	
la få	 ->1	r->1	
la fö	l->2	r->41	
la ge	m->5	n->1	
la gi	l->1	v->1	
la gl	ä->1	
la go	d->3	
la gr	a->1	u->10	ä->2	
la gå	r->1	
la ha	 ->1	d->1	m->2	n->7	r->6	t->1	v->1	
la he	l->1	
la hi	n->2	
la hj	ä->2	
la ho	n->1	p->3	s->1	
la hu	r->2	v->1	
la hä	n->1	
la hå	l->1	
la hö	g->5	
la i 	E->1	d->1	e->1	f->1	g->1	i->1	m->1	o->1	p->1	t->1	
la id	e->3	é->2	
la ig	e->1	
la in	 ->4	,->1	b->1	d->2	f->1	i->4	l->1	n->1	o->2	r->1	s->13	t->6	v->4	
la is	ä->1	
la jo	r->3	
la ju	r->2	
la jä	m->2	
la ka	m->3	n->3	t->3	
la kl	a->2	i->2	y->1	
la kn	o->1	y->1	
la ko	l->1	m->13	n->24	r->2	s->7	
la kr	a->6	
la kv	a->3	
la kä	n->1	
la kö	l->1	
la la	g->4	n->1	r->1	
la le	d->5	
la li	k->2	n->1	v->4	
la lo	k->1	
la lä	m->1	n->6	
la lö	f->1	s->3	
la ma	j->1	k->1	n->1	r->7	x->1	
la me	d->37	n->1	r->2	
la mi	g->5	n->3	s->2	t->6	
la mo	d->2	t->2	
la mu	r->1	
la my	c->1	n->31	
la mä	n->3	
la må	s->4	
la mö	j->4	t->1	
la na	t->1	
la ne	o->1	r->1	
la ni	m->1	v->8	
la no	r->1	t->1	
la nu	v->1	
la ny	a->3	
la nä	r->1	t->3	
la nå	g->1	
la nö	d->1	
la ob	a->3	
la oc	h->61	
la od	d->1	
la of	e->1	
la oj	ä->1	
la ol	i->3	j->2	
la om	 ->46	.->3	b->2	r->13	s->7	v->1	
la op	a->1	e->2	
la or	g->5	i->1	s->1	
la os	s->5	
la pa	r->24	
la pe	n->1	r->2	
la pl	a->1	ä->1	
la po	l->15	
la pr	e->2	i->6	o->15	
la pu	n->1	
la på	 ->6	p->1	
la ra	d->1	m->2	p->1	
la re	f->2	g->26	k->1	l->1	n->1	s->4	
la ri	k->1	s->2	
la ro	,->1	
la ru	t->1	
la rä	d->1	t->15	
la rö	r->3	
la sa	k->1	m->23	
la se	k->3	
la si	d->2	g->15	n->18	t->7	
la sj	ä->1	ö->4	
la sk	a->10	e->1	i->8	o->1	r->2	u->1	y->2	ä->2	
la sl	a->3	u->1	
la sn	e->1	
la so	c->2	m->15	
la sp	e->5	ö->1	
la st	a->4	o->2	r->6	y->1	ä->2	ö->14	
la su	b->1	m->1	
la sv	å->1	
la sy	f->1	n->1	s->6	
la sä	g->1	k->1	t->3	
la så	 ->2	d->2	
la ta	 ->1	l->2	
la te	r->1	x->2	
la ti	d->11	l->9	
la tj	ä->11	
la to	l->2	n->1	
la tr	a->6	e->1	o->1	y->2	
la ty	n->1	p->1	
la tä	v->1	
la un	d->4	i->7	
la up	p->11	
la ur	h->1	
la ut	 ->2	b->3	g->3	k->1	l->1	s->5	t->2	v->14	
la va	l->1	p->1	r->4	
la ve	r->5	t->5	
la vi	d->1	k->3	l->4	n->1	s->4	
la vä	d->1	g->1	r->7	s->1	v->1	
la vå	r->10	
la än	d->4	
la är	 ->4	.->1	
la å 	m->1	
la åk	l->2	
la år	e->1	l->1	
la ås	i->1	
la åt	e->4	g->6	
la ön	s->1	
la öp	p->1	
la ös	t->1	
la öv	e->4	r->1	
la!He	r->1	
la" s	o->1	
la" v	a->1	
la".B	a->1	
la".H	i->1	
la"; 	ö->1	
la, a	t->1	
la, c	o->1	
la, d	e->1	
la, f	ö->1	
la, h	a->1	ö->1	
la, i	n->2	
la, k	a->1	
la, l	å->1	
la, m	o->1	
la, n	e->1	ä->1	
la, o	c->3	
la, p	å->1	
la, r	a->1	e->1	
la, s	o->2	t->1	
la, v	i->1	
la, ä	v->1	
la.Bi	l->1	
la.De	 ->1	s->2	t->8	
la.Dä	r->1	
la.He	l->1	r->1	
la.I 	d->1	
la.Ja	g->3	
la.Ko	m->1	
la.Me	n->2	
la.Nä	r->1	
la.Sm	å->1	
la.Vi	 ->4	
la.Öv	e->1	
la:Fö	r->1	
la?Av	s->1	
la?De	 ->1	n->1	t->1	
laams	 ->1	
labor	a->3	
lacer	a->15	i->2	
lacio	 ->7	,->3	.->2	:->1	s->2	
lad a	t->12	
lad e	l->1	
lad f	ö->2	
lad h	ä->1	
lad i	n->1	
lad l	e->1	
lad m	a->1	e->1	
lad o	c->1	
lad p	e->1	
lad r	e->2	
lad s	o->1	t->1	
lad ö	v->4	
lad, 	m->1	
lada 	o->1	ö->2	
ladak	i->1	
ladda	d->1	
ladde	 ->2	
lade 	1->1	4->1	V->1	a->6	d->6	e->1	f->4	i->7	j->3	k->4	l->2	m->9	n->1	o->19	p->3	r->5	s->5	u->3	v->1	ö->1	
lades	 ->17	
lafra	n->1	
lag -	 ->2	
lag 1	 ->2	,->2	0->5	1->1	2->1	3->1	5->1	7->1	8->2	9->2	
lag 2	,->2	2->3	3->1	6->1	
lag 3	 ->1	4->1	8->3	
lag 4	 ->1	.->2	3->1	4->1	5->3	
lag 5	,->2	
lag 6	 ->2	
lag a	n->2	t->4	v->8	
lag b	e->4	i->1	ö->4	
lag d	e->1	ä->2	
lag e	l->1	n->2	t->1	
lag f	r->19	ö->16	
lag g	e->4	r->1	ä->1	å->1	
lag h	a->10	e->1	ä->4	
lag i	 ->18	n->5	
lag j	a->1	
lag k	a->6	o->1	
lag l	a->1	
lag m	e->1	o->1	å->1	
lag n	i->1	u->1	ä->2	
lag o	c->15	m->19	s->1	
lag p	å->2	
lag r	ö->3	
lag s	k->7	o->52	p->1	t->1	y->2	å->1	
lag t	a->1	i->57	o->1	y->1	
lag u	n->2	
lag v	a->1	e->1	i->3	
lag ä	r->4	
lag å	t->1	
lag ö	v->1	
lag, 	d->3	e->2	f->4	g->1	h->1	i->2	l->2	m->4	n->1	o->4	s->8	t->2	u->2	v->4	
lag. 	H->1	
lag.)	F->2	H->1	
lag..	 ->1	
lag.B	e->1	
lag.D	e->6	i->1	ä->2	
lag.F	r->2	ö->3	
lag.H	e->4	
lag.I	 ->2	
lag.J	a->6	
lag.K	o->1	
lag.L	å->1	
lag.M	e->1	å->1	
lag.P	a->1	
lag.S	y->1	
lag.T	i->1	
lag.U	n->1	
lag.V	a->1	i->2	å->1	
lag; 	s->1	
lag?D	e->1	
lag?F	i->1	r->1	
laga 	2->1	a->3	d->3	n->1	
laga!	F->1	
laga.	D->1	F->1	
lagad	e->2	
lagan	 ->2	d->5	s->3	
lagar	 ->26	,->4	.->4	e->21	m->14	n->3	ä->1	
lagat	 ->1	
lagd 	a->1	i->1	o->1	p->1	
lagd,	 ->1	
lagda	 ->6	.->1	
lagel	s->3	
lagen	 ->67	,->5	.->8	s->3	
lager	.->1	k->1	
laget	 ->51	,->5	.->11	:->1	s->3	
lagfö	r->5	
lagg 	d->1	f->1	i->1	m->1	o->1	s->1	
lagg,	 ->7	
lagg.	D->1	F->1	K->1	M->1	N->1	
lagg;	 ->1	
lagga	 ->2	d->2	n->1	
lagge	n->2	
laggn	i->1	
laggo	r->1	
lagit	 ->8	.->3	s->5	
lagli	g->18	
lagna	 ->15	.->1	
lagni	n->17	
lagom	 ->1	å->3	
lagor	 ->2	?->1	n->2	
lagos	k->1	
lagra	n->1	r->1	
lagre	n->1	
lags 	a->1	f->2	i->2	o->1	p->1	r->2	s->3	u->2	v->1	
lagsd	e->1	
lagsf	ö->1	
lagsk	r->1	
lagst	a->1	i->127	
lagt 	4->1	a->3	e->1	f->28	i->1	m->1	n->10	s->1	
lagt,	 ->1	
lagte	x->2	
lagts	 ->26	
lai L	a->7	
lak s	a->1	
lakta	r->1	
lakti	g->24	
lam f	ö->2	
lam l	i->1	
lam, 	s->1	
lamen	t->600	
lamer	a->2	
lamod	 ->2	
lampo	r->1	
lamsk	y->4	
lamt 	u->1	
lan 1	5->1	9->5	
lan 8	 ->2	
lan C	E->1	e->1	
lan D	a->1	
lan E	r->1	u->9	
lan G	a->1	
lan H	a->1	
lan I	s->9	
lan P	a->1	o->2	
lan S	P->1	y->2	
lan a	k->1	l->1	r->2	v->1	
lan b	e->2	
lan c	h->1	
lan d	e->30	i->1	r->1	
lan e	k->2	m->1	n->4	t->1	
lan f	a->2	o->1	r->2	ö->15	
lan g	e->1	o->1	
lan h	j->1	ö->1	
lan i	t->1	
lan k	a->1	l->1	o->8	u->1	v->4	ö->3	
lan l	e->1	o->3	ä->2	
lan m	e->14	o->1	ä->1	
lan n	a->4	
lan o	c->4	l->3	r->1	s->1	
lan p	a->4	e->2	o->1	r->1	
lan r	a->1	e->14	i->1	å->3	
lan s	e->1	k->1	o->2	t->7	v->1	y->2	å->1	
lan t	j->1	r->1	
lan u	n->2	p->1	t->5	
lan v	e->5	i->2	
lan Ö	s->1	
lan ä	g->1	r->1	
lan" 	g->1	
lan".	R->1	
lan, 	a->1	o->2	s->1	t->1	ä->1	
lan. 	D->1	
lan.D	e->2	
lan.E	n->1	
lan.I	 ->1	l->1	
lan.J	a->1	
lan.S	l->1	
lan.U	n->1	
lan.V	i->1	
lan: 	A->1	
lan?H	e->1	
lanNä	s->1	
lana 	h->1	o->1	
lana,	 ->2	
lanca	,->1	
land 	-->4	8->1	E->1	S->1	T->1	a->27	b->4	d->17	e->6	f->4	g->4	h->7	i->14	k->5	l->2	m->9	n->4	o->22	p->2	r->2	s->29	t->7	u->5	v->7	ä->10	ö->1	
land)	,->1	
land,	 ->31	
land.	D->4	E->1	G->1	I->6	J->5	K->1	L->1	M->2	N->2	O->2	S->1	U->1	V->1	Å->1	
landa	 ->5	d->9	r->3	t->1	
lande	 ->144	!->1	,->10	.->14	;->1	n->42	r->2	s->1	t->69	v->2	
landn	i->10	
lands	 ->10	,->1	b->42	k->2	m->9	p->3	v->1	ä->1	
landv	i->2	
lanen	 ->7	,->1	.->4	s->1	
laner	 ->18	,->1	.->2	a->37	i->20	n->7	
lanet	 ->1	,->1	.->1	
lang,	 ->1	
lange	r->1	s->6	
lanhö	j->4	
lanke	s->1	
lankl	a->1	
lanko	.->1	
lankt	 ->1	
lanli	g->1	
lanni	v->1	
lans 	-->1	a->1	i->1	m->6	o->1	s->5	v->1	
lans,	 ->2	
lanse	n->10	r->12	
lansl	a->1	
lanst	a->5	o->2	
lansv	a->1	
lanså	t->1	
lansö	v->1	
lanta	t->1	
lante	n->4	r->3	
lanti	n->1	q->1	
lantk	u->1	
lantl	i->1	
lanto	r->1	
lanös	t->19	
lappa	 ->1	
lapph	e->3	
lappj	a->1	
lapps	s->1	
lappv	e->2	
lar "	ö->1	
lar -	 ->4	
lar 2	6->1	
lar a	l->2	n->2	t->3	v->18	
lar b	e->1	y->1	å->1	ö->1	
lar d	e->27	o->1	ä->3	
lar e	m->1	n->4	t->2	
lar f	i->1	l->1	r->9	ö->13	
lar g	i->2	
lar h	a->1	e->3	ä->1	å->1	
lar i	 ->16	n->14	
lar j	a->3	u->1	
lar k	a->1	o->3	
lar l	e->1	i->1	
lar m	a->2	e->16	i->6	y->1	å->1	
lar n	a->2	u->1	ä->3	
lar o	c->17	m->96	r->1	
lar p	o->2	r->1	å->7	
lar r	e->2	ä->3	
lar s	a->2	i->8	k->3	o->20	p->2	å->4	
lar t	i->5	j->1	
lar u	n->3	p->2	t->2	
lar v	a->1	e->2	i->4	ä->1	å->2	
lar ä	r->5	v->3	
lar å	t->1	
lar, 	a->1	b->1	d->5	e->3	g->2	i->2	k->2	l->1	m->5	o->2	s->1	u->1	v->1	ä->1	å->2	
lar.B	l->1	
lar.D	e->10	
lar.E	f->1	
lar.F	ö->2	
lar.I	 ->2	n->2	
lar.J	a->7	
lar.K	o->1	
lar.M	e->2	
lar.V	i->4	
lar: 	F->1	
lar; 	i->1	
lar?K	o->1	
lar?N	a->1	
lara 	a->5	d->4	e->1	f->5	h->3	m->3	o->7	p->1	r->2	t->2	u->1	v->1	ö->1	
lara,	 ->1	
lara.	D->1	V->1	
larad	 ->1	e->4	
larar	 ->29	
laras	 ->5	
larat	 ->4	s->1	
larbe	t->1	
lare 	4->1	a->1	b->3	e->3	f->3	h->5	i->2	k->1	m->2	o->4	r->1	s->5	v->1	
lare,	 ->8	
lare.	D->2	K->1	
laren	 ->3	)->2	,->4	.->5	
larfo	r->1	
larfä	r->1	
largö	r->17	
larhe	t->12	
larin	g->24	
laris	e->1	k->2	
larla	g->3	
larlä	g->2	
larmr	a->2	
larms	i->2	
larn 	-->1	s->1	
larna	 ->40	,->4	.->10	?->1	s->5	
lars 	o->2	
larst	o->1	
lart 	-->1	a->35	b->3	e->1	f->12	h->2	i->7	l->1	n->1	o->10	p->1	s->5	t->1	u->2	v->1	ä->3	
lart,	 ->2	
lart.	M->1	
lart:	 ->1	
larte	c->4	x->3	
larti	d->2	
larve	r->1	
lary 	o->1	
las a	v->7	
las b	o->1	
las d	e->3	
las e	f->3	l->1	n->6	
las h	ä->1	
las i	 ->12	n->4	
las k	o->2	
las l	i->1	
las m	e->3	
las n	ä->1	å->1	
las o	c->6	f->1	m->4	
las p	å->9	
las s	a->2	o->2	å->2	
las t	i->9	
las u	n->5	p->1	t->2	
las v	a->1	i->1	å->2	
las y	t->2	
las ö	g->1	
las, 	b->1	e->1	h->1	m->1	o->1	r->1	s->1	u->1	
las.B	l->1	
las.D	e->3	ä->1	
las.K	o->2	
las.T	a->1	
las: 	e->1	
lashu	s->1	
lasia	t->2	
lasie	n->4	
laspe	k->1	
lass 	e->1	f->1	
lassa	s->1	
lasse	n->2	r->1	
lassi	f->9	g->1	s->5	
lassp	e->1	
last 	f->2	m->1	s->1	ä->1	
last!	D->1	
last,	 ->2	
last-	 ->1	
last.	D->1	
lasta	d->3	n->1	r->1	s->1	
laste	 ->2	n->4	
lasti	n->1	
lastn	i->6	
lat "	K->1	e->1	
lat B	r->1	
lat a	n->3	r->1	t->5	
lat d	e->3	
lat e	n->4	r->1	
lat f	r->1	å->1	ö->3	
lat g	e->1	å->1	ö->1	
lat h	a->2	ö->1	
lat i	 ->2	n->2	
lat k	ö->1	
lat m	y->1	
lat n	ä->1	ö->1	
lat o	m->7	s->2	
lat p	å->1	
lat s	i->2	o->1	å->1	
lat u	t->3	
lat v	ä->1	
lat ö	v->1	
lat, 	a->1	i->1	o->2	s->1	
lat.H	e->1	
lat.I	 ->1	
lat.V	a->1	
later	 ->1	a->13	
lath 	h->1	n->1	o->1	
lath,	 ->1	
latio	n->19	
lativ	 ->6	a->2	t->7	
latla	n->1	
laton	s->1	
lator	e->2	
lats 	-->2	S->2	a->4	d->2	f->4	i->7	m->1	o->2	p->1	s->1	t->2	u->6	v->1	
lats,	 ->7	
lats.	D->2	F->1	K->1	
latse	n->5	r->14	
latta	 ->1	
laude	 ->1	
lausu	l->6	
lautr	e->2	
lavan	o->2	
lavar	.->1	s->1	
laver	e->1	
lavie	n->1	
lavta	l->1	
law, 	s->1	
law.M	e->1	
layab	e->1	
layed	 ->2	
lbacè	t->1	
lbaka	 ->35	.->4	?->1	d->3	g->4	v->4	
lbaks	 ->1	
lban 	s->1	
lbane	r->5	
lbani	e->1	
lbank	e->7	s->1	
lbans	k->4	
lbar 	e->2	o->1	p->2	s->2	t->1	u->12	
lbara	 ->6	
lbarh	e->2	
lbart	 ->16	,->1	.->2	
lbefo	l->2	
lbelo	p->1	
lbert	 ->1	
lberä	k->1	
lbes 	a->1	ä->1	
lbesl	u->1	
lbest	ä->4	å->1	
lbild	n->1	
lbloc	k->1	
lbord	a->3	
lbran	s->1	
lbrig	h->1	
lbrin	g->4	
lbrot	t->1	
lbund	e->11	n->4	
lbyrå	k->1	
ld Wi	d->1	
ld av	 ->3	
ld be	k->1	t->2	
ld bo	m->1	
ld fr	å->5	
ld fu	n->1	
ld i 	f->1	v->1	
ld in	o->1	t->1	
ld kl	a->1	
ld ko	m->1	n->1	
ld ku	l->1	
ld ma	n->1	
ld me	d->1	
ld mi	t->1	
ld oc	h->2	
ld pa	r->1	
ld pe	r->1	
ld po	l->1	
ld pu	b->1	
ld på	 ->1	
ld re	g->2	
ld ro	l->1	
ld so	m->1	
ld ta	n->1	
ld ti	l->1	
ld to	n->1	
ld up	p->2	
ld är	 ->1	
ld åt	a->1	
ld, d	e->1	ä->1	
ld, k	o->1	
ld, m	a->1	e->2	
ld, o	c->3	
ld, s	o->1	
ld.De	t->1	
ld.Fö	r->1	
ld.Ja	g->2	
ld.Nu	 ->1	
lda b	e->1	
lda d	e->1	j->1	o->1	
lda e	k->1	n->3	
lda f	a->2	o->1	r->1	ö->5	
lda i	 ->3	n->3	
lda k	o->1	ä->1	
lda l	a->1	ä->1	
lda m	e->4	i->1	å->2	
lda n	a->1	
lda o	c->1	m->1	
lda p	a->3	o->1	r->1	
lda r	a->1	e->3	ä->1	ö->1	
lda s	k->2	o->1	t->4	ä->3	
lda t	i->1	o->1	r->2	
lda v	i->2	
lda ä	r->1	
lda å	t->3	
lda, 	m->3	s->2	
lda.D	e->1	
lda.E	t->1	
lda.H	e->1	
lda.J	a->2	
lda.Ä	r->1	
lda?F	r->1	
ldade	 ->3	
ldage	n->1	
ldand	e->6	
ldar 	a->1	d->2	e->1	r->1	s->1	
ldas 	i->4	r->1	t->1	
ldas,	 ->1	
ldas.	I->1	
ldas?	H->1	
ldast	e->1	
ldat 	k->1	
ldate	r->2	
ldats	 ->2	
ldbel	ä->1	
ldbes	t->1	
lde B	u->1	
lde K	i->1	
lde a	t->1	
lde d	e->5	
lde e	n->2	t->2	
lde f	r->2	ö->2	
lde h	a->1	
lde j	o->1	
lde m	e->1	
lde n	ä->1	å->1	
lde o	c->1	
lde t	r->1	
lde u	n->1	
lde å	r->1	
lde, 	u->1	
lde.E	u->1	
ldela	d->4	r->4	t->5	
ldele	s->23	
ldeln	i->3	
ldelt	a->3	
ldemo	k->16	
lden 	-->2	a->2	f->3	g->2	h->1	i->3	m->2	o->3	p->1	s->5	u->2	ä->1	
lden,	 ->9	
lden.	H->1	I->1	J->2	
lden:	 ->1	
lden?	V->1	
ldens	 ->4	
lder 	a->2	e->1	m->1	r->1	s->2	
lder.	 ->1	B->1	D->1	
lderd	o->2	
ldern	 ->2	a->1	
ldes 	A->1	a->1	b->1	d->3	i->4	m->1	
ldes.	I->1	
ldet 	m->1	
ldet,	 ->1	
ldez,	 ->1	
ldez-	k->2	
ldgrä	n->1	
ldhet	 ->7	e->3	s->13	
ldig 	a->1	f->1	n->1	
ldiga	 ->10	.->1	n->3	
ldige	s->1	
ldigh	e->15	
ldigt	 ->21	
ldiox	i->5	
ldire	k->17	
ldist	r->1	
ldjur	,->1	
ldnin	g->66	
ldoms	t->1	
ldra 	e->1	r->1	s->1	
ldrad	e->3	
ldrag	e->1	
ldrar	 ->1	
ldrat	s->2	
ldre 	e->1	f->2	ä->2	
ldre,	 ->1	
ldre.	D->1	
ldrig	 ->32	
ldsam	 ->2	m->1	
ldsde	l->1	
ldsek	o->1	
ldsfr	å->1	
ldsha	n->6	
ldskr	i->6	
ldsli	g->1	
ldsma	r->1	
ldsni	v->1	
ldsom	s->1	
ldsut	t->1	
ldta 	j->1	
ldtag	i->1	
le - 	o->1	
le Eu	r->3	
le Ki	n->1	
le al	l->3	
le an	t->3	
le at	t->18	
le av	s->1	
le ba	r->3	
le be	a->1	g->1	h->3	s->1	t->2	v->1	
le bi	d->1	
le bl	i->5	
le bé	b->1	
le bö	r->2	
le de	 ->4	l->1	n->3	s->2	t->18	
le do	c->3	
le dä	r->8	
le då	 ->2	
le el	i->1	
le em	e->1	
le en	 ->4	g->1	
le ev	e->1	
le fa	k->1	
le fi	n->2	
le fr	a->2	ä->1	å->1	
le få	 ->4	
le fö	l->1	r->19	
le ge	 ->1	n->1	
le go	d->1	
le gr	a->1	
le gä	l->2	r->5	
le gå	 ->1	
le gö	r->5	
le ha	 ->14	m->1	n->2	r->1	
le he	n->1	
le hä	n->1	r->2	v->1	
le i 	a->1	f->1	m->2	o->1	p->1	
le in	f->2	k->1	n->6	r->2	s->1	t->8	
le ja	g->44	
le ka	n->1	
le ko	m->4	n->1	r->1	
le kr	ä->2	
le ku	n->56	
le kä	n->1	
le le	d->3	v->1	
le lä	g->1	
le ma	n->2	
le me	d->2	
le mo	t->1	
le na	t->1	
le ni	 ->1	
le nu	 ->1	
le nä	r->1	
le oc	h->5	k->7	
le of	r->1	
le ol	j->1	
le pa	r->2	s->1	
le pl	a->1	
le po	s->1	
le på	 ->2	
le re	a->1	d->1	
le rä	c->1	
le rå	d->1	
le rö	s->1	
le sa	n->1	
le se	 ->1	
le sj	ä->1	
le sk	a->4	e->1	
le sl	u->2	
le so	m->3	p->1	
le sp	e->1	
le st	r->1	å->2	
le sv	a->1	
le sä	g->1	k->1	r->1	t->1	
le så	l->6	
le sö	n->1	
le t.	e->1	
le ta	 ->4	c->1	
le ti	l->5	
le tr	o->1	
le tv	i->1	ä->1	
le un	d->3	
le up	p->4	
le ur	h->2	v->1	
le ut	?->1	g->1	s->1	t->1	v->1	ö->1	
le va	n->1	r->36	
le ve	r->2	
le vi	 ->8	a->1	d->2	l->69	s->1	
le vä	c->1	n->1	r->1	
le än	d->1	
le är	 ->2	
le äv	e->1	
le åt	e->1	m->1	
le ön	s->2	
le, o	c->1	m->2	
le-de	-->2	
le.Ja	g->1	
le.Vi	 ->1	
led i	 ->1	
led m	e->1	
leda 	a->2	d->4	e->7	f->5	i->2	m->3	o->3	p->1	t->30	
leda,	 ->1	
ledam	o->71	ö->83	
ledan	d->14	
ledar	e->7	f->1	n->5	s->1	
ledas	 ->5	,->1	
ledda	 ->3	
ledde	 ->13	s->7	
leder	 ->38	,->2	
ledes	 ->44	
ledig	h->1	
ledni	n->74	
leds 	b->1	i->1	r->1	u->1	å->1	
ledse	n->2	
ledst	j->2	
lefan	t->1	
lefon	,->1	
lega 	B->3	E->2	F->6	H->1	J->3	K->1	L->1	M->1	N->2	R->2	S->1	a->1	b->1	d->1	f->2	k->1	s->2	t->1	v->4	
lega!	 ->1	D->1	J->1	Ä->1	
lega,	 ->3	
lega.	J->1	
legad	.->1	e->1	
legal	 ->4	a->7	i->2	t->9	
legan	 ->16	
legas	 ->2	
legat	 ->3	i->16	
lege.	O->1	
lege?	H->1	
leger	 ->34	!->65	,->14	.->4	:->1	a->3	i->1	n->8	s->1	
legie	r->3	t->2	
legit	i->18	
legiu	m->3	
legor	 ->1	i->1	s->2	
lehan	d->3	
leido	s->2	
lejda	 ->1	
lejdo	s->1	
lekas	t->1	
leken	 ->1	,->1	
leker	 ->1	
lekom	m->3	
lekon	o->4	
leksa	k->1	
lekte	r->3	
lekti	o->5	v->11	
lektr	i->1	o->9	
lektu	e->3	
lekty	r->1	
leler	s->3	
lella	 ->2	
lellt	 ->3	
lelse	 ->7	,->1	n->1	
lem -	 ->1	
lem a	v->2	
lem d	e->2	
lem e	f->2	n->1	
lem f	ö->3	
lem h	a->2	ä->1	
lem i	 ->10	n->3	
lem k	a->1	o->1	
lem m	e->12	
lem n	i->1	ä->3	
lem o	c->6	m->1	
lem p	å->1	
lem s	o->17	
lem u	r->1	
lem v	a->1	i->2	
lem ä	r->4	
lem ö	v->1	
lem, 	a->1	b->1	e->1	g->1	m->2	o->3	p->2	u->1	v->2	
lem. 	M->1	
lem..	 ->1	
lem.A	l->1	
lem.D	e->5	ä->1	
lem.F	ö->1	
lem.H	e->2	
lem.I	n->1	
lem.J	a->3	
lem.M	å->1	
lem.P	r->1	
lem.S	l->1	o->1	
lem.V	e->1	i->2	
lem: 	A->1	
lem; 	d->2	
lem?M	e->1	
lemat	i->5	
lemen	 ->16	,->1	t->20	
lemet	 ->41	,->3	.->3	s->1	
lemik	 ->1	
lemlä	s->1	
lemma	 ->2	:->1	r->14	
lemom	r->3	
lemsk	a->2	
lemsl	a->9	ä->27	
lemsr	e->1	
lemss	t->284	
len B	r->1	
len E	r->1	
len a	l->1	n->1	t->4	v->21	
len b	e->5	r->1	ö->1	
len d	ä->1	å->2	
len e	f->2	l->1	r->1	
len f	r->5	ö->11	
len g	e->1	o->1	
len h	a->8	
len i	 ->26	n->7	
len k	a->1	o->3	ä->1	
len m	e->8	å->1	
len n	u->1	ä->1	
len o	c->12	m->1	
len p	å->2	
len s	j->1	k->4	l->1	n->1	o->11	
len t	a->1	i->5	
len u	n->2	t->4	
len v	i->3	
len ä	l->1	n->1	r->2	
len å	s->1	t->2	
len ö	v->1	
len" 	i->1	o->1	
len",	 ->1	
len, 	1->2	8->1	V->1	d->6	e->1	f->1	h->1	i->2	j->1	k->1	m->2	n->1	o->5	s->3	t->1	u->1	v->1	ä->1	
len. 	V->1	
len.A	l->1	
len.D	e->9	ä->1	
len.E	t->1	
len.H	e->3	
len.I	 ->1	n->1	
len.J	a->3	
len.K	a->1	o->1	v->1	
len.M	a->1	e->4	
len.R	e->1	
len.S	k->1	t->1	
len.T	y->1	
len.U	t->1	
len.V	a->1	i->3	
len?Ä	r->1	
lenFr	å->2	
lena 	f->1	k->1	r->1	s->1	
lena,	 ->1	
lenar	s->4	å->1	
lenni	e->5	u->2	
lens 	b->2	d->2	e->1	o->2	r->1	s->1	u->1	ö->1	
lensk	a->1	
lenti	n->1	
lenum	 ->4	.->1	
lenÄr	a->1	
lenät	 ->1	
leote	 ->1	
ler -	 ->3	
ler 2	0->1	
ler 7	3->1	
ler 8	0->1	
ler 9	0->1	
ler A	l->2	z->1	
ler D	a->1	
ler E	M->1	u->7	
ler F	i->1	ö->3	
ler I	t->1	
ler J	a->1	
ler L	y->1	
ler M	e->1	
ler N	e->1	
ler P	V->1	a->1	
ler R	a->1	u->1	
ler S	c->2	h->1	k->1	y->1	
ler T	o->1	u->2	
ler U	S->1	r->1	
ler a	k->1	l->8	n->19	r->3	t->33	v->9	
ler b	a->2	e->12	i->4	l->5	o->1	r->4	u->1	å->1	ö->1	
ler c	i->2	
ler d	a->2	e->101	i->1	o->2	u->3	ä->2	å->2	ö->1	
ler e	f->3	g->1	j->7	k->4	m->5	n->27	r->4	t->13	u->1	x->1	
ler f	a->5	e->1	i->4	l->5	o->5	r->21	u->1	å->2	ö->54	
ler g	e->9	l->1	o->3	r->5	y->1	å->1	ö->2	
ler h	a->7	e->5	j->1	o->1	u->4	ä->2	ö->1	
ler i	 ->13	c->1	f->1	g->1	m->1	n->53	
ler j	a->3	o->1	ä->1	
ler k	a->8	e->1	l->1	n->1	o->18	r->7	v->4	ä->3	ö->1	
ler l	a->4	e->4	i->4	o->1	ä->6	å->4	
ler m	a->7	e->27	i->19	o->2	u->1	y->4	ä->2	å->1	ö->3	
ler n	a->1	e->2	o->1	u->1	y->2	ä->5	å->8	
ler o	a->1	b->1	c->26	f->1	k->1	l->1	m->20	r->4	s->5	ö->1	
ler p	a->4	e->2	o->2	r->7	u->1	å->26	
ler r	a->4	e->5	i->3	ä->2	å->1	ö->1	
ler s	a->6	e->4	i->15	j->2	k->6	l->2	m->1	o->21	p->2	t->12	u->1	v->3	y->2	ä->5	å->2	ö->2	
ler t	.->1	a->2	i->14	j->2	o->2	r->7	u->2	v->2	
ler u	n->5	p->2	t->13	
ler v	a->12	e->3	i->15	ä->2	å->5	
ler Ö	s->2	
ler ä	l->1	n->10	r->6	v->4	
ler å	r->1	t->7	
ler ö	k->1	p->1	r->1	v->4	
ler, 	a->1	b->1	e->1	g->1	h->1	k->1	m->4	n->1	o->2	s->2	t->3	u->1	v->1	
ler-r	e->1	
ler.A	v->1	
ler.D	e->6	
ler.E	f->1	
ler.F	å->1	ö->2	
ler.H	e->2	
ler.J	a->3	
ler.K	a->1	
ler.M	e->1	ä->1	
ler.O	m->1	
ler.R	e->1	
ler.Ä	n->1	
ler; 	d->1	
ler?P	å->1	
lera 	-->1	2->1	L->1	a->13	b->2	d->4	e->8	f->10	g->11	h->10	i->1	k->4	l->3	m->8	n->2	o->10	p->4	s->9	t->5	u->2	Ö->2	ä->2	å->5	ö->1	
lera"	.->1	
lera,	 ->1	
lera.	D->1	
lerad	 ->5	e->7	
leran	d->1	s->11	
lerar	 ->19	!->1	
leras	 ->15	,->3	.->3	
lerat	 ->7	s->3	
lerer	a->7	
leri 	a->1	f->2	o->1	
lerie	t->1	
lerin	g->25	
lerkä	n->3	
lermo	,->1	
lerna	 ->35	,->6	.->10	s->1	
lers 	j->1	l->1	
lerst	a->1	
lersu	n->3	
lerta	l->6	
lerti	d->67	
lerår	i->12	
les G	i->1	
les a	t->1	v->1	
les e	g->1	l->1	
les f	ö->8	
les h	a->1	i->1	
les i	 ->1	
les j	u->1	
les k	l->1	
les n	y->4	
les p	å->1	
les r	i->2	o->1	ä->3	
les s	j->1	l->1	o->1	p->1	t->1	ä->1	
les t	v->1	
les u	t->2	
les.H	u->1	
les.V	a->1	
les; 	o->1	
lesa 	b->1	
lesam	m->5	
lesar	e->1	
lese 	i->1	
leska	t->1	
lesma	n->1	
lesmä	n->1	
lesnå	l->4	
lesta	 ->25	
lesti	n->22	
lesät	t->2	
let -	 ->1	
let A	l->1	
let E	U->1	
let T	V->1	
let V	e->1	o->1	
let a	n->1	r->1	t->8	v->5	
let b	l->1	o->1	å->1	ö->1	
let d	e->3	
let e	f->2	n->3	u->2	
let f	e->1	i->2	o->1	r->12	ö->25	
let g	e->1	ä->2	å->1	
let h	a->6	j->1	o->2	ä->2	
let i	 ->21	n->5	
let j	u->1	
let k	a->1	e->1	o->2	r->2	
let l	e->2	i->1	
let m	e->19	å->3	
let n	a->1	ä->1	
let o	c->9	l->2	m->9	
let p	o->1	
let r	e->3	i->1	ä->2	
let s	a->1	k->4	l->1	o->3	p->1	t->4	
let t	a->1	i->10	j->1	ä->2	
let u	n->1	p->1	
let v	a->1	e->4	i->1	
let Ö	s->1	
let ä	r->10	
let å	t->1	
let ö	v->1	
let!P	r->1	
let, 	a->3	d->1	e->1	f->1	h->1	i->1	k->1	m->6	o->4	p->1	s->5	u->3	v->3	
let. 	D->1	
let.)	R->1	
let.A	v->2	
let.D	e->11	
let.F	r->1	
let.H	e->2	
let.I	 ->1	n->1	
let.J	a->7	
let.K	o->1	
let.N	ä->1	
let.O	r->1	
let.S	o->1	t->1	
let.T	r->1	
let.U	n->1	
let.V	i->4	
let: 	d->1	
letar	 ->1	
lets 	B->1	a->1	f->1	k->1	m->1	s->1	
lett 	e->2	f->1	o->1	s->2	t->8	
lette	r->13	
letts	 ->6	,->1	.->3	
leum 	v->1	
leuro	p->3	
lev a	n->1	v->2	
lev d	j->1	ä->1	
lev f	a->1	ö->1	
lev i	n->2	
lev k	v->1	
lev o	b->2	c->1	
lev t	v->1	
lev u	n->1	
leva 	d->1	e->2	f->1	h->1	i->4	l->1	m->2	n->1	p->1	s->1	u->1	v->1	
leva,	 ->1	
leva?	N->1	
levan	d->3	t->9	
levde	 ->2	
leveb	r->1	
level	 ->1	s->1	
lever	 ->12	.->1	a->3	e->4	
levis	i->1	
levna	d->12	
levs 	o->1	s->2	
levt 	d->1	e->2	i->1	
lewoo	d->2	
lex f	l->1	
lex.J	a->1	
lexa,	 ->1	
lexan	d->2	
lexib	e->11	i->10	l->6	
lext 	o->1	
lez o	c->1	
lf Hi	t->2	
lf-Ma	t->2	
lfabe	t->1	
lfede	r->1	
lfen 	o->1	ä->1	
lfen.	I->1	Ä->1	
lferi	e->1	
lfing	e->1	
lfkri	g->1	
lfoga	 ->5	r->1	
lfond	e->15	
lford	-->1	o->2	
lfram	g->3	
lfred	s->27	
lfrih	e->2	
lfråg	a->2	o->7	
lfstr	ö->3	
lfte 	g->1	
lften	 ->3	
lfunk	t->2	
lfunn	a->1	
lfäll	e->87	i->10	
lfärd	 ->1	,->2	;->1	s->5	
lfång	s->4	
lfölj	a->2	e->1	
lför 	E->1	d->2	
lför.	D->1	
lföra	 ->1	s->1	
lförb	u->4	
lföre	t->7	
lförf	a->2	
lförl	i->4	
lförs	a->2	i->2	t->1	v->2	ä->7	
lförv	a->2	
lgado	,->1	
lgari	e->1	
lgeme	n->1	
lgen 	t->1	
lgeri	e->1	
lgien	 ->5	,->2	?->1	s->1	
lgisk	 ->2	a->6	
lgivn	i->1	
lgjor	t->1	
lgodo	s->1	
lgrip	a->1	e->1	
lgrun	d->2	
lgäng	l->21	
lgång	 ->19	,->1	a->1	e->4	
lgåvo	r->1	
lgöra	 ->1	n->1	
lhand	a->43	
lhava	r->1	
lhave	t->1	
lhavs	l->1	o->1	
lhelm	s->1	
lhet 	a->1	f->2	i->1	k->1	m->1	o->1	s->1	u->1	ä->1	å->1	
lhet,	 ->7	
lhet.	N->1	
lhet?	 ->1	
lhete	n->1	
lhets	k->1	p->1	s->1	
lhjär	t->8	
lhoek	 ->1	
lhör 	d->1	e->1	i->1	n->1	
lhöra	 ->2	n->1	
lhöri	g->1	
li - 	e->1	
li 19	9->4	
li 20	0->3	
li ak	t->1	
li al	l->2	
li an	n->1	s->1	
li at	t->4	
li av	f->1	g->1	
li be	g->1	s->1	v->1	
li br	a->1	
li bä	t->1	
li de	n->1	t->2	
li do	m->2	
li ef	f->2	
li en	 ->18	
li et	t->11	
li fl	e->2	
li fr	å->1	
li fä	r->1	
li fö	r->9	
li ga	r->1	
li ha	r->1	
li he	l->1	
li ju	s->1	
li kl	a->3	
li ko	m->1	
li le	v->1	
li li	k->2	
li lä	t->1	
li me	d->5	r->6	
li mi	g->1	n->1	
li my	c->4	n->1	
li mö	j->3	
li nä	r->1	
li nå	g->2	
li nö	d->1	j->1	
li ob	l->1	
li om	 ->1	
li ot	y->1	
li pl	a->1	
li pr	e->2	
li ri	k->1	
li sl	u->1	
li st	e->1	o->1	ö->1	
li su	b->1	
li sv	å->1	
li sy	n->1	
li sä	m->1	
li så	 ->1	
li tv	u->3	
li un	d->1	
li va	k->1	
li ve	r->2	
li vå	r->1	
li äm	n->1	
li öv	e->2	
li!Ja	g->1	
li, e	n->1	
li, m	e->1	
li, o	c->1	
li.Ut	v->1	
lia-R	o->1	
lians	 ->3	e->4	
libak	t->1	
liban	e->1	
libbi	g->1	
liber	a->29	
libi 	n->1	
lic -	 ->1	
lican	t->1	
licen	s->1	
licer	a->15	i->1	
licie	n->2	
licit	.->1	e->1	
lick 	a->1	b->1	e->1	f->1	
lick,	 ->1	
lick.	H->1	K->1	
licka	 ->2	
lickb	a->5	
licke	n->1	t->9	
licko	r->1	
licy,	 ->1	
licya	v->1	
licyd	e->1	
licyf	ö->1	
lida 	s->1	
lidan	d->2	
lidar	i->30	
lider	 ->7	a->1	i->2	
lidit	 ->3	
lien 	e->2	f->2	h->3	o->3	t->1	ä->1	
lien,	 ->5	
lien.	E->1	M->1	
liens	 ->1	k->17	
lient	i->1	
lier 	e->1	m->1	s->2	
liera	d->1	
liern	a->1	
liest	r->1	
lific	e->14	
lifik	a->1	
lig a	c->1	n->2	r->1	s->2	t->4	v->1	
lig b	e->7	i->1	y->1	
lig d	e->13	i->1	
lig e	f->1	k->1	l->3	u->1	x->1	
lig f	a->1	o->1	r->9	ö->19	
lig g	a->1	r->7	
lig h	a->3	i->2	j->2	ä->2	
lig i	 ->2	n->12	
lig j	o->1	ä->1	
lig k	a->3	o->14	u->2	
lig l	a->4	ö->3	
lig m	a->6	e->3	i->1	o->2	å->1	
lig n	e->1	i->3	o->1	y->1	ä->2	
lig o	c->15	f->2	m->4	n->1	r->1	
lig p	o->5	r->3	å->1	
lig r	a->2	e->7	i->2	y->1	ä->1	å->2	
lig s	a->2	e->5	i->4	k->3	o->3	t->5	u->1	v->1	y->2	ä->2	
lig t	e->1	i->12	o->1	
lig u	p->6	t->14	
lig v	ä->2	
lig y	r->1	
lig å	k->1	s->1	
lig ö	v->2	
lig!H	a->1	
lig, 	a->1	e->1	i->1	n->1	o->2	s->5	v->2	
lig. 	F->1	S->1	
lig.D	e->2	
lig.G	e->1	r->1	
lig.J	a->4	
lig.O	c->3	
lig.V	i->2	
lig: 	d->2	
lig?D	e->1	
lig?H	u->1	
liga 	-->3	3->1	a->20	b->30	c->1	d->13	e->13	f->94	g->15	h->12	i->21	k->27	l->21	m->35	n->6	o->66	p->27	r->66	s->88	t->16	u->12	v->12	y->1	ä->13	å->11	ö->9	
liga,	 ->18	
liga.	(->1	D->2	E->1	F->3	I->2	M->1	N->2	P->2	S->1	V->3	
liga/	h->1	
liga;	 ->1	
liga?	F->1	
ligad	e->1	
ligan	d->5	
ligar	e->67	
ligas	 ->2	,->2	t->6	
ligat	o->14	s->2	
ligen	 ->454	,->18	.->3	:->1	s->1	t->4	
ligga	 ->13	n->10	
ligge	r->86	
liggj	o->12	
liggö	r->21	
lighe	t->333	
lighå	l->2	
ligie	r->1	
ligiö	s->4	
ligse	k->1	
ligt 	-->2	:->1	D->1	E->1	G->1	I->1	K->1	S->1	T->1	a->110	b->16	d->20	e->23	f->55	g->43	h->17	i->26	j->2	k->14	l->8	m->60	n->7	o->42	p->22	r->6	s->86	t->19	u->15	v->30	y->1	ä->5	å->1	ö->3	
ligt!	L->1	M->1	
ligt,	 ->30	
ligt.	D->9	E->1	F->5	G->1	H->5	I->1	J->6	L->1	M->8	N->1	O->3	P->1	S->2	U->1	V->9	Ö->1	
ligt:	 ->1	
ligt;	 ->1	
ligtv	i->101	
lihop	.->1	
lik h	a->1	
lik m	i->1	
lik p	o->1	å->1	
lik.D	e->1	
lik: 	v->1	
lika 	E->1	a->4	b->12	d->4	e->3	f->12	g->7	h->4	i->9	k->8	l->9	m->14	n->8	p->11	r->9	s->18	t->5	u->5	v->11	ä->7	å->3	ö->1	
lika,	 ->1	
lika.	D->1	I->1	J->1	
likab	e->1	
likad	a->2	
likal	y->1	
likan	e->5	s->1	
likar	 ->3	t->2	
likas	å->2	
liken	 ->10	s->1	
liker	,->1	n->3	
likgi	l->2	
likhe	t->35	
likna	n->19	r->2	
likni	n->44	
likri	k->3	
likso	m->47	
likst	ä->2	
likt 	a->3	b->1	d->2	e->1	h->2	i->2	k->1	l->1	m->2	s->1	
likt,	 ->1	
likt.	D->1	O->1	
likta	d->4	
likte	l->13	n->9	r->6	
liktf	ö->1	
likti	g->5	
likvä	l->3	r->5	
lilla	 ->4	
lillf	i->1	
lilli	!->1	
liman	g->3	
limat	 ->1	.->1	e->7	f->4	p->1	
limen	t->1	
limin	e->3	ä->3	
limso	l->1	
lin 1	9->1	
lin b	e->1	
lin f	r->1	ö->1	
lin i	 ->1	
lin n	ä->1	
lin o	c->4	
lin s	t->1	
lin u	n->1	
lin, 	f->1	o->2	
lin.L	i->1	
lin.O	m->1	
linar	b->1	
linba	n->1	
linda	 ->1	.->2	
lindr	a->4	
lindu	s->56	
line 	f->1	
liner	i->2	n->1	
linfr	å->1	
ling 	(->2	a->23	e->2	f->5	g->1	h->2	i->13	k->6	l->2	m->3	n->1	o->16	p->1	r->2	s->15	u->1	v->3	ä->2	
ling,	 ->25	
ling.	 ->1	D->7	F->2	H->2	I->3	J->3	K->1	M->3	N->2	O->3	V->2	
linga	n->1	r->75	
linge	n->89	
lings	-->3	a->4	b->3	c->3	f->42	g->1	k->6	l->1	m->5	n->1	o->1	p->29	r->8	s->8	t->1	u->4	ä->1	
linis	t->2	
linje	 ->11	.->2	n->3	r->77	
linko	n->2	
linor	n->1	
linri	k->5	
linrå	d->1	
linsb	u->1	
lint 	b->1	
linto	n->1	
lintr	e->1	
linär	a->4	
liote	k->2	
lippe	r->2	
lir E	u->2	
lir a	l->3	n->2	t->4	v->1	
lir b	i->1	r->1	ä->1	
lir d	e->12	i->2	
lir e	n->7	t->3	
lir f	o->1	r->2	ö->3	
lir g	r->1	
lir h	a->1	j->1	o->1	
lir i	 ->2	n->3	
lir j	a->1	u->1	
lir k	o->1	
lir l	a->1	e->1	u->1	ä->2	
lir m	e->4	i->1	y->2	å->1	ö->3	
lir n	a->1	e->1	å->2	ö->1	
lir o	f->1	n->1	t->1	u->1	
lir r	a->1	e->1	ä->1	
lir s	a->2	e->2	k->1	o->1	t->3	v->2	ä->1	å->1	
lir t	i->4	ä->1	
lir u	t->2	
lir v	a->1	e->2	i->1	
lir ä	n->1	
lir å	s->1	
lir ö	v->1	
lir, 	g->1	i->1	
lir: 	O->1	
lirar	 ->1	
lirta	n->1	
lis f	o->1	
lis, 	d->1	
lis.V	i->1	
lis; 	a->1	
lisab	e->1	
lisak	a->1	
lisat	i->1	
lisen	 ->4	s->1	
liser	.->1	a->42	i->37	
lisio	n->3	
lisiä	r->1	
lisk 	m->1	o->1	r->1	ä->1	
lisk,	 ->1	
lisk.	O->1	
liska	 ->17	,->1	
liske	 ->1	
liskt	 ->1	
lism 	e->1	o->3	s->2	ä->1	
lism.	I->2	M->1	
lism?	V->1	
lisme	n->3	
lismy	n->2	
lissa	m->1	
lisse	r->1	
lisst	y->1	
lista	 ->7	,->1	.->6	?->1	N->1	n->47	
liste	 ->2	n->1	r->24	
listg	r->3	
listi	g->2	s->35	
listk	o->1	
listp	a->5	
lists	 ->1	
lisvä	s->1	
lit -	 ->1	
lit a	n->1	t->1	
lit b	o->1	
lit e	n->2	r->1	
lit f	a->1	r->1	
lit h	ö->1	
lit i	 ->1	
lit m	i->1	
lit o	f->2	
lit p	å->2	
lit s	i->1	j->1	t->2	
lit t	y->1	
lit ö	v->1	
lit, 	v->1	
lita 	o->1	p->2	s->1	u->1	
litad	e->1	
litan	o->1	
litar	 ->9	i->4	
litat	.->1	i->6	
lite 	b->1	e->1	i->1	m->1	s->1	
liten	 ->20	.->2	
liter	-->1	i->1	s->1	
litet	 ->52	!->1	,->10	.->7	?->1	e->25	s->11	
litic	a->1	
litik	 ->110	!->1	"->1	,->28	.->24	?->2	e->136	o->6	s->1	
litio	n->14	
litis	k->223	
litli	g->5	
lits 	d->1	h->1	i->2	
lits.	D->1	M->1	
litte	r->8	
littr	a->2	i->2	
litär	 ->2	a->3	e->1	
liv f	r->1	ö->1	
liv i	 ->1	
liv k	o->1	
liv o	a->1	c->1	
liv s	i->1	o->1	
liv t	i->1	
liv, 	s->3	t->1	
liv.A	v->1	
liv.D	e->1	
liv.I	 ->1	
liv.M	e->1	
liv.V	i->1	
liva 	d->1	e->1	f->1	
livad	e->1	
livan	d->8	
livas	 ->4	,->1	.->1	
livat	 ->1	s->3	
livet	 ->12	"->1	,->3	.->6	s->3	
livie	r->1	
livit	 ->26	
livsc	y->3	
livsd	u->2	
livsk	r->1	v->5	
livsm	e->85	i->3	
livsu	p->1	
livsv	i->1	
lixtr	a->1	
lj Li	b->1	
lj om	 ->1	
lj öv	e->1	
lj, o	m->1	
lj, ä	v->1	
lj.Vi	 ->1	
lja -	 ->1	
lja F	N->1	
lja H	a->1	
lja M	a->1	
lja a	n->8	t->8	
lja b	e->12	o->1	ö->5	
lja c	i->1	
lja d	e->6	
lja e	f->1	k->1	l->1	n->5	r->3	t->1	
lja f	o->1	r->13	u->1	ä->1	ö->7	
lja g	e->3	r->4	ö->10	
lja h	a->8	u->1	ä->2	ö->2	
lja i	 ->2	
lja k	n->1	o->2	r->1	
lja l	y->1	ä->2	
lja m	e->1	
lja n	y->1	ä->2	
lja o	c->5	
lja p	e->1	å->7	
lja r	e->1	i->1	ä->3	
lja s	a->1	e->2	i->3	l->1	o->2	v->1	ä->20	
lja t	a->18	i->6	v->1	
lja u	n->5	p->10	r->1	t->5	
lja v	a->3	e->4	i->1	å->1	
lja y	t->1	
lja ö	v->1	
lja, 	f->1	g->1	h->1	p->1	t->1	
lja..	.->1	
lja.J	a->1	
lja.M	i->1	
lja.T	r->1	
ljade	 ->3	
ljakt	i->4	l->14	
ljan 	a->4	f->4	g->1	i->1	o->1	u->1	
ljan,	 ->1	
ljana	l->1	
ljand	e->46	
ljar 	a->2	r->1	s->1	u->1	
ljar.	M->1	
ljarb	a->1	
ljard	 ->1	e->14	
ljare	 ->3	.->2	n->2	
ljarn	a->6	
ljas 	a->4	f->5	o->2	u->1	
ljas,	 ->1	
ljas.	H->2	V->1	
ljat 	a->2	o->1	s->2	
ljats	 ->2	,->1	
ljd a	v->18	
ljd.J	a->1	
ljde 	d->1	p->1	u->1	
ljder	 ->10	n->6	
ljdes	 ->2	
ljdri	k->1	
ljdsk	a->2	
ljdåt	g->1	
lje- 	o->1	
ljebe	f->1	
ljebo	l->4	
ljebä	l->10	
ljedo	m->1	
ljefa	d->1	
ljefö	r->2	
ljein	d->3	
ljejo	r->3	
ljeko	k->1	n->1	
ljeli	n->1	
ljels	e->3	
ljemä	s->1	
ljer 	a->2	d->3	e->1	f->1	g->1	h->2	i->2	m->3	o->4	p->2	r->1	s->12	u->1	v->3	
ljer,	 ->4	
ljer.	D->1	
ljera	d->11	t->5	
ljern	a->4	
ljesk	a->1	
ljest	a->1	
ljeta	n->9	
ljetr	a->1	u->1	
ljeut	s->2	
ljeåt	e->1	
ljflö	d->1	
ljkon	t->2	
ljnin	g->13	
ljon 	i->1	
ljone	r->63	
ljont	a->1	
ljs a	v->1	
ljs k	a->1	
ljs u	p->2	
ljs, 	f->1	
ljt i	 ->1	
ljt u	t->1	
ljt v	i->1	
ljts 	t->1	u->1	
ljudd	a->1	
ljude	r->1	
ljudl	i->1	
ljuge	r->1	
ljus 	p->1	
ljus.	I->1	
ljuse	t->8	
ljö f	ö->2	
ljö i	 ->1	
ljö k	a->1	
ljö m	o->1	
ljö s	a->1	o->1	
ljö v	i->1	
ljö!D	e->1	
ljö, 	f->7	h->1	l->1	s->1	u->1	
ljö- 	o->2	
ljö.D	e->2	å->1	
ljö.M	e->1	
ljö.U	n->1	
ljö.V	i->1	
ljöan	p->1	s->2	
ljöav	t->1	
ljöbe	l->1	s->2	
ljöbr	o->1	
ljöde	p->1	
ljödi	r->1	
ljöer	 ->3	n->1	
ljöfa	k->1	r->1	
ljöfr	å->4	
ljöfö	r->4	
ljöin	f->1	
ljöka	s->1	t->10	
ljöko	n->6	
ljökr	a->8	
ljökv	a->1	
ljöla	g->1	
ljömi	n->1	
ljömä	s->11	
ljömå	l->3	
ljön 	e->2	f->1	h->1	i->1	o->6	p->1	s->1	t->1	ä->1	
ljön!	D->1	
ljön,	 ->9	
ljön.	D->3	E->1	J->1	L->1	M->1	U->1	V->2	
ljöno	r->2	
ljöns	 ->2	
ljöom	r->4	
ljöov	ä->1	
ljöpe	r->1	
ljöpo	l->8	
ljöpr	o->4	
ljöpå	v->1	
ljörå	d->1	
ljörö	r->2	
ljöse	k->1	
ljösi	d->1	
ljösk	a->2	y->11	ä->2	
ljöst	ö->1	
ljösy	n->6	
ljöut	s->1	
ljövä	n->7	r->2	
lk at	t->1	
lk bl	i->1	
lk bo	r->1	
lk ha	r->1	
lk i 	E->1	f->1	
lk oc	h->2	
lk re	a->1	
lk sk	a->1	
lk so	m->2	
lk tv	i->1	
lk up	p->1	
lk, d	e->1	
lk.At	t->1	
lk.De	t->1	
lk.Me	n->1	
lk.Oc	h->1	
lk.Vi	 ->3	l->1	
lka a	v->1	
lka b	e->1	l->1	
lka d	e->8	
lka e	f->1	k->1	m->1	
lka f	a->1	r->2	ö->6	
lka g	a->2	e->2	r->1	
lka i	n->2	
lka j	a->1	
lka k	a->2	o->9	r->3	u->2	
lka l	a->2	i->1	ä->1	
lka m	a->1	e->1	o->1	y->1	å->1	ö->1	
lka n	i->1	y->1	
lka o	f->2	l->1	m->1	
lka p	l->1	r->3	
lka r	ö->1	
lka s	i->1	k->1	l->1	t->4	v->3	ä->1	
lka t	e->1	y->1	ä->1	
lka u	n->2	t->2	
lka v	e->2	i->3	
lka ä	r->8	v->1	
lka å	t->7	
lka ö	v->1	
lkade	 ->1	
lkan 	h->1	i->1	s->1	
lkan.	D->3	O->1	
lkar 	d->3	
lkarn	a->2	
lkas 	d->1	m->1	o->1	s->1	u->1	v->1	
lkas,	 ->1	
lkas.	M->1	
lkast	a->2	
lkats	 ->1	
lkemi	s->1	
lken 	a->1	b->2	d->3	f->5	g->1	h->3	i->9	j->4	k->3	l->3	m->2	n->1	r->2	s->8	t->1	u->5	v->1	å->2	
lken,	 ->1	
lkens	 ->4	
lkest	e->1	
lket 	-->1	B->1	E->2	P->1	V->1	a->3	b->4	d->9	e->4	f->20	g->8	h->7	i->15	j->8	k->5	l->3	m->6	n->5	o->7	p->3	r->7	s->24	t->3	u->4	v->17	ä->17	
lket,	 ->1	
lket.	V->1	
lket:	 ->1	
lketi	n->2	
lkets	 ->4	
lkfro	n->1	
lkgru	p->2	
lkhäl	s->9	
lklap	p->1	
lklar	a->2	
lklig	.->1	
lklin	g->1	
lknin	g->57	
lkoho	l->1	
lkoml	i->5	
lkomm	a->1	e->10	
lkomn	a->42	
lkomr	ö->6	
lkoms	t->3	
lkons	t->1	
lkonv	e->1	
lkor 	-->1	a->1	f->16	h->1	i->1	o->1	s->4	t->1	u->1	v->1	ä->1	
lkor,	 ->5	
lkor.	D->3	E->1	G->1	T->1	Ö->1	
lkora	n->1	
lkore	n->21	
lkorl	i->2	
lkpar	t->10	
lkreg	e->1	
lkrep	u->3	
lkret	s->4	
lkrit	i->1	
lkrät	t->1	
lks f	r->1	
lks s	o->1	u->1	
lksty	r->1	
lkswa	g->1	
lksäg	n->1	
lkurs	e->1	
lkval	d->2	
lkvot	 ->1	
lkyrk	o->1	
lkänd	a->2	
lkänn	a->9	
lkänt	 ->1	
lköpa	r->2	
ll "M	i->1	
ll - 	n->1	r->1	s->1	
ll 10	 ->1	
ll 15	 ->1	
ll 19	3->1	5->1	9->1	
ll 2 	0->1	
ll 2,	4->1	6->1	
ll 25	 ->1	
ll 3 	0->1	
ll 30	 ->1	
ll 4 	p->1	
ll 50	 ->1	
ll 7,	4->1	
ll 70	0->1	
ll 75	 ->1	
ll 77	 ->1	
ll 83	 ->1	
ll 85	 ->1	
ll 9 	m->1	
ll 91	 ->1	
ll 94	 ->1	,->1	
ll Al	b->1	
ll Ba	r->1	
ll Bo	u->2	
ll Br	y->2	
ll Ch	i->1	
ll Co	n->1	
ll Di	m->1	
ll EG	 ->1	-->2	
ll EU	 ->2	-->1	.->1	:->2	
ll Ef	t->1	
ll Eu	r->25	
ll Fr	a->3	
ll Fö	r->4	
ll Ge	n->1	
ll Gr	e->1	
ll Ir	l->1	
ll Ka	r->1	u->1	
ll Ki	n->1	r->2	
ll Ko	s->9	
ll Ku	l->1	
ll Lo	r->2	
ll Mc	N->1	
ll Mi	c->1	
ll Mo	r->2	
ll Ni	e->2	
ll OL	F->1	
ll PP	E->1	
ll Pa	l->1	t->2	
ll Pu	r->1	
ll Ra	p->1	
ll Sc	h->1	
ll So	l->3	
ll St	.->1	r->1	
ll Sy	r->1	
ll Th	e->1	
ll Ti	b->1	
ll Tr	e->1	
ll Ty	s->2	
ll Ve	r->1	
ll Wa	l->1	s->1	
ll Wi	l->1	
ll Wu	r->1	
ll ab	s->1	
ll ac	c->1	
ll ag	e->1	
ll al	d->1	l->33	
ll an	d->4	f->1	l->1	m->1	n->1	p->1	s->11	t->3	v->10	
ll ap	p->1	
ll ar	b->8	m->1	t->4	
ll at	t->275	
ll av	 ->23	g->2	k->1	l->1	m->1	s->8	t->1	v->1	
ll ba	c->1	g->1	l->1	n->2	r->11	s->1	
ll be	 ->6	d->5	f->2	g->5	h->9	k->1	m->1	r->2	s->12	t->33	v->3	
ll bi	b->2	d->3	l->2	
ll bl	i->23	o->2	
ll bo	r->3	t->3	
ll br	a->1	i->1	o->1	ä->1	ö->1	
ll bu	d->1	
ll by	g->2	
ll bä	r->3	t->2	
ll bå	d->2	
ll bö	d->1	r->11	
ll ca	 ->1	
ll ce	n->1	
ll ci	t->2	
ll da	g->1	
ll de	 ->70	b->4	c->1	f->1	l->9	m->10	n->87	r->5	s->12	t->82	
ll di	a->3	r->17	s->8	
ll do	c->2	m->2	
ll dr	a->1	i->1	y->1	
ll du	m->1	
ll dä	r->16	
ll då	 ->3	
ll ef	t->3	
ll eg	e->3	
ll ek	o->2	
ll el	l->3	
ll em	e->2	i->1	
ll en	 ->106	b->1	d->2	e->1	t->1	
ll er	 ->3	,->4	:->1	b->1	f->1	h->1	i->2	s->1	t->1	
ll et	t->31	
ll eu	r->3	
ll ex	e->45	i->1	
ll fa	l->1	m->1	s->1	t->7	
ll fe	b->1	l->2	
ll fi	c->1	n->5	s->1	
ll fl	e->1	y->2	
ll fo	n->3	r->8	
ll fr	a->9	e->2	i->3	u->1	ä->7	å->19	
ll fu	l->5	n->8	
ll fy	l->2	
ll fä	r->1	s->1	
ll få	 ->9	n->1	r->1	
ll fö	l->23	r->129	
ll ga	g->3	m->2	r->2	
ll ge	 ->10	m->8	n->12	s->2	
ll gi	s->1	
ll gl	ä->1	
ll go	d->10	
ll gr	a->7	u->12	
ll gä	l->7	r->7	
ll gå	 ->9	.->1	n->2	
ll gö	r->23	
ll ha	 ->39	.->1	m->1	n->21	r->6	v->14	
ll he	d->1	l->3	m->2	n->1	r->4	
ll hi	n->3	
ll hj	ä->5	
ll ho	n->1	p->1	
ll hu	m->1	r->4	
ll hä	n->2	r->3	
ll hå	l->2	
ll hö	g->4	r->3	
ll i 	E->1	M->1	a->3	d->8	e->1	f->5	g->1	i->1	l->2	m->4	o->1	s->1	u->1	v->4	
ll ic	k->1	
ll id	é->1	
ll in	b->1	d->3	f->7	g->3	l->5	n->2	o->3	r->5	s->5	t->48	
ll is	r->1	
ll ja	g->107	n->1	
ll jo	r->1	
ll ju	 ->4	l->1	s->1	
ll jä	m->2	
ll ka	l->1	m->3	n->5	s->1	t->1	
ll kl	a->4	
ll kn	y->1	
ll ko	l->4	m->53	n->22	r->3	
ll kr	a->1	i->3	ä->2	
ll ku	l->1	n->56	
ll kv	e->1	
ll kä	r->2	
ll kö	k->1	
ll la	g->1	n->2	
ll le	d->5	
ll li	g->5	k->2	v->5	
ll lu	c->1	
ll ly	c->3	d->1	f->1	s->2	
ll lä	g->4	m->6	r->1	s->1	
ll lå	t->3	
ll lö	s->1	
ll ma	j->2	k->4	n->11	r->3	
ll me	d->24	l->2	n->1	r->2	t->1	
ll mi	d->1	g->3	l->1	n->17	s->1	t->2	
ll mo	b->1	t->4	
ll mu	s->1	
ll my	c->4	n->3	
ll mä	r->1	
ll må	l->3	n->4	s->3	
ll mö	j->3	t->2	
ll na	c->4	t->10	
ll ni	 ->3	v->7	
ll no	r->1	
ll nu	 ->3	
ll ny	 ->2	a->3	l->1	t->5	
ll nä	m->4	r->5	s->4	
ll nå	 ->1	g->10	
ll nö	d->2	
ll oa	c->1	
ll oc	h->45	k->26	
ll oe	n->1	
ll of	f->2	
ll oi	g->1	
ll oj	ä->1	
ll ol	i->3	y->3	
ll om	 ->6	f->9	l->1	r->4	s->2	v->1	
ll op	t->1	
ll or	d->2	g->2	o->3	ä->1	
ll os	s->4	
ll oä	n->2	
ll pa	r->9	s->1	
ll pe	n->3	r->5	
ll pi	l->1	
ll pl	a->2	
ll po	l->5	
ll pr	e->6	i->5	o->8	
ll pu	n->2	
ll på	 ->4	l->1	m->1	p->3	s->2	t->1	v->1	
ll ra	m->1	t->1	
ll re	d->3	f->1	g->12	k->3	p->1	s->11	v->2	
ll ri	k->4	s->1	
ll ro	l->1	
ll ry	m->1	
ll rä	c->3	k->1	t->16	
ll rå	d->20	
ll rö	r->1	s->1	
ll sa	k->2	m->9	n->1	t->1	
ll se	 ->15	s->2	
ll si	g->3	m->1	n->13	s->12	t->6	
ll sj	ä->2	ö->4	
ll sk	a->11	e->4	i->5	j->2	o->3	r->1	u->3	y->7	ö->2	
ll sl	u->15	å->2	
ll sm	å->2	
ll sn	a->1	
ll so	c->2	l->2	m->30	
ll sp	e->3	ä->1	
ll st	a->4	i->1	o->13	r->5	y->1	ä->4	å->42	ö->3	
ll su	b->4	s->1	v->1	
ll sv	a->2	
ll sy	n->1	s->5	
ll sä	g->39	k->4	n->2	r->4	
ll så	 ->3	d->2	
ll sö	r->1	
ll ta	 ->17	c->21	l->12	s->3	
ll te	n->1	r->1	x->1	
ll ti	d->3	l->16	t->2	
ll to	l->1	t->1	
ll tr	a->2	e->4	o->5	ä->3	
ll tu	r->1	
ll tv	i->1	ä->1	å->6	
ll ty	c->1	d->1	
ll tä	c->1	n->1	
ll u-	l->1	
ll un	d->11	i->3	
ll up	p->19	
ll ur	s->1	v->1	
ll ut	a->3	b->2	f->4	g->3	n->1	o->1	r->2	s->5	t->7	v->7	ö->2	
ll va	d->10	l->1	p->1	r->43	
ll ve	r->12	t->6	
ll vi	 ->40	c->1	d->9	k->1	l->6	s->10	
ll vo	l->1	r->2	
ll vä	g->1	l->2	n->2	r->1	s->1	
ll vå	r->15	
ll yr	k->2	
ll yt	t->3	
ll Ös	t->1	
ll äg	n->1	
ll än	 ->6	d->12	
ll är	 ->12	?->1	
ll äv	e->5	
ll åk	l->1	
ll år	 ->2	
ll ås	t->2	
ll åt	a->2	e->12	g->3	s->1	t->1	
ll ök	a->5	n->1	
ll ön	s->1	
ll öp	p->3	
ll ös	t->1	
ll öv	e->15	
ll!He	r->1	
ll!Ja	g->1	
ll", 	s->1	v->1	
ll".I	 ->1	
ll, a	t->2	v->1	
ll, b	e->1	
ll, d	e->1	v->1	ä->1	
ll, e	f->1	r->1	u->1	
ll, f	r->1	ö->2	
ll, h	a->1	u->1	ä->1	
ll, i	 ->4	
ll, j	a->1	u->1	
ll, k	a->1	
ll, m	e->7	o->1	
ll, n	a->1	ä->2	å->1	
ll, o	c->12	
ll, p	å->1	
ll, r	ö->1	
ll, s	o->5	å->2	ö->1	
ll, t	o->1	
ll, u	n->1	t->2	
ll, v	a->3	i->2	
ll, ä	n->1	v->2	
ll, å	t->2	
ll- o	c->4	
ll. D	e->1	
ll. o	c->1	
ll.An	g->1	
ll.Av	s->1	
ll.Bi	l->1	
ll.De	 ->1	n->2	t->18	
ll.Dä	r->1	
ll.En	l->2	
ll.Et	t->1	
ll.Fi	n->2	
ll.Fr	å->1	
ll.Fö	r->2	
ll.Ha	r->1	
ll.He	r->3	
ll.Hä	r->1	
ll.I 	A->1	d->1	f->1	o->1	
ll.In	t->1	
ll.Ja	g->11	
ll.Ko	m->2	s->1	
ll.Me	d->1	n->1	
ll.Må	l->1	
ll.Om	 ->1	
ll.Or	k->1	
ll.Pr	o->1	
ll.På	 ->1	
ll.Re	s->1	
ll.Sa	n->1	
ll.Sm	å->1	
ll.So	m->1	
ll.Så	 ->1	s->1	
ll.Ta	n->1	
ll.Tä	n->1	
ll.Ut	m->1	
ll.Vi	 ->8	
ll.Vo	n->1	
ll.Vå	r->1	
ll.Än	 ->1	
ll: "	h->1	
ll: e	n->1	
ll: j	a->1	
ll?. 	(->1	
ll?Da	g->1	
ll?Hu	r->1	
ll?Ja	g->1	
ll?Ko	l->1	
lla -	 ->1	
lla A	l->1	
lla E	U->2	u->2	
lla F	ö->1	
lla H	i->1	
lla P	a->1	
lla a	g->1	k->1	l->3	n->15	r->3	s->7	t->25	v->6	
lla b	a->2	e->21	i->7	l->1	o->4	r->1	u->1	ö->2	
lla d	e->94	i->9	o->6	r->1	
lla e	f->1	g->2	k->1	l->4	m->2	n->16	r->7	t->4	u->6	v->2	
lla f	a->17	i->3	l->1	o->11	r->23	å->2	ö->27	
lla g	e->2	l->1	o->3	r->8	
lla h	a->15	i->1	j->2	o->3	u->3	ä->1	å->1	ö->5	
lla i	 ->5	d->1	n->25	s->1	
lla j	o->3	u->2	ä->1	
lla k	a->8	l->3	n->2	o->25	r->6	v->2	ä->1	
lla l	a->6	e->2	i->3	o->1	ä->6	ö->2	
lla m	a->5	e->30	i->7	o->2	u->1	y->17	ä->2	å->2	ö->3	
lla n	e->2	i->9	o->1	u->1	y->1	ä->2	å->1	ö->1	
lla o	c->22	d->1	l->4	m->20	r->4	s->4	
lla p	a->15	e->2	l->1	o->13	r->12	u->1	å->3	
lla r	a->4	e->27	i->3	o->1	ä->14	ö->1	
lla s	a->7	e->2	i->21	j->4	k->8	l->4	o->15	p->3	t->22	u->1	v->1	y->5	ä->4	å->3	
lla t	a->3	e->2	i->8	j->9	o->3	r->8	y->1	ä->1	
lla u	n->3	p->8	t->12	
lla v	a->6	e->8	i->6	ä->4	å->7	
lla ä	n->3	r->2	
lla å	k->2	r->1	s->1	t->6	
lla ö	n->1	p->1	v->3	
lla!H	e->1	
lla, 	f->1	h->1	i->2	k->1	m->1	n->1	o->2	p->1	r->1	s->2	
lla.D	e->5	ä->1	
lla.H	e->1	
lla.J	a->1	
lla.V	i->2	
lla:F	ö->1	
llad 	e->1	m->1	p->1	r->1	s->1	
llade	 ->4	s->1	
llamt	 ->1	
llan 	1->5	8->2	C->2	D->1	E->10	G->1	H->1	I->9	P->3	S->3	a->5	b->2	c->1	d->31	e->7	f->10	g->2	h->2	i->1	k->17	l->6	m->14	n->4	o->5	p->8	r->18	s->10	t->2	u->5	v->5	Ö->1	ä->1	
llan"	 ->1	
llan,	 ->3	
llan.	E->1	I->1	
lland	e->145	
llanl	i->1	
llann	i->1	
llans	t->7	
llant	e->1	i->1	
llanö	s->19	
llar 	"->1	a->1	d->5	f->1	i->1	l->1	o->1	p->2	s->3	
llar,	 ->3	
llar.	K->1	
llar;	 ->1	
llare	 ->1	,->1	n->3	
llarn	 ->2	a->2	
llas 	a->3	d->1	e->7	i->4	k->1	m->2	n->2	o->4	p->3	s->1	t->3	u->6	v->3	ö->1	
llas,	 ->4	
llas.	D->1	K->1	
llast	e->1	
llat 	"->2	d->2	n->1	
llava	r->1	
llbak	a->51	s->1	
llbar	 ->19	a->1	h->1	t->5	
llbes	t->1	
llbil	d->1	
llbor	d->3	
llbri	n->4	
lld a	v->1	
lld b	o->1	
lld p	a->1	å->1	
lld t	i->1	
llda 	f->1	i->1	m->3	o->1	s->1	t->3	v->1	
llda,	 ->4	
llda.	D->1	E->1	H->1	J->2	Ä->1	
lldas	 ->2	
llde 	B->1	K->1	a->1	d->5	e->2	f->4	h->1	n->2	o->1	t->1	u->1	å->1	
lldel	a->10	e->23	n->3	
lldes	 ->8	.->1	
lldhe	t->23	
lldra	g->1	
lle -	 ->1	
lle E	u->3	
lle K	i->1	
lle a	l->3	n->3	t->18	v->1	
lle b	a->3	e->9	i->1	l->5	ö->2	
lle d	e->28	o->3	ä->8	å->2	
lle e	l->1	m->1	n->5	v->1	
lle f	a->1	i->2	r->4	å->4	ö->20	
lle g	e->2	o->1	r->1	ä->7	å->1	ö->5	
lle h	a->18	e->1	ä->4	
lle i	 ->6	n->20	
lle j	a->44	
lle k	a->1	o->6	r->2	u->56	ä->1	
lle l	e->4	ä->1	
lle m	a->2	e->2	o->1	
lle n	a->1	i->1	u->1	ä->1	
lle o	c->10	f->1	l->1	
lle p	a->2	l->1	å->2	
lle r	e->2	ä->1	å->1	ö->1	
lle s	a->1	e->1	j->1	k->5	l->2	o->4	p->1	t->3	v->1	ä->4	å->6	ö->1	
lle t	.->1	a->5	i->5	r->1	v->2	
lle u	n->3	p->4	r->3	t->6	
lle v	a->37	e->2	i->81	ä->3	
lle ä	n->1	r->1	v->1	
lle å	t->2	
lle ö	n->2	
lle, 	o->3	
lle.J	a->1	
llega	 ->36	!->4	,->3	.->1	l->9	n->16	s->2	
llege	r->127	
llegi	e->2	u->2	
llego	r->4	
lleha	n->3	
llekt	i->10	u->3	
llele	r->3	
llell	a->2	t->3	
llels	e->9	
llen 	a->7	b->2	d->3	e->1	f->5	g->1	h->3	i->12	k->3	m->1	o->7	p->1	s->10	t->1	u->3	v->1	ä->1	å->2	ö->1	
llen"	 ->1	
llen,	 ->10	
llen.	A->1	D->4	E->1	H->2	I->1	J->2	K->1	M->3	R->1	S->1	T->1	V->1	
llena	 ->4	,->1	r->1	
llenn	i->7	
llens	 ->2	
llenÄ	r->1	
ller 	-->3	2->1	7->1	8->1	9->1	A->3	D->1	E->8	F->4	I->1	J->1	L->1	M->1	N->1	P->2	R->2	S->4	T->3	U->2	a->71	b->26	c->2	d->112	e->66	f->88	g->22	h->20	i->67	j->5	k->41	l->21	m->61	n->18	o->46	p->36	r->16	s->71	t->28	u->20	v->36	Ö->2	ä->14	å->8	ö->7	
ller,	 ->6	
ller.	D->1	F->1	H->2	J->2	M->1	O->1	R->1	Ä->1	
ller;	 ->1	
llera	 ->18	d->3	r->3	s->9	t->2	
llerk	ä->3	
llern	a->5	
llert	i->67	
lles 	a->1	h->1	i->1	j->1	r->1	s->1	
llesa	m->5	
llet 	-->1	A->1	V->1	a->7	b->3	d->2	e->2	f->34	g->2	h->9	i->23	j->1	k->2	l->1	m->3	n->1	o->13	r->4	s->8	t->8	u->1	v->4	Ö->1	ä->4	ö->1	
llet!	P->1	
llet,	 ->17	
llet.	 ->1	)->1	A->1	D->8	I->1	J->5	K->1	N->1	O->1	S->2	T->1	U->1	V->4	
llet:	 ->1	
llets	 ->3	
lleur	o->2	
llfin	g->1	
llfog	a->6	
llfre	d->27	
llfun	k->1	
llfäl	l->97	
llfär	d->1	
llföl	j->3	
llför	 ->3	.->1	a->2	b->3	l->4	s->3	v->1	
llgjo	r->1	
llgod	o->1	
llgri	p->2	
llgän	g->21	
llgån	g->25	
llgåv	o->1	
llgör	a->1	
llhan	d->43	
llhet	 ->1	,->2	
llhör	 ->4	a->3	i->1	
lli h	a->1	
lli!J	a->1	
llian	s->7	
llibe	r->1	
llier	a->1	
llig 	a->1	f->1	i->1	n->1	o->1	p->1	u->2	v->1	
lliga	 ->16	,->2	.->1	r->3	
llige	n->5	
lligh	e->25	
lligs	e->1	
lligt	 ->24	,->1	.->1	
lliho	p->1	
llind	u->1	
lling	 ->1	
llise	r->2	
llisi	o->3	
llit 	-->1	a->2	b->1	e->3	f->2	h->1	i->1	m->1	o->2	p->1	s->4	t->1	ö->1	
llit,	 ->1	
llite	t->1	
llits	 ->4	.->2	
llive	t->1	
llkas	t->1	
llkla	r->2	
llkom	l->5	m->4	s->2	
llkor	 ->29	,->4	.->7	a->1	e->21	l->2	
llkän	n->9	
llmak	t->1	
llmos	o->1	
llmyn	d->2	
llmän	 ->18	g->1	h->47	n->42	t->17	
llmär	k->1	
llmät	a->1	e->1	
llmöj	l->2	
llmös	s->1	
llmöt	e->3	
llna,	 ->1	
llnad	 ->10	:->1	e->33	
llnin	g->140	
llnis	c->1	
llnär	m->6	
llo g	o->1	
llo i	 ->1	
llo o	c->1	
llo r	e->1	
llo å	t->1	
llobb	y->2	
lloja	l->2	
lloke	r->1	
llolj	a->1	
llomr	å->1	
llor 	f->2	h->2	i->2	k->1	m->1	o->4	s->1	t->1	v->2	ä->2	
llor,	 ->5	
llor.	D->4	F->1	H->1	J->1	M->2	O->1	V->1	Ä->1	
llorg	a->1	
llorn	a->5	
llpol	i->1	
llra 	b->2	f->1	h->1	s->3	v->2	
llran	d->1	
llre 	H->1	a->1	b->1	h->1	s->1	v->1	
llrin	g->1	
llris	k->1	
llräc	k->75	
llrät	t->6	
lls C	E->1	
lls a	l->2	n->2	t->1	v->2	
lls b	e->2	l->1	
lls d	e->3	r->1	
lls e	n->1	
lls f	u->1	
lls h	a->11	u->1	ä->1	
lls i	 ->7	n->10	
lls k	u->1	
lls m	e->2	
lls n	å->1	
lls o	c->1	l->1	
lls p	å->5	
lls s	a->2	k->3	o->2	
lls t	i->2	r->1	v->1	
lls u	t->3	
lls v	a->3	i->3	ä->1	
lls ä	n->1	r->2	
lls å	s->1	t->1	
lls ö	v->1	
lls, 	f->1	g->1	o->1	p->1	
lls.D	e->3	
lls.F	ö->1	
lls.H	a->1	
lls.N	u->1	
lls.T	a->1	
lls.U	n->1	
lls.Y	t->1	
lls?V	i->1	
llsam	h->1	m->31	
llsat	s->1	t->2	
llsbe	d->1	
llse 	a->13	
llsek	o->3	
llsfö	r->1	
llsha	n->1	
llsid	i->1	
llska	p->9	
llsko	t->1	
llskr	i->2	
llskt	.->1	
llsky	n->1	
llsli	g->1	
llslu	t->1	
llslö	s->1	
llsme	d->1	
llsmä	n->1	s->2	
llsom	g->1	
llsri	k->2	
llsse	r->1	
llsst	r->3	
llsti	l->7	
llsto	l->3	
llstr	ö->4	
llstu	d->1	
llstä	n->41	
llstå	n->22	
llsva	r->3	
llsvi	l->1	
llsvä	r->1	
llsyn	t->2	
llsys	t->3	
llsäm	n->1	
llsät	t->4	
llt -	 ->1	
llt 1	8->1	
llt a	n->9	t->10	v->4	
llt b	e->4	i->1	l->2	o->1	u->1	ä->1	ö->2	
llt d	e->39	o->1	r->1	ä->1	
llt e	f->1	k->1	n->2	r->1	t->1	
llt f	a->2	e->1	i->5	l->2	o->1	r->3	ö->24	
llt g	e->3	i->1	o->2	y->1	ä->1	
llt h	a->1	ä->1	
llt i	 ->13	n->15	
llt k	a->4	o->11	r->1	u->2	ä->1	
llt l	ä->1	
llt m	e->12	i->3	o->1	å->1	
llt n	a->1	ä->4	å->1	ö->1	
llt o	c->11	f->2	m->3	r->1	s->2	
llt p	a->1	l->1	o->2	r->2	å->7	
llt r	e->2	i->2	
llt s	a->10	e->9	i->3	j->1	k->6	o->7	t->12	v->2	y->1	ä->3	å->1	ö->1	
llt t	i->4	r->2	v->1	
llt u	n->4	p->2	r->1	t->13	
llt v	a->3	i->5	ä->5	å->2	
llt y	t->1	
llt ä	n->2	r->7	
llt å	t->1	
llt ö	p->1	v->2	
llt, 	a->1	b->2	d->1	e->1	f->1	j->1	m->1	o->3	s->1	t->1	u->1	v->2	ä->1	
llt.D	e->5	
llt.H	e->1	
llt.M	a->1	e->1	
llt.V	i->2	
llt: 	a->1	
llt; 	d->1	
llta 	ä->1	
lltag	a->1	
lltal	a->1	
lltfl	e->1	
lltfö	r->39	
lltid	 ->74	,->2	.->1	
lltih	o->1	
lltin	g->5	
lltjä	m->3	
lltme	r->1	
lltro	 ->1	
llträ	d->7	
llts 	-->1	a->1	f->1	i->2	m->1	o->1	t->1	ä->1	
llts:	 ->1	
lltsa	m->1	
lltse	d->3	
lltså	 ->61	,->2	
lluti	o->1	
lluts	k->14	
llval	.->1	
llvar	 ->6	,->1	.->4	e->1	l->62	
llver	k->87	
llvid	a->1	
llvil	l->1	
llväg	a->8	
llvän	t->1	
llvär	d->2	
llväx	t->20	
lly f	ö->1	
lly! 	G->1	
lly.A	n->1	
llybe	t->1	
llys 	b->1	
llywo	o->1	
llägg	 ->6	,->1	a->8	s->3	
llägn	a->2	
llämp	a->99	l->11	n->67	
lländ	a->2	
llång	 ->4	
llåt 	m->10	
llåta	 ->8	s->5	
llåte	n->3	r->16	t->1	
llåtl	i->3	
llåtn	a->6	
llåts	 ->3	
llösa	 ->1	
llösn	i->1	
lm de	n->1	
lm, h	a->1	
lm.He	r->1	
lmajo	r->1	
lmakt	e->1	
lman 	F->1	I->2	f->1	o->3	
lman!	 ->224	A->1	D->2	E->2	J->6	M->1	S->1	T->2	U->1	V->2	
lman,	 ->157	
lman:	 ->1	
lmann	e->11	
lmans	k->9	
lmar 	B->2	
lmast	e->1	
lmede	l->2	
lmedv	e->1	
lmen 	C->1	
lment	 ->1	a->1	
lmer 	o->1	
lmoso	r->1	
lmsha	v->1	
lmynd	i->2	
lmän 	a->1	d->2	f->2	g->2	o->2	p->1	r->2	å->6	
lmäng	i->1	
lmänh	e->47	
lmänn	a->39	e->1	y->2	
lmänt	 ->16	,->1	
lmärk	e->2	
lmäss	i->2	
lmäta	s->1	
lmäte	r->1	
lmåen	d->2	
lmöjl	i->2	
lmöss	o->1	
lmöte	s->3	
ln "u	t->1	
ln at	t->1	
ln fö	r->3	
ln i 	d->1	f->1	
ln ko	n->1	
ln me	d->1	
ln oc	h->2	
ln om	 ->1	
ln ti	l->5	
ln är	 ->2	
ln, d	ä->1	
ln, h	a->1	
ln.De	t->1	
lna k	o->1	
lna, 	m->1	
lnad 	b->1	f->2	i->2	m->4	s->1	
lnad:	 ->1	
lnade	n->3	r->30	
lning	 ->72	,->7	.->19	?->1	a->17	e->41	s->55	
lnisc	h->1	
lns l	a->2	
lnärm	e->1	n->5	
lo go	d->1	
lo gå	n->1	
lo i 	d->1	
lo må	l->1	
lo oc	h->3	
lo re	s->1	
lo åt	e->1	
lo, W	y->1	
lo, s	e->1	o->1	
loakl	u->1	
lobal	 ->1	a->4	i->5	t->2	
lobby	a->1	g->2	i->2	m->1	n->3	v->1	
locka	 ->2	d->2	n->2	
lockb	i->1	
locke	r->2	t->1	
lod t	a->1	ä->1	
loden	 ->2	
lodla	r->1	
log a	t->1	v->1	
log b	e->2	
log e	n->1	r->1	t->1	
log f	a->1	
log i	 ->3	
log m	e->9	å->1	
log o	m->1	
log s	o->4	t->1	
log t	i->1	
log v	i->1	
log ä	r->1	
log å	t->1	
log, 	o->1	v->1	
log.D	a->1	
log.F	r->1	ö->1	
log.H	a->1	
log.J	a->2	
log.N	ä->1	
loge 	f->1	
loge,	 ->1	
logen	 ->7	.->1	
logi 	-->1	o->2	
logik	 ->1	,->2	.->3	e->2	
login	,->1	
logis	k->33	
logs 	a->1	i->1	p->1	t->1	
lojal	a->2	i->5	
lok o	c->1	
loka 	h->1	
lokal	 ->7	a->31	i->3	p->1	t->2	
lokas	t->1	
loker	i->1	
lokt 	d->2	s->2	v->1	
lolad	d->1	
lolja	,->1	
lomat	e->1	i->10	
lomet	e->1	
lomma	.->1	
lommo	r->2	
lområ	d->1	
lomst	r->3	
lomäs	s->1	
lonap	r->2	
lonia	l->1	
lonmä	s->1	
looij	-->1	
lopp 	-->1	a->2	h->2	i->1	s->1	
lopp,	 ->1	
lopp.	.->1	
loppe	n->4	t->8	
lor f	r->1	ö->1	
lor h	a->3	
lor i	n->2	
lor k	a->1	
lor m	e->2	
lor o	c->6	m->1	
lor s	a->1	å->1	
lor t	i->2	
lor v	i->2	
lor ä	r->2	
lor, 	b->1	e->1	i->1	o->1	s->2	
lor.D	e->3	ä->1	
lor.F	r->1	
lor.H	u->1	
lor.J	a->2	
lor.M	e->2	
lor.O	c->1	
lor.V	i->1	
lor.Ä	v->1	
lora 	1->1	i->1	o->1	s->1	
lorad	 ->2	e->3	
lorar	 ->4	
lorat	 ->4	,->1	.->2	s->1	
loren	z->19	
lorga	n->1	
lorna	 ->3	,->1	s->1	
lors 	b->1	h->1	
lors.	V->1	
los f	ö->1	
los o	c->4	
losio	n->1	
losiv	 ->1	
losof	i->5	
loss 	d->1	
lossa	l->1	
lossn	i->1	
lot i	 ->1	
loten	 ->1	
lotpr	o->2	
lott 	h->1	o->1	
lotta	 ->2	,->1	d->3	n->1	s->1	
lotto	r->1	
lotts	p->1	
lov a	t->1	
lov i	n->1	
lova 	a->2	
lovad	e->4	
lovak	i->1	
lovar	 ->1	
lovat	 ->5	.->1	s->1	
loven	s->1	
lovo 	o->1	
lovor	d->2	
lovvä	r->2	
lovyt	t->1	
loyds	 ->1	
lp at	t->1	
lp av	 ->26	
lp de	 ->1	
lp fr	å->3	
lp fö	r->3	
lp ni	 ->1	
lp oc	h->2	
lp på	 ->1	
lp sk	a->1	
lp so	m->1	
lp ti	l->5	
lp vi	d->2	
lp öv	e->1	
lp, d	å->1	
lp, m	e->1	
lp.De	t->1	
lp.Hä	r->1	
lp.I 	a->1	
lp.Ja	g->1	
lp.Vi	 ->1	
lpa W	a->1	
lpa a	n->1	
lpa d	e->5	
lpa f	ö->2	
lpa g	e->1	
lpa h	o->1	
lpa i	n->1	
lpa k	o->2	
lpa l	a->1	
lpa m	e->2	i->1	ä->4	ö->1	
lpa o	f->2	s->1	
lpa p	e->1	
lpa s	o->1	å->1	
lpa t	i->7	
lpa v	å->1	
lpand	e->3	
lpare	 ->1	
lpark	 ->2	e->4	
lparl	a->1	
lpatr	i->1	
lpe p	å->1	
lpen 	i->1	s->1	ä->2	
lper 	d->1	
lpern	a->1	
lpes 	e->1	
lplan	.->1	
lplig	t->1	
lpoli	s->1	t->44	
lprob	l->1	
lprod	u->2	
lprog	r->1	
lps.J	u->1	
lpt t	i->1	
lpta.	D->1	
lpte 	t->1	
lpunk	t->2	
lpvil	l->1	
lra b	ä->2	
lra f	l->1	
lra h	ö->1	
lra s	e->2	t->1	
lra v	i->1	ä->1	
lrand	e->1	
lrapp	o->1	
lre H	i->1	
lre a	t->1	
lre b	ö->1	
lre h	a->1	
lre s	e->1	
lre v	e->1	
lrege	r->1	
lregl	e->4	
lresu	l->1	r->3	
lrika	 ->4	
lrikt	a->1	
lring	e->1	
lrisk	,->1	
lroll	,->1	
lrum 	f->1	
lryck	n->1	
lräck	l->75	
lräke	n->1	
lräkn	i->1	
lrätt	 ->3	a->3	e->4	s->1	
ls CE	N->1	
ls al	k->1	l->2	
ls an	s->1	t->1	
ls ar	b->3	
ls at	t->4	
ls av	 ->4	s->1	
ls ba	r->1	
ls be	f->1	n->1	
ls bl	i->1	
ls de	 ->1	n->1	t->1	
ls dr	a->1	
ls dä	r->1	
ls en	 ->1	
ls ex	i->1	
ls fa	l->1	m->1	
ls fi	s->1	
ls fr	i->1	
ls fu	l->1	
ls fö	r->3	
ls ga	l->1	
ls ha	f->1	r->10	
ls he	k->1	
ls hu	r->1	
ls hä	r->1	
ls i 	a->3	d->2	f->1	n->1	
ls il	l->1	
ls in	f->1	g->2	i->2	t->7	
ls ko	m->1	
ls ku	n->1	
ls kv	i->1	
ls li	v->2	
ls me	d->2	s->1	
ls mi	l->3	
ls mä	n->2	
ls må	n->1	
ls nå	g->1	
ls oc	h->3	k->1	
ls ol	i->1	
ls or	d->2	
ls pr	e->2	i->1	o->1	
ls på	 ->5	
ls sa	m->1	t->1	
ls se	m->1	
ls sk	a->3	u->1	
ls so	l->1	m->2	
ls st	ö->1	
ls ti	l->6	
ls tr	o->1	
ls tv	i->1	
ls up	p->1	
ls ut	,->3	
ls va	r->3	t->1	
ls vi	 ->1	d->2	
ls vä	g->2	
ls än	n->1	
ls är	 ->2	
ls år	 ->1	.->1	
ls ås	t->1	
ls åt	 ->1	a->1	g->1	
ls öv	e->1	
ls, f	o->1	
ls, g	e->1	
ls, o	c->1	
ls, p	å->1	
ls- o	c->1	
ls.De	n->1	t->3	
ls.Fö	r->1	
ls.Ha	n->1	
ls.Nu	 ->1	
ls.Ta	n->1	
ls.Un	d->1	
ls.Yt	t->1	
ls?Vi	l->1	
lsa k	o->1	
lsa o	c->11	
lsa p	å->1	
lsa s	t->1	
lsa t	i->1	
lsa, 	d->2	e->1	
lsa.H	e->1	
lsace	 ->1	.->2	
lsamh	e->1	
lsamm	a->31	
lsan 	h->1	
lsan,	 ->2	
lsan.	S->1	
lsar 	k->1	
lsats	e->1	
lsatt	a->1	e->1	s->1	
lsavg	ö->1	
lsbed	r->1	
lsbur	n->1	
lsdom	s->1	
lsdrä	n->1	
lse -	 ->3	
lse a	t->16	v->11	
lse b	e->1	
lse d	e->2	
lse e	l->1	
lse f	r->1	ö->15	
lse g	e->2	i->1	
lse h	a->3	
lse i	 ->3	n->2	
lse j	a->2	u->1	
lse k	a->2	o->3	
lse m	e->14	o->1	
lse n	o->2	ä->2	
lse o	c->12	m->5	
lse p	å->2	
lse r	e->1	
lse s	k->1	o->16	t->1	ä->1	å->1	
lse t	i->2	
lse u	n->1	
lse v	i->1	
lse ä	r->3	
lse ö	v->4	
lse, 	d->1	e->2	i->2	j->1	k->1	m->3	t->1	u->1	
lse- 	o->1	
lse.B	e->1	
lse.D	e->5	
lse.E	f->1	t->1	
lse.J	a->3	
lse.K	o->1	
lse.L	å->1	
lse.M	e->1	i->1	
lse.N	i->1	
lse.S	a->1	k->1	
lse.V	i->2	
lseak	t->1	
lseby	g->1	
lsefu	l->11	
lsehi	n->1	
lseko	n->5	
lsekr	e->2	
lsekt	o->6	
lsele	d->2	
lselö	s->3	
lsemö	n->1	
lsen 	-->1	1->1	a->20	f->5	h->1	i->2	k->1	m->2	o->3	s->1	t->1	v->2	ä->1	
lsen,	 ->3	
lsen.	A->1	G->1	J->1	N->1	Ä->1	
lsenl	i->2	
lsens	 ->4	
lseom	r->1	
lser 	-->2	a->4	b->1	e->3	f->12	g->3	h->2	i->4	k->2	m->4	n->1	o->12	p->3	s->26	t->5	u->2	ä->2	
lser!	D->1	
lser,	 ->19	
lser.	B->1	D->5	I->2	K->2	S->1	T->1	V->1	
lser:	 ->1	
lseri	k->1	
lsern	a->52	
lsers	 ->1	
lseut	v->1	
lsevi	s->2	
lsexp	o->1	
lsfal	l->1	
lsfas	e->1	
lsflo	t->2	
lsfrå	g->2	
lsför	h->1	s->1	
lshan	t->2	
lshin	d->1	
lsidi	g->1	
lsign	e->1	
lsike	.->1	
lsind	u->2	
lsing	f->20	
lsitu	a->1	
lsk-f	r->1	
lska 	"->1	d->1	g->1	i->1	k->2	l->1	m->1	n->1	o->1	s->1	v->3	
lska.	J->1	
lska:	 ->1	
lskan	d->2	
lskap	.->1	a->1	e->6	l->1	
lskar	 ->1	
lskat	t->3	
lsken	 ->1	
lskif	t->1	
lskni	n->1	
lskom	m->1	
lskon	s->1	t->1	
lskot	t->1	
lskri	s->2	v->2	
lskro	t->2	v->2	
lskt 	e->1	l->1	
lskt.	J->1	
lskul	t->1	
lskva	l->1	
lskyd	d->4	
lskyn	d->1	
lsköp	a->1	
lslag	s->5	
lslig	a->1	
lslog	i->1	
lslut	a->1	
lslös	n->1	t->1	
lsmed	b->1	
lsmyn	d->9	
lsmän	 ->1	g->1	
lsmäs	s->4	
lsnin	g->2	
lsnyh	e->1	
lso- 	o->1	
lsoci	a->1	
lsoef	f->1	
lsomg	i->1	
lsomr	å->2	
lson 	k->1	o->1	s->1	v->1	
lson.	N->1	
lsore	l->1	
lsorg	a->3	
lsori	s->1	
lsosk	y->1	
lsovå	d->1	r->2	
lspar	t->1	
lspla	t->2	
lspol	i->2	
lspri	s->1	
lspro	c->1	d->1	g->1	
lspun	k->6	
lsrik	a->2	
lsruh	e->2	
lsrun	d->1	
lssek	t->1	
lsser	v->1	
lssid	a->1	
lssjö	f->1	
lssti	l->1	
lsstr	ö->3	
lsstö	d->1	
lssys	t->1	
lssäk	e->43	
lst a	n->1	t->1	
lst b	e->1	
lst f	ö->1	
lst h	a->1	
lst i	 ->1	l->1	n->4	
lst k	o->1	
lst l	a->1	
lst m	o->1	å->2	
lst n	o->1	
lst p	r->1	å->1	
lst r	e->1	
lst s	e->2	k->3	o->1	y->1	
lst t	v->2	
lst u	t->1	
lst v	a->1	i->3	
lst ä	r->1	
lst, 	d->2	e->2	f->1	h->1	i->1	
lst. 	A->1	
lst.A	c->1	
lst.D	e->1	
lst.F	ö->1	
lst.V	i->1	
lstat	e->5	s->2	
lster	 ->1	
lstho	m->3	
lstil	l->9	
lstol	 ->1	e->1	p->1	s->1	
lstor	 ->1	,->1	a->38	t->1	
lstru	k->1	
lströ	m->4	
lstud	i->1	
lstvi	s->1	
lstän	d->41	
lstån	d->28	
lstöd	 ->1	e->1	
lsumm	a->1	
lsuta	n->3	
lsuts	l->1	
lsvar	a->4	
lsvil	l->1	
lsvär	d->1	
lsväs	e->1	
lsyn.	E->1	
lsynt	 ->2	
lsyst	e->6	
lsämn	e->1	
lsätt	a->2	e->1	n->120	
lsöka	n->6	
lt - 	e->1	s->1	
lt 18	0->1	
lt 27	 ->1	
lt 70	0->1	
lt 95	 ->1	
lt EU	 ->1	-->2	.->1	
lt St	o->1	
lt Su	d->1	
lt ab	s->1	
lt ad	m->1	
lt ak	t->1	
lt al	l->1	
lt an	g->1	n->3	s->8	t->1	v->1	
lt ar	b->1	
lt at	t->22	
lt av	 ->3	s->2	t->1	
lt be	 ->1	f->1	h->2	k->1	r->2	t->5	
lt bi	d->1	
lt bl	a->1	i->1	
lt bo	r->1	
lt br	a->1	
lt bu	d->2	
lt bä	t->1	
lt bö	r->3	
lt de	 ->11	b->1	l->1	m->1	n->2	t->32	
lt di	r->1	
lt do	k->1	
lt dr	a->2	
lt dä	r->2	
lt ef	t->3	
lt ek	o->1	
lt el	l->1	
lt en	 ->2	d->1	i->2	k->19	s->1	
lt er	 ->1	k->1	
lt et	t->5	
lt fa	l->2	r->2	
lt fe	l->1	
lt fi	n->5	s->1	
lt fl	e->3	
lt fo	r->1	
lt fr	a->2	e->1	u->1	å->3	
lt fä	s->1	
lt få	g->1	
lt fö	r->42	
lt ge	m->1	n->4	
lt gi	c->1	
lt gl	a->1	
lt go	d->5	
lt gy	n->1	
lt gä	l->3	
lt ha	n->6	r->3	
lt he	r->1	
lt hä	n->2	
lt i 	E->4	F->2	K->1	a->1	d->5	e->2	l->4	o->1	s->6	t->2	u->1	v->2	ö->2	
lt il	l->1	
lt im	p->1	
lt in	f->4	o->3	s->2	t->14	v->1	
lt jo	r->1	
lt ju	r->1	
lt ka	m->1	n->2	p->1	
lt kl	a->16	
lt ko	m->9	n->3	r->8	
lt kr	ä->1	
lt ku	l->1	n->1	
lt kä	n->3	r->1	
lt li	g->1	
lt lo	g->1	
lt ly	s->1	
lt lä	m->1	
lt me	d->18	l->1	n->1	r->2	
lt mi	l->1	n->1	s->2	
lt mo	n->1	t->1	
lt my	c->1	
lt mä	r->1	
lt må	n->2	s->1	
lt na	t->1	
lt no	g->1	r->1	t->1	
lt ny	 ->1	a->1	l->1	
lt nä	m->1	r->7	
lt nå	g->2	
lt nö	d->3	
lt oa	c->3	
lt oc	h->31	
lt of	t->1	ö->1	
lt ol	y->1	
lt om	 ->6	e->1	ö->1	
lt or	e->2	i->1	o->1	
lt os	s->2	y->1	
lt ot	i->1	
lt ov	ä->1	
lt pa	r->1	s->1	
lt pl	a->4	
lt po	l->1	s->1	
lt pr	o->2	ä->1	
lt pu	n->2	
lt på	 ->16	
lt ra	k->1	
lt re	d->2	
lt ri	k->6	s->1	
lt rä	t->8	
lt sa	k->2	m->9	t->1	
lt se	 ->2	d->2	t->9	
lt si	g->2	n->1	t->1	
lt sj	ä->2	
lt sk	a->3	r->1	u->3	y->1	
lt sn	a->1	
lt so	m->10	
lt sp	a->1	
lt st	a->4	o->1	ö->11	
lt sv	a->2	
lt sy	f->1	
lt sä	g->1	k->3	n->2	t->9	
lt så	d->1	
lt sö	k->1	
lt ta	c->2	
lt ti	l->16	
lt tr	e->1	y->1	ä->1	
lt tv	å->1	
lt ty	d->4	
lt un	d->4	
lt up	p->9	
lt ur	 ->1	
lt ut	 ->4	,->4	.->4	e->1	n->1	t->3	
lt va	d->5	n->2	r->1	
lt vi	a->1	d->1	k->10	l->4	s->4	
lt vä	g->1	r->1	s->3	
lt vå	r->4	
lt yt	t->1	
lt än	 ->1	d->3	
lt är	 ->7	e->1	l->1	
lt äv	e->1	
lt åt	 ->2	a->1	
lt åv	i->1	
lt öp	p->1	
lt öv	e->11	
lt, a	t->1	
lt, b	r->1	ö->1	
lt, d	e->1	
lt, e	t->1	
lt, f	ö->2	
lt, j	a->1	
lt, m	e->3	
lt, o	c->5	m->1	
lt, s	o->1	
lt, t	y->1	
lt, u	t->1	
lt, v	a->1	i->1	
lt, ä	v->1	
lt, å	t->1	
lt. D	e->1	
lt.De	l->1	t->9	
lt.En	l->1	
lt.He	r->2	
lt.Hä	r->1	
lt.I 	m->1	
lt.Ja	g->2	
lt.Ma	n->1	
lt.Me	d->1	
lt.Om	 ->1	
lt.Un	d->1	
lt.Va	d->3	
lt.Vi	 ->3	
lt: a	t->1	
lt; d	e->2	
lt?Ja	g->1	
lta f	u->1	
lta i	 ->12	n->1	
lta o	c->2	m->1	
lta p	å->2	
lta s	t->1	
lta u	t->1	
lta ä	r->1	v->1	
lta ö	v->2	
lta, 	o->2	s->1	
ltaga	n->24	r->1	
ltagi	t->6	
ltakt	i->1	
ltala	 ->1	
ltali	g->2	
ltar 	d->1	i->8	v->1	
ltare	,->1	
ltas 	a->1	
ltat 	a->5	b->1	f->2	h->1	i->5	k->1	m->1	o->2	s->8	u->2	v->2	ä->1	
ltat,	 ->6	
ltat.	 ->1	D->1	E->1	H->1	I->2	J->2	K->1	O->1	
ltat:	 ->1	
ltat?	.->1	J->1	
ltate	n->16	t->28	
ltati	n->1	o->2	
ltatl	i->1	
ltatt	a->7	
ltatö	v->6	
ltbas	i->1	
lte k	ä->1	
lte v	i->1	
lte, 	d->1	s->1	
lten 	d->1	f->3	i->1	s->1	t->1	
lten!	 ->2	
lten,	 ->1	
lten.	D->3	T->1	
ltena	 ->1	
ltenb	e->4	
ltene	r->18	
ltens	 ->3	
lter 	s->1	t->1	
ltera	d->3	n->1	r->4	
ltern	a->12	
ltesi	s->3	
ltet 	d->1	f->1	o->1	v->1	ä->1	
ltet"	,->1	
ltet.	 ->1	J->1	S->1	
ltfle	r->1	
ltför	 ->39	
lthen	 ->3	,->1	s->2	
lthet	 ->2	
ltibe	t->1	
ltid 	a->9	b->7	d->1	f->6	g->2	h->12	i->2	k->5	l->1	m->2	n->4	o->1	p->1	r->2	s->4	t->4	u->1	v->3	y->1	ä->6	
ltid,	 ->2	
ltid.	O->1	
ltida	 ->1	
ltide	r->1	
ltids	s->1	
ltiet	n->3	
ltig 	i->2	o->1	
ltiga	 ->7	
ltigh	e->12	
ltigt	 ->4	
ltiho	p->1	
ltila	t->1	
ltill	v->17	
ltima	t->1	
ltina	t->5	
lting	 ->2	,->1	.->2	
ltisk	a->1	
ltjäm	t->3	
ltmer	 ->1	
ltnin	g->48	
ltog 	1->1	i->1	
lton.	H->1	
ltraf	i->1	
ltral	i->1	
ltrap	e->1	
ltrer	a->1	
ltro 	t->1	
lträd	a->1	e->6	
lts -	 ->1	
lts a	v->1	
lts f	ö->1	
lts i	 ->2	
lts m	e->1	
lts o	c->1	m->1	
lts p	å->1	
lts s	å->1	
lts t	i->1	
lts u	t->1	
lts ä	n->1	
lts.K	o->1	
lts: 	v->1	
ltsam	m->1	
ltsed	a->3	
ltsit	u->1	
ltså 	E->1	a->5	b->2	d->2	e->4	f->5	g->1	i->11	k->1	l->1	m->2	p->2	r->3	s->11	t->5	v->5	
ltså,	 ->2	
ltur 	2->20	b->2	d->1	f->2	h->1	i->4	o->2	p->1	s->4	u->1	v->1	ä->2	
ltur,	 ->11	
ltur-	 ->1	
ltur.	O->1	T->1	V->1	
ltur?	M->1	
ltura	k->1	n->1	r->6	
lture	l->28	n->30	r->6	
lturf	o->1	
lturh	i->1	
lturo	m->1	
lturp	o->5	r->3	
lturs	e->5	
lturu	t->1	
ltäck	a->4	
lucka	 ->1	"->1	,->1	
lucko	r->2	
luddi	g->2	
luder	a->4	
luftb	u->1	
lufto	m->1	
luför	a->1	
lugn 	o->1	
lugna	 ->2	d->1	n->1	s->1	
lukar	 ->2	
lukas	.->1	
lukt 	p->1	
lukta	r->1	
lump 	a->2	s->1	
lump.	D->1	
lumra	 ->1	
lunch	t->1	
lunda	 ->12	.->1	r->1	
lundr	i->1	
lunta	r->4	
lunto	r->1	
lupsk	h->1	
lural	i->1	
luras	 ->1	
lurat	 ->1	
lures	 ->1	
lus a	n->1	
lus t	r->1	
lusiv	 ->1	a->1	e->17	t->1	
lussa	 ->1	s->1	
lust 	s->1	
lust.	V->1	
lustb	r->1	
luste	n->2	r->5	
lut -	 ->1	
lut 8	8->2	
lut 9	4->1	
lut a	n->1	t->4	v->2	
lut b	e->3	o->1	ö->2	
lut d	i->1	
lut e	n->2	
lut f	a->1	o->1	r->5	ö->3	
lut g	o->1	
lut h	a->4	
lut i	 ->7	n->9	
lut k	a->2	o->1	
lut l	a->1	y->1	ä->1	å->1	
lut m	e->1	y->1	ö->1	
lut n	r->1	ö->10	
lut o	c->6	m->20	
lut p	l->1	å->10	
lut r	e->1	
lut s	e->1	k->1	o->12	t->1	ä->1	
lut t	a->1	i->1	
lut u	n->1	t->3	
lut v	a->1	i->2	
lut ä	n->1	r->3	
lut å	s->1	
lut, 	a->1	f->1	h->3	i->2	o->3	s->2	t->1	v->1	
lut. 	D->1	
lut.D	e->2	å->1	
lut.F	r->1	
lut.I	n->1	
lut.N	a->2	
lut.O	c->1	
lut.S	k->1	
lut.T	v->1	
lut.V	a->1	
lut; 	d->1	
luta 	a->2	d->4	e->2	f->2	g->2	i->1	k->1	m->6	o->12	p->1	r->1	s->6	u->1	v->1	Ö->2	
luta,	 ->5	
lutad	,->1	.->18	e->11	
lutaf	r->10	
lutan	 ->3	,->2	d->26	v->1	
lutap	o->1	
lutar	 ->8	.->1	
lutas	 ->8	p->2	
lutat	 ->11	s->3	
lutau	n->3	
lutbe	t->2	
lutbi	l->3	
luten	 ->9	,->2	.->3	s->1	
luter	 ->8	
lutet	 ->50	,->2	.->1	?->1	s->1	
lutfö	r->9	
lutgi	l->8	
lutha	n->1	
luthe	r->1	
lutio	n->101	
lutit	 ->3	s->1	
lutko	m->1	
lutli	g->72	
lutna	 ->8	,->3	.->4	
lutni	n->40	
lutpe	r->1	
lutre	s->3	
luts 	k->1	
lutsa	m->14	t->41	
lutsc	e->1	
lutsf	a->11	ö->1	
lutsk	o->14	
lutsp	r->4	
lutsr	ä->1	
lutst	a->1	
lutve	c->2	r->1	
lutän	d->5	
lux, 	n->1	
lv an	s->1	
lv ar	b->1	
lv at	t->3	
lv be	s->1	
lv bi	d->1	
lv da	g->1	
lv fr	å->2	
lv fö	r->3	
lv go	d->1	
lv ha	r->2	
lv hö	r->1	
lv i 	d->1	e->1	s->1	
lv ko	m->1	
lv me	d->2	
lv oc	h->1	k->2	
lv sa	m->1	
lv se	 ->1	
lv sk	a->1	
lv so	m->3	
lv sä	g->1	
lv ta	 ->1	
lv ti	m->2	
lv un	d->1	
lv ut	a->1	
lv va	r->1	
lv ve	r->1	
lv är	 ->3	
lv år	 ->1	
lv, h	e->2	y->1	
lv, m	e->2	
lv.De	t->1	
lv.Ja	g->1	
lv.Ko	m->1	
lv.Vi	 ->1	
lva E	u->1	
lva a	n->1	v->1	
lva b	e->2	j->1	o->1	ä->1	
lva d	a->1	e->2	
lva f	ö->1	
lva h	a->1	
lva i	 ->1	
lva k	a->2	u->1	ä->3	
lva l	a->1	
lva m	å->1	
lva o	c->3	m->1	
lva r	e->1	
lva s	k->1	o->1	t->2	y->1	
lva t	i->3	
lva u	n->1	
lva v	e->27	ä->1	
lva ä	r->2	
lva å	r->2	
lva, 	d->1	i->1	s->1	
lva.D	e->1	
lva.L	å->1	
lva.N	ä->1	
lva.O	m->1	
lva.V	å->1	
lval.	S->1	
lvand	e->1	
lvar 	e->1	i->1	o->1	s->2	ä->1	
lvar,	 ->1	
lvar.	I->1	N->1	S->1	V->1	
lvare	t->1	
lvarl	i->62	
lvbes	t->3	
lvbio	g->1	
lvbär	a->1	
lver 	o->1	u->1	
lver,	 ->1	
lvera	 ->2	d->6	r->1	
lverk	 ->13	,->1	.->1	a->76	e->8	n->12	s->2	
lvers	i->1	
lvet 	o->1	
lvfal	l->2	
lvför	t->1	
lvhjä	l->1	r->1	
lvida	 ->1	
lvill	i->1	
lvini	s->1	
lvis 	A->1	a->2	b->1	d->3	e->3	f->5	g->2	i->2	k->1	m->1	n->1	o->4	p->1	r->1	s->3	v->1	ä->3	å->2	ö->1	
lvis,	 ->2	
lvkla	r->20	
lvkos	t->1	
lvmil	j->1	
lvnin	g->3	
lvoff	e->1	
lvoly	m->1	
lvplå	g->1	
lvrak	 ->1	.->2	?->1	e->2	
lvsty	m->1	r->6	
lvstä	n->8	
lvsäk	e->1	
lvt d	i->1	
lvt h	a->2	
lvt k	o->1	
lvt s	o->1	
lvt å	r->2	
lvtid	s->1	
lvtim	m->2	
lvväg	s->2	
lväga	 ->1	.->1	g->6	
lvägg	i->3	
lvänd	a->1	
lvänn	e->1	
lvänt	 ->1	
lvärd	i->2	
lväxt	 ->7	,->2	.->2	b->1	e->8	
lvår 	k->1	
lvåre	t->2	
lvårs	s->2	
lvö, 	f->1	
lvö.D	e->1	
lvön 	s->1	
ly fö	r->1	
ly åt	e->1	
ly! G	e->1	
ly, k	a->1	v->1	
ly.An	d->1	
ly.Vi	 ->1	
lybet	ä->1	
lycka	 ->12	,->1	.->1	?->1	d->13	n->13	s->24	t->20	
lyckl	i->9	
lycko	r->16	s->1	
lycks	b->1	d->3	f->2	r->2	ö->1	
lyckö	n->5	
lyda 	u->2	
lydan	d->1	
lydel	s->2	
lyder	 ->3	
lyft 	f->2	
lyfta	 ->4	n->2	
lyfte	r->2	
lyfto	r->3	
lyg, 	h->1	
lyga 	m->1	
lygan	d->1	
lygbl	a->1	
lyger	 ->1	
lyget	 ->1	
lygkr	a->1	
lygni	n->1	
lygpl	a->4	
lygsa	m->4	
lygtr	a->2	
lykta	 ->1	
lykte	n->2	r->1	
lykti	n->13	
lym a	t->1	
lym o	m->1	
lymen	 ->1	
lymer	 ->1	
lympi	c->1	s->1	
lyr f	r->1	
lys -	 ->1	
lys a	v->16	
lys b	e->1	
lys f	a->1	ö->1	
lys g	e->1	
lys i	 ->1	
lys j	a->1	
lys o	c->2	
lys s	o->1	
lys v	i->1	
lys, 	a->1	d->1	u->1	v->1	
lys.D	e->2	
lys.F	r->1	
lys.G	e->1	
lys.H	ä->1	
lys?D	e->1	
lys?I	 ->1	
lysa 	o->2	u->3	
lysan	d->4	
lysat	o->2	
lysen	 ->5	
lyser	 ->2	.->1	a->15	
lysni	n->4	
lyssn	a->28	i->1	
lyst 	f->1	m->1	
lytan	d->12	
lytel	s->1	
lytt 	ö->1	
lytt.	J->1	
lytta	 ->6	r->3	s->1	t->1	
lyttn	i->4	
lyver	i->1	
lywoo	d->1	
lz en	 ->1	
lz sa	d->2	
lzen.	J->1	
lzman	n->2	
läcka	 ->2	d->1	
läcke	r->1	
läcko	r->1	
läckt	 ->2	e->1	
läder	 ->19	a->1	i->2	
lädja	 ->4	n->3	s->1	
lädje	 ->7	
läds 	d->1	m->1	r->1	å->2	ö->1	
lägar	n->1	
läge 	d->2	g->1	m->2	s->3	ä->1	
läge,	 ->1	
läge.	H->1	V->1	
lägen	 ->2	,->1	h->12	
läger	,->1	
läges	b->1	r->2	
läget	 ->16	,->1	.->2	
lägg 	f->1	g->1	h->2	i->4	k->1	l->1	s->1	t->4	u->4	v->1	
lägg,	 ->1	
lägg.	F->1	
lägga	 ->92	,->1	n->76	s->11	
lägge	n->2	r->39	t->2	
läggn	i->27	
läggs	 ->17	,->1	b->1	f->1	k->1	
lägli	g->1	
lägna	 ->6	,->2	
lägre	 ->8	.->2	n->1	
lägse	n->2	t->4	
lägsn	a->5	
lägst	a->1	
läkar	e->3	k->2	
läkem	e->1	
läkta	d->1	r->2	
läkte	t->1	
läkti	n->1	
lämna	 ->26	d->6	n->2	r->19	s->10	t->18	
lämni	n->5	
lämpa	 ->40	d->1	n->2	r->9	s->42	t->6	
lämpl	i->60	
lämpn	i->68	
lända	 ->1	r->2	t->1	
lände	r->184	t->1	
länds	k->26	
länga	s->1	
längd	 ->2	e->2	
länge	 ->35	
längn	i->3	
längr	e->62	
längs	 ->2	
längt	a->1	
länka	 ->2	
länni	n->1	
länt.	J->1	
läpad	e->1	
läpp 	a->1	k->1	
läpp,	 ->1	
läpp.	D->1	
läppa	 ->4	n->2	
läppe	n->3	r->1	t->1	
läpph	ä->1	
läpps	r->1	
läppt	e->3	
lär e	x->1	
lära 	f->1	k->1	o->1	s->3	å->1	
lärar	e->2	
lärde	 ->1	
lärdo	m->7	
lärli	n->1	
läroa	n->1	
läros	a->1	
lärt 	g->1	o->1	s->1	
läs t	e->1	
läs u	n->1	
läs y	t->1	
läsa 	k->1	o->1	v->1	
läsba	r->2	
läser	 ->6	
läsfr	ä->1	
läsku	n->1	
läsni	n->2	
läst 	D->1	d->1	e->2	
lästa	n->1	
läste	 ->1	
lät d	ä->1	
lät m	i->1	
lät s	i->1	k->1	o->1	
lätt 	a->3	f->1	k->1	l->1	s->1	t->2	
lätt.	A->1	K->1	
lätta	 ->20	d->2	r->17	
lättf	ö->1	
lätti	l->2	
lättn	a->1	
lättv	i->2	
läxan	?->1	
läxat	 ->1	
läxor	.->1	
lå Eu	r->1	
lå at	t->6	
lå ba	s->1	
lå el	l->1	
lå en	 ->3	
lå fa	s->6	
lå ih	o->1	
lå ko	m->3	n->1	
lå me	d->1	r->1	
lå nå	g->1	
lå pr	i->1	
lå rå	d->1	
lå sa	m->1	
lå si	g->1	
lå va	d->1	k->1	
lå ve	m->1	
lå vi	s->1	
låda 	f->1	
lådef	ö->1	
låder	 ->1	)->7	a->3	
låend	e->1	
låg a	r->1	
låg d	e->1	
låg h	ö->1	
låg i	n->1	
låg n	i->2	
låg t	i->1	
låga 	g->1	k->1	t->1	v->1	ö->1	
låger	i->1	
lågt 	s->1	v->1	
lånan	d->1	
lånbo	k->1	
lång 	a->2	e->1	i->1	l->1	o->3	p->1	r->2	s->10	t->11	v->2	
lång,	 ->1	
lång.	N->1	
långa	 ->10	
långd	r->1	
långf	r->1	ä->1	
långr	a->1	
långs	a->6	i->7	
långt	 ->34	.->3	g->11	i->4	
långv	a->6	
lånin	g->1	
lår B	a->1	
lår a	t->6	v->1	
lår d	e->1	ä->2	
lår e	n->2	r->1	t->3	
lår f	r->1	
lår i	 ->3	n->1	
lår j	a->4	
lår k	o->2	
lår m	a->1	e->1	
lår n	o->1	
lår r	e->1	
lår s	j->1	n->1	
lår t	i->1	
lår v	a->1	i->5	
lår ä	r->2	
lår".	J->1	
lår. 	E->1	
lår.M	a->1	
lår?S	o->1	
lås a	t->2	v->1	
lås b	l->2	
lås d	e->2	
lås e	n->1	
lås g	e->1	ö->1	
lås i	 ->11	
lås m	o->1	
lås p	å->1	
lås t	i->2	
lås.D	e->1	
låser	 ->3	
låss 	m->1	
låst 	s->1	
låsta	 ->2	
låt e	r->1	
låt m	i->15	
låt o	s->8	
låta 	E->1	J->1	a->2	b->3	d->10	e->2	f->2	h->1	j->1	k->1	l->1	m->4	n->1	o->2	p->2	r->2	s->4	t->1	
låtan	d->3	
låtas	 ->6	
låten	 ->4	h->2	
låter	 ->20	,->1	.->1	v->1	
låtet	 ->1	
låtit	 ->2	s->1	
låtli	g->5	
låtna	 ->5	.->1	
låts 	e->1	f->1	m->1	å->1	
låtsa	s->2	
lécha	r->1	
löden	a->1	
lödet	 ->2	
lödig	t->1	
löfte	 ->3	n->8	
löjad	e->1	
löjan	d->1	
löjar	 ->3	
löjas	.->1	
löjev	ä->3	
lökmo	d->1	
lömma	 ->13	:->1	
lömme	r->2	
lömsk	a->1	
lömt 	A->1	a->1	b->1	e->1	
lön f	ö->1	
lönar	 ->1	
lönas	,->1	
löne-	 ->1	
lönea	r->1	
löner	 ->1	
lönsa	m->5	
lönt 	a->1	
lönta	g->3	
löpa 	e->1	u->1	
löpan	d->6	
löper	 ->9	.->1	
löpt 	u->5	
löpte	 ->2	
lörda	g->1	
lös -	 ->1	
lös d	e->1	
lös e	n->1	
lös k	ä->1	
lös s	u->1	
lös.D	e->1	
lösa 	d->9	e->2	f->1	g->2	h->1	i->1	k->2	m->4	n->1	o->2	p->6	s->2	u->2	v->3	
lösa,	 ->3	
lösa.	F->1	I->1	M->1	
lösar	 ->1	
lösas	 ->5	.->1	
löser	 ->1	i->3	
löses	 ->1	
lösgö	r->1	
löshe	t->44	
lösni	n->52	
lösry	c->1	
löst 	d->2	f->1	i->2	o->2	p->1	r->1	v->1	
löst,	 ->1	
lösta	 ->3	,->1	.->2	
löste	s->1	
lösts	.->1	
löt a	t->1	
löt d	e->1	
löt v	i->1	
lötsl	i->4	
lövsk	o->1	
løn, 	i->1	m->1	
m "Eq	u->1	
m "Eu	r->1	
m "Ku	l->1	
m "Kv	i->1	
m "nå	g->1	
m "or	m->1	
m "va	l->1	
m "öp	p->1	
m - K	a->1	
m - a	t->4	
m - e	t->1	
m - i	n->1	
m - k	o->1	
m - m	e->2	
m - o	c->1	m->2	
m - p	r->1	
m - s	o->1	y->1	
m - t	r->1	
m - v	a->1	i->1	
m 1 0	0->1	
m 150	 ->1	
m 16 	0->1	
m 198	6->1	
m 199	7->1	9->1	
m 20 	m->1	p->1	å->1	
m 28 	p->1	
m 3-l	i->2	
m 314	 ->1	
m 35 	m->2	
m 350	 ->1	
m 40 	m->1	å->1	
m 400	 ->1	
m 45 	c->1	
m 50 	p->1	
m 5b-	o->1	
m 6,0	7->1	
m 80 	ä->1	
m Agu	s->1	
m Ahe	r->1	
m Ala	v->1	
m Alp	e->1	
m Amo	k->1	
m Ams	t->2	
m Apa	r->1	
m Atl	a->1	
m BSE	 ->1	
m Bar	a->1	
m Bel	g->1	
m Ber	e->1	g->3	t->1	
m Bla	k->1	
m Bow	i->1	
m Bri	t->1	
m Bry	s->1	
m CEN	:->1	
m Cey	h->1	
m Coc	i->1	
m Cox	 ->1	
m Da 	C->1	
m Dal	a->1	
m Dan	m->2	
m De 	g->1	
m Det	 ->1	
m Dim	i->1	
m Dut	r->1	
m EG-	d->3	
m EMU	:->1	
m EU 	I->1	d->1	f->1	h->2	k->3	o->1	s->2	
m EU,	 ->1	
m EU-	e->1	i->1	
m EU.	A->1	D->1	R->1	
m EU:	s->3	
m Ehu	d->1	
m Ell	e->1	
m Eri	k->1	
m Eti	o->1	
m Eur	o->73	
m FBI	 ->1	
m FPÖ	 ->1	
m Flo	r->1	
m Fra	n->2	
m För	b->1	e->3	
m GUS	P->1	
m Gal	e->1	
m Gen	e->2	
m Gol	a->1	
m Goo	d->1	
m Gre	k->2	
m Hai	d->3	
m Hat	z->2	
m Hed	k->1	
m Hit	l->1	
m INT	E->1	
m Ind	i->1	
m Irl	a->1	
m Isr	a->1	
m Ita	l->2	
m Jon	a->1	c->1	
m Jör	g->2	
m Kau	k->1	
m Kos	o->4	
m Kou	c->1	
m Lan	g->6	
m Lib	e->1	
m Llo	y->1	
m Mal	t->1	
m Mar	i->1	
m McC	a->1	
m McN	a->1	
m Ned	e->1	
m Off	i->1	
m PPE	-->1	
m Pak	i->1	
m Pal	a->1	
m Pay	s->1	
m Por	t->1	
m Pow	e->3	
m Pro	d->1	
m Rac	k->1	
m Ric	h->1	
m Rot	h->1	
m SEK	 ->1	
m Sch	e->2	r->1	
m Sei	x->2	
m Sjä	t->1	
m Sko	t->1	
m Spe	n->1	
m Syr	i->1	
m Tam	m->1	
m The	a->3	
m Tib	e->2	
m Tor	r->1	
m Tot	a->1	
m Tur	k->4	
m Vär	l->1	
m Wal	e->2	
m Wie	n->1	
m a p	r->1	
m abs	o->2	
m acc	e->1	
m adv	o->2	
m age	n->1	r->2	
m agr	o->1	
m ald	r->1	
m all	 ->3	a->29	i->1	m->3	t->16	v->5	
m alt	e->1	
m amb	u->1	
m ame	r->1	
m and	r->10	
m anf	ö->2	
m ang	e->3	
m ank	o->1	
m anl	ö->2	
m ann	a->2	
m ano	n->1	
m ans	e->3	j->1	l->3	t->3	v->14	ö->1	
m ant	a->6	i->3	o->4	
m anv	ä->8	
m app	l->1	
m arb	e->17	
m arg	u->1	
m arm	é->1	
m arr	e->1	
m art	i->2	
m asy	l->5	
m att	 ->398	
m av 	A->1	B->1	E->4	F->1	P->1	a->1	b->1	c->2	d->7	e->6	f->6	g->1	k->5	l->1	m->2	o->1	p->1	r->1	s->3	t->2	u->3	v->2	
m av,	 ->1	
m avf	a->2	
m avg	i->2	r->1	ö->4	
m avk	l->1	u->1	
m avl	i->1	o->1	
m avs	e->3	k->1	l->5	t->1	
m avt	a->1	
m avv	i->2	
m b) 	i->1	
m bak	d->1	g->1	
m bal	a->1	
m ban	d->1	
m bar	a->3	
m bea	k->2	
m bed	r->7	ö->1	
m bef	i->5	o->1	r->2	ä->1	
m beg	r->2	ä->2	å->3	
m beh	a->9	o->11	ö->10	
m bek	a->3	r->2	v->2	ä->3	
m bel	a->1	
m bem	y->1	
m beo	r->1	
m ber	 ->1	ä->2	ö->12	
m bes	e->1	i->1	k->7	l->6	t->10	v->1	ä->1	ö->1	
m bet	a->7	e->1	o->2	r->3	t->1	y->3	ä->3	
m bev	i->6	
m bid	r->7	
m bil	a->1	i->1	
m bin	d->1	
m bio	s->1	
m bit	e->1	
m bl.	a->2	
m bla	n->2	
m ble	v->2	
m bli	r->4	
m bly	.->1	
m bor	 ->4	d->7	g->1	
m bos	a->1	ä->1	
m bot	t->1	
m bri	s->1	t->2	
m bro	m->1	t->3	
m bru	k->1	
m bry	r->1	t->1	
m brå	d->3	
m bud	g->4	
m byg	g->1	
m byr	å->1	
m bär	 ->5	
m bät	t->2	
m båd	a->2	e->3	
m böc	k->1	
m bör	 ->12	j->2	
m böt	e->1	
m c) 	l->1	
m can	c->1	
m cen	t->1	
m cha	r->1	
m cho	c->1	
m cor	p->2	
m dag	 ->1	a->1	e->1	l->2	o->3	
m dam	m->1	
m de 	1->1	P->1	a->10	b->6	d->3	e->13	f->9	g->8	h->8	i->13	k->9	l->3	m->6	n->9	o->8	p->2	r->8	s->15	t->7	u->4	v->11	y->1	ä->5	å->1	
m de,	 ->1	
m deb	a->3	
m dec	e->1	
m def	i->3	
m del	a->2	e->1	n->1	t->3	
m dem	 ->2	o->4	
m den	 ->117	,->1	.->2	n->29	
m der	a->3	
m des	s->36	
m det	 ->214	,->3	.->8	?->1	a->3	t->67	
m dia	l->1	
m dif	f->1	
m dik	t->1	
m dio	x->1	
m dip	l->1	
m dir	e->7	
m dis	k->7	p->1	
m djä	v->1	
m dog	.->1	
m dom	i->1	s->4	
m dra	b->9	r->3	
m dri	c->1	f->1	v->1	
m dry	g->1	
m du 	ä->1	
m dub	b->1	
m dyk	e->1	
m där	 ->4	,->1	.->1	f->5	i->1	
m då 	a->1	f->2	h->1	o->1	v->1	
m dål	i->2	
m död	a->1	
m döe	n->1	
m döl	j->1	
m döm	t->1	
m eff	e->3	
m eft	e->10	
m ege	n->5	
m egn	a->1	
m ej 	l->1	
m eko	n->5	
m el-	S->4	
m ele	k->1	
m ell	e->5	
m eme	l->1	
m emo	t->17	
m en 	P->1	S->1	a->10	b->6	c->2	d->10	e->12	f->16	g->6	h->3	i->4	j->1	k->13	l->5	m->13	n->9	o->7	p->7	r->13	s->21	t->3	u->9	v->7	y->1	ä->1	ö->3	
m enb	a->1	
m end	a->6	
m ene	r->5	
m enh	e->1	
m enl	i->4	
m eno	r->1	
m ens	 ->1	a->1	k->1	
m er 	b->1	f->1	t->1	
m era	 ->4	
m erf	a->1	
m erk	ä->1	
m ers	ä->1	
m ert	 ->5	
m erö	v->1	
m etc	.->1	
m ett	 ->124	,->1	
m eur	o->10	
m ex 	a->1	
m exa	k->1	m->1	
m exc	e->2	
m exe	m->9	
m exp	o->1	
m fad	d->1	
m fak	t->3	
m fal	l->7	
m far	l->1	
m fas	c->1	t->10	
m fat	t->9	
m fem	 ->2	
m fic	k->1	
m fin	a->9	n->30	
m fis	k->4	
m fjo	r->1	
m fla	g->1	
m fle	r->6	
m fly	g->1	k->1	r->1	t->2	
m fod	e->1	
m fol	k->2	
m fon	d->1	
m for	d->4	s->2	t->12	
m fos	s->1	
m fra	m->27	n->2	
m fre	d->6	
m fri	 ->1	h->6	s->1	
m fru	 ->2	
m frä	m->1	
m frå	g->6	n->13	
m ful	l->1	
m fun	d->1	g->3	
m fus	k->1	
m fyl	l->1	
m fyr	a->1	
m fäl	l->1	
m fär	d->1	
m får	 ->6	
m fåt	t->3	
m föl	j->7	l->1	
m för	 ->109	.->1	b->12	d->7	e->55	f->5	h->5	k->1	l->11	m->2	n->7	o->8	r->2	s->40	t->8	u->7	v->7	
m gam	l->1	
m gar	a->5	
m gav	s->1	
m ge 	d->1	f->1	
m gem	e->19	
m gen	e->3	o->11	
m ger	 ->10	
m ges	 ->4	
m get	t->1	
m gic	k->1	
m gil	l->1	t->1	
m giv	i->1	
m gjo	r->10	
m glo	b->1	
m god	 ->1	k->7	
m gra	n->1	t->1	
m gri	p->2	
m gru	n->11	p->2	
m grä	n->2	
m gäl	l->22	
m gån	g->1	
m går	 ->9	
m gåt	t->2	
m göm	m->1	
m gör	 ->30	s->6	
m ha 	e->1	
m had	e->4	
m ham	n->3	
m han	 ->17	d->19	k->1	s->4	t->1	
m har	 ->147	m->5	
m has	t->1	
m hav	e->2	
m hed	r->1	
m hel	a->2	h->4	s->43	t->3	
m her	r->3	
m het	s->1	
m hin	d->2	
m hit	 ->1	t->11	
m hjä	l->3	r->3	
m hob	b->1	
m hon	 ->10	
m hot	a->1	e->2	
m hum	a->2	
m hur	 ->28	u->4	
m hys	e->1	
m häl	s->2	
m hän	d->10	g->6	t->1	v->1	
m här	 ->11	.->3	j->2	r->2	
m häv	d->4	
m hål	l->8	
m hår	t->1	
m hög	 ->1	a->1	r->1	s->1	
m hör	 ->3	
m i B	e->1	r->1	
m i C	e->1	
m i E	U->1	u->1	
m i G	u->1	
m i H	e->1	
m i N	e->1	
m i T	a->2	u->1	y->1	
m i U	r->1	
m i a	l->1	n->1	
m i b	e->1	å->1	ö->1	
m i d	a->19	e->15	
m i e	n->2	t->2	
m i f	a->2	i->1	l->2	o->1	r->10	ö->2	
m i g	r->1	
m i h	a->1	e->2	u->1	ä->1	ö->2	
m i k	a->1	
m i l	i->1	
m i m	a->1	o->13	å->1	
m i n	o->1	y->1	
m i o	c->2	r->1	
m i p	a->3	l->1	r->3	
m i r	e->3	å->1	
m i s	a->1	e->2	i->7	j->2	l->1	t->6	y->1	
m i t	i->2	r->1	
m i u	n->1	
m i v	a->1	e->2	i->3	å->1	
m i Ö	s->1	
m i å	r->1	
m i ö	v->1	
m ick	e->4	
m idé	n->1	
m ifa	l->1	
m ifr	å->1	
m ige	n->1	
m ihå	g->1	
m in 	p->1	
m inb	e->1	
m ind	i->3	u->3	
m inf	o->5	r->1	ö->12	
m ing	e->8	i->1	å->2	
m ini	t->2	
m ink	o->1	
m inl	e->9	
m inn	e->29	
m ino	m->8	
m inr	e->1	i->1	ä->5	
m ins	p->1	t->3	
m int	e->105	r->3	
m inv	a->2	o->1	
m isr	a->1	
m jag	 ->134	,->2	
m jor	d->6	
m ju 	M->1	m->1	ä->3	
m jus	t->9	
m jäm	f->1	l->1	
m jär	n->1	
m kam	m->1	
m kan	 ->53	d->1	i->1	s->3	
m kap	i->2	t->2	
m kar	a->1	t->4	
m kem	i->1	
m kla	r->1	s->1	
m koa	l->1	
m kod	e->1	
m kol	l->4	
m kom	 ->2	m->139	p->5	
m kon	c->2	f->1	k->21	s->4	t->3	v->1	
m kor	r->2	t->8	
m kos	t->6	
m kra	f->1	v->2	
m kri	n->1	t->5	
m krä	v->18	
m kul	t->7	
m kun	n->1	
m kur	s->1	
m kva	n->1	
m kvi	n->1	
m kän	n->5	s->1	
m kär	n->6	
m köp	e->1	
m kör	s->1	
m lad	e->4	
m lag	e->1	s->6	t->8	
m lan	d->2	
m led	a->13	d->8	e->8	n->1	
m leg	i->1	
m let	a->1	
m lev	e->6	
m lib	e->2	
m lig	g->16	
m lik	a->1	n->1	s->3	
m lit	e->1	t->1	
m liv	s->16	
m lju	s->1	
m lok	a->1	
m lyc	k->2	
m lyd	e->1	
m lyf	t->1	
m lyk	t->1	
m lys	s->1	
m läc	k->1	
m läg	e->1	g->7	
m läk	a->1	
m läm	n->7	p->4	
m län	d->2	g->3	
m lät	t->1	
m låg	 ->1	a->1	
m lån	g->2	
m löp	e->1	
m lös	n->4	
m mai	n->1	
m maj	o->2	
m mak	r->1	
m man	 ->96	,->1	n->1	
m mar	k->5	
m max	i->1	
m med	 ->33	b->8	d->2	e->2	f->1	g->3	l->17	v->2	
m mel	l->3	
m men	 ->3	a->2	
m mer	 ->6	v->1	
m mes	t->1	
m mil	i->1	j->8	
m min	 ->10	a->2	d->1	i->5	s->1	
m mis	s->4	
m mit	t->1	
m mod	e->3	
m mot	 ->2	i->2	o->1	p->1	s->7	
m mus	i->1	
m myc	k->9	
m myn	d->8	
m män	n->4	s->9	
m mär	k->1	
m måh	ä->1	
m mål	 ->2	
m mån	a->1	g->4	
m mås	t->32	
m möj	l->52	
m nar	k->1	
m nat	i->3	u->6	
m naz	i->3	
m ned	e->1	g->1	
m neg	a->1	
m nek	a->1	
m ni 	a->1	b->1	f->5	g->1	h->5	i->5	k->7	n->3	o->1	p->1	r->2	s->9	t->4	v->18	ä->1	
m ni,	 ->5	
m ni.	D->1	
m nio	 ->1	
m nor	m->2	
m nu 	a->1	f->4	g->1	h->5	i->2	l->1	m->1	p->1	r->2	t->1	u->1	v->1	ä->4	
m num	e->1	
m ny 	l->1	
m nya	 ->2	
m nyl	i->2	
m nys	s->1	
m nyt	t->1	
m näm	n->5	
m när	 ->10	i->1	
m näs	t->1	
m någ	o->16	r->14	
m nöd	v->1	
m nöt	k->1	
m oac	c->1	
m obe	g->1	h->1	
m och	 ->72	
m ock	s->19	u->1	
m off	e->1	r->2	
m oft	a->4	
m oge	n->1	
m oli	k->3	
m olj	e->2	
m oly	c->1	
m om 	6->1	E->1	H->1	S->1	a->2	b->1	d->9	e->1	f->1	g->1	i->2	j->1	k->3	l->1	m->3	n->1	r->3	s->1	t->1	u->2	v->4	
m omb	e->1	
m ome	d->1	
m omf	a->4	ö->1	
m oml	o->1	
m omr	å->8	ö->2	
m oms	ä->1	
m omö	j->1	
m onö	d->1	
m ord	e->2	f->8	v->1	
m ori	e->1	
m oro	a->1	n->1	
m ors	a->3	
m oss	 ->1	,->2	.->1	
m oti	l->1	
m par	l->24	t->1	
m pek	a->2	
m pen	n->1	s->1	
m per	s->3	
m pla	c->1	n->3	
m pol	i->6	
m pos	i->1	
m poä	n->1	
m pra	k->2	
m pre	s->3	
m pri	n->3	o->3	s->1	
m pro	b->3	d->2	g->3	j->3	
m pub	l->1	
m pum	p->1	
m pun	k->2	
m på 	-->1	7->1	a->5	b->1	d->12	e->6	f->2	g->4	h->1	k->1	l->1	m->1	n->4	o->1	r->1	s->4	t->4	v->2	
m på.	D->1	
m påg	å->1	
m påm	i->1	
m påp	e->1	
m påt	a->1	v->1	
m påv	e->8	
m rad	i->1	
m ram	 ->1	e->51	
m rap	p->1	
m ras	i->2	
m rat	i->1	
m red	a->34	u->1	
m ref	o->9	
m reg	e->15	i->5	l->5	
m rek	o->1	
m rel	a->6	e->1	i->1	
m rep	u->1	
m res	a->1	e->1	o->6	p->5	t->1	u->2	
m ret	o->1	
m rev	i->2	
m rik	t->5	
m rim	l->2	
m ris	k->8	
m rol	l->1	
m rul	l->2	
m rus	t->1	
m ryg	g->1	
m rys	s->1	
m räc	k->1	
m räk	e->1	
m rät	t->14	
m råd	 ->1	d->1	e->32	g->1	s->1	
m rör	 ->13	
m rös	t->3	
m röv	a->1	
m s.k	.->1	
m sad	e->3	
m sag	t->4	
m sak	 ->2	e->2	n->3	
m sam	a->3	b->1	l->4	m->17	o->2	t->7	v->1	
m san	n->1	
m sat	t->2	
m sch	a->1	
m sed	a->5	
m seg	l->3	
m sek	t->2	
m sen	a->1	
m ser	 ->5	
m sex	 ->1	
m sin	 ->4	a->2	
m sit	t->6	u->2	
m sju	k->1	n->1	
m sjä	l->1	
m sjö	f->1	
m ska	d->4	l->63	p->8	t->4	
m ske	r->8	t->4	
m ski	l->2	s->1	
m skj	u->1	
m sko	g->3	l->1	n->1	
m skr	e->1	i->1	o->2	ä->3	
m sku	l->27	
m sky	d->5	
m skö	t->1	
m slo	g->1	
m slu	t->7	
m små	 ->3	
m sna	b->1	r->1	
m sne	d->1	
m soc	i->2	
m sol	i->1	
m som	 ->130	,->1	l->1	
m spe	c->6	l->1	n->2	
m spo	n->1	
m spr	i->2	å->1	
m sta	d->1	r->4	t->10	
m ste	l->1	
m sti	m->1	
m sto	r->2	
m str	a->5	i->1	u->5	
m sty	r->3	
m stä	l->10	n->1	r->3	
m stå	l->2	n->4	r->21	
m stö	d->13	r->1	t->1	
m sub	s->2	v->2	
m sva	r->3	
m syf	t->9	
m syn	d->2	
m sys	s->5	t->5	
m säg	e->1	s->1	
m säk	e->16	r->1	
m sär	s->3	
m sät	t->1	
m så 	a->2	b->1	f->1	i->2	k->1	m->5	o->2	s->2	v->1	ä->2	
m såd	a->8	
m sål	e->1	
m såt	i->1	
m sök	e->1	
m sör	j->2	
m t.e	x->2	
m t.o	.->1	
m tag	i->2	
m tal	a->5	r->1	
m tan	k->2	
m tar	 ->6	
m tas	 ->5	
m tax	-->1	
m tib	e->1	
m tid	 ->2	e->1	i->8	t->1	
m til	l->112	
m tio	t->1	
m tjä	n->3	
m tog	 ->2	s->3	
m tol	e->2	k->3	
m tra	g->1	n->16	
m tre	 ->5	t->1	
m tro	r->1	t->1	
m trä	d->5	
m tur	i->1	
m tve	k->1	
m två	 ->4	n->1	
m tyc	k->2	
m tyd	e->3	l->2	
m tyn	g->1	
m tys	k->1	
m tyv	ä->2	
m täc	k->2	
m tän	k->1	
m täp	p->1	
m und	e->20	
m uni	o->22	
m upp	 ->1	b->1	e->2	f->6	g->2	k->1	l->2	m->5	n->2	r->4	s->9	t->1	
m ur 	E->1	e->1	
m urs	p->1	ä->6	
m ut 	a->1	
m ut.	J->1	
m uta	n->5	r->2	
m utb	i->5	
m utd	e->1	
m ute	s->1	
m utf	o->1	ö->6	
m utg	i->1	å->3	ö->7	
m uti	f->1	
m utj	ä->1	
m utl	a->1	ä->1	
m utm	a->1	ä->1	
m utn	y->1	
m utr	i->2	
m uts	e->2	k->3	t->6	ä->1	
m utt	a->2	j->10	r->2	
m utv	e->8	i->4	ä->1	
m utö	v->1	
m vad	 ->16	
m vag	a->1	
m val	 ->1	d->1	t->1	u->1	
m van	 ->3	l->1	
m var	 ->23	a->1	f->2	i->5	j->7	k->2	
m ved	e->1	
m vel	a->1	
m vem	 ->2	
m ver	k->20	
m vet	e->5	
m vi 	a->28	b->14	d->9	e->6	f->13	g->11	h->38	i->37	j->4	k->22	l->6	m->9	n->7	o->2	r->3	s->23	t->14	u->7	v->16	ä->7	å->1	ö->3	
m vi,	 ->3	
m vi?	.->1	
m via	 ->1	
m vid	 ->10	t->3	
m vik	t->2	
m vil	j->1	k->17	l->21	
m vin	d->1	
m vis	a->9	e->1	s->12	t->2	
m vit	b->5	
m von	 ->3	
m vor	e->2	
m vrä	k->1	
m vux	i->1	
m väc	k->3	
m väg	e->1	r->3	
m väl	j->3	l->1	
m vän	t->2	
m vär	l->1	
m väs	e->1	
m vår	 ->9	a->4	t->6	
m yrk	e->1	
m ytt	e->3	r->1	
m Öst	e->4	
m äge	r->2	
m ägn	a->1	
m ägt	 ->1	
m än 	e->1	h->1	i->1	m->1	o->1	r->1	
m änd	r->12	å->5	
m änn	u->4	
m änt	l->3	
m är 	-->1	1->1	a->21	b->10	d->17	e->17	f->11	g->2	h->5	i->13	k->6	l->6	m->14	n->5	o->8	p->8	r->5	s->14	t->7	u->6	v->9	y->2	ä->3	
m är,	 ->1	
m äte	r->1	
m äve	n->15	
m åkl	a->1	
m åkt	e->1	
m åla	g->1	
m åli	g->1	
m år 	b->1	e->1	f->1	h->1	s->4	
m år,	 ->1	
m år.	D->2	
m åre	n->3	t->2	
m års	 ->1	r->1	
m åsa	t->1	
m åsi	k->1	
m åst	a->1	
m åsy	f->4	
m åte	r->17	
m åtg	ä->7	
m åtm	i->1	
m öar	n->1	
m öka	d->1	r->1	t->1	
m ökn	i->1	
m öms	e->1	
m öns	k->1	
m öpp	e->5	n->2	
m öro	n->1	
m öst	e->2	
m öve	r->23	
m övr	i->1	
m!Den	n->1	
m!Det	 ->1	
m!Men	 ->1	
m!Tro	r->1	
m".De	t->1	
m) om	 ->1	
m); a	n->1	
m, Ku	l->1	
m, al	d->1	l->1	
m, an	n->1	s->1	
m, at	t->4	
m, av	 ->1	
m, bl	a->1	
m, bå	d->1	
m, bö	r->2	
m, de	n->3	s->1	t->7	
m, dä	r->1	
m, då	 ->1	
m, ef	t->5	
m, en	 ->1	l->2	
m, et	t->1	
m, ex	e->1	
m, fi	n->1	
m, fr	a->1	u->1	ä->1	
m, fö	r->3	
m, ge	n->1	
m, gr	u->1	
m, ha	r->3	
m, he	r->2	
m, hu	r->1	
m, i 	S->1	d->1	h->1	l->1	v->1	
m, id	r->1	
m, in	k->1	
m, ja	g->1	
m, ju	 ->1	s->1	
m, ka	n->2	
m, kr	o->1	
m, kv	i->1	
m, le	d->1	
m, me	d->4	n->8	
m, na	z->1	
m, ni	 ->1	
m, nä	r->2	
m, nå	g->1	
m, oc	h->20	
m, om	 ->1	
m, op	p->1	
m, or	g->1	
m, pr	i->1	
m, på	 ->3	g->1	
m, re	g->1	
m, sa	m->1	
m, se	x->1	
m, so	m->7	
m, sp	o->1	
m, sä	r->2	
m, så	 ->4	d->1	
m, ti	l->1	
m, tr	å->1	
m, up	p->1	
m, ut	a->6	i->1	ö->1	
m, va	d->1	l->1	r->1	
m, ve	t->1	
m, vi	a->1	d->1	l->7	
m, än	d->1	
m, är	 ->3	
m, äv	e->5	
m, åt	m->1	
m- oc	h->1	
m-el-	S->1	
m. De	t->1	
m. Dä	r->1	
m. Då	 ->1	
m. Ho	n->1	
m. Hu	r->1	
m. Ma	n->1	
m. av	s->2	
m. de	 ->1	
m. i 	e->1	
m. än	n->1	
m. är	 ->1	
m.(Ap	p->1	
m., d	e->1	
m.. F	r->1	
m..(F	R->1	
m.All	a->1	
m.Att	 ->1	
m.Av 	e->1	
m.Avb	r->1	
m.Avs	e->1	
m.Bet	ä->1	
m.Bud	g->1	
m.De 	a->1	k->1	s->1	ä->2	
m.Den	 ->5	n->2	
m.Des	s->2	
m.Det	 ->20	t->4	
m.Där	 ->1	f->4	
m.EG-	d->1	
m.EKS	G->1	
m.En 	s->1	
m.Eur	o->1	
m.Exp	e->1	
m.Fru	 ->5	
m.För	 ->3	
m.Gen	o->2	
m.Gör	 ->1	
m.Her	r->10	
m.Hur	 ->1	u->1	
m.I d	e->2	
m.I n	o->1	
m.I r	e->1	
m.Inf	ö->1	
m.Ino	m->1	
m.Jag	 ->17	
m.Kom	m->1	
m.Kos	t->1	
m.Kul	t->1	
m.Låt	 ->1	
m.Man	 ->1	
m.Med	 ->3	
m.Men	 ->8	,->1	
m.Mån	g->1	
m.Nat	u->1	
m.Nej	,->1	
m.Ni 	t->1	
m.Nu 	v->1	
m.När	 ->3	
m.Någ	r->1	
m.OMR	Ö->1	
m.Och	 ->4	
m.Om 	d->1	n->1	
m.Pro	b->2	
m.Ref	o->1	
m.Res	t->1	
m.Råd	e->1	
m.Sam	t->1	
m.Slu	t->2	
m.Som	 ->2	
m.Sta	t->2	
m.Syf	t->1	
m.Så 	j->1	
m.Til	l->1	
m.Tro	t->1	
m.Tyv	ä->1	
m.Ur 	d->1	
m.Vad	 ->1	
m.Vem	s->1	
m.Vi 	a->1	b->1	h->5	k->4	m->2	t->1	u->1	v->1	
m.Vid	 ->2	
m.Vil	k->1	
m.m.O	c->1	
m.Änd	r->1	
m.Är 	d->1	
m/rik	e->1	
m: As	t->1	
m: Nä	r->1	
m: de	 ->1	n->1	
m: du	b->1	
m: en	 ->1	
m: pa	r->1	
m; de	t->2	
m?Det	t->1	
m?Jag	 ->1	
m?Men	a->1	
m?Vil	k->2	
mI. f	ö->1	
ma - 	j->1	p->1	
ma 16	7->1	
ma Br	y->1	
ma Eu	r->1	
ma Ha	i->2	
ma Ma	a->1	
ma al	l->2	
ma am	b->1	
ma an	d->1	s->1	
ma ar	b->1	t->1	v->1	
ma at	t->15	
ma av	 ->1	s->1	
ma be	f->1	g->1	l->1	s->1	t->1	
ma bi	l->2	
ma bo	r->4	
ma br	o->1	
ma bä	t->1	
ma da	g->1	
ma de	 ->7	b->5	f->1	m->1	n->3	s->1	t->4	
ma di	m->1	
ma dr	a->1	
ma en	 ->6	
ma er	 ->1	
ma et	t->3	
ma eu	r->2	
ma fa	l->1	
ma fi	s->1	
ma fr	a->6	e->1	å->4	
ma fö	l->1	r->16	
ma gr	u->1	
ma gä	l->2	
ma gå	r->1	
ma ha	d->1	n->1	r->1	
ma hi	t->2	
ma ho	s->1	
ma hu	r->1	
ma hä	f->1	n->1	r->1	
ma hå	l->1	
ma hö	g->1	
ma i 	E->1	F->1	a->1	d->5	e->1	h->1	k->1	s->1	
ma i.	N->1	S->1	
ma if	a->1	r->1	
ma ig	å->1	
ma ih	å->14	
ma in	 ->5	o->3	r->1	s->4	t->2	
ma iv	e->1	
ma jo	r->5	
ma ka	n->1	r->1	
ma kl	i->1	
ma ko	k->1	m->1	n->4	s->1	
ma kr	a->4	i->1	
ma ku	l->2	
ma kä	r->1	
ma la	n->2	
ma li	n->1	
ma lä	n->1	
ma lå	n->2	
ma lö	s->1	
ma ma	j->1	r->1	s->1	
ma me	d->17	
ma mi	n->1	
ma mo	n->1	t->1	
ma mä	n->1	
ma må	l->5	
ma mö	j->2	
ma na	m->1	
ma ni	v->1	
ma nä	m->2	r->2	
ma nå	g->3	
ma oc	h->4	
ma om	 ->5	s->2	
ma or	d->1	g->3	o->1	
ma os	s->1	
ma pa	r->1	
ma pe	r->2	
ma po	l->5	
ma pr	i->2	o->4	
ma pu	n->1	
ma på	 ->7	.->1	p->1	
ma re	a->1	g->2	s->6	
ma ri	k->4	s->1	
ma ro	l->1	
ma rä	t->2	
ma sa	k->13	
ma si	g->1	n->1	t->1	
ma sk	a->1	u->1	ä->2	
ma sl	u->1	
ma sn	a->1	
ma so	m->9	r->1	
ma st	a->1	i->1	r->4	ä->1	å->48	
ma su	m->1	
ma sv	å->2	
ma sy	n->1	s->1	
ma sä	g->1	t->17	
ma så	 ->1	
ma te	x->1	
ma ti	l->12	
ma ty	c->1	p->1	
ma un	i->1	
ma up	p->2	
ma ut	k->9	m->1	r->1	v->1	
ma va	l->5	r->1	
ma vi	d->1	l->4	
ma vä	r->1	
ma vå	g->1	r->1	
ma är	 ->3	
ma år	,->1	s->1	
ma ås	i->1	
ma åt	 ->1	g->1	
ma öv	e->9	
ma, a	t->1	
ma, d	e->1	v->1	å->1	
ma, f	r->1	ö->1	
ma, m	e->1	
ma, o	c->1	
ma, s	å->1	
ma, u	t->1	
ma.De	t->1	
ma.He	r->2	
ma.Ja	g->4	
ma.Om	 ->1	
ma.Or	s->1	
ma.Vi	d->1	
ma: a	n->1	
ma: u	n->1	
maceu	t->1	
mad o	c->1	
made 	f->1	h->1	i->1	k->1	u->4	v->1	
mades	 ->1	
maffä	r->1	
mage 	s->1	
mager	 ->1	
magh 	m->1	
magin	ä->1	
magna	.->1	
magni	t->1	
magog	e->1	i->3	
mail 	m->1	
mains	t->7	
maj 1	9->3	
maj 2	0->1	
maj f	ö->1	
maj, 	o->1	
maj.J	a->1	
maj.T	o->1	
major	i->41	
makol	o->1	
makro	e->5	f->1	
makt 	-->1	a->1	f->6	i->3	m->1	o->2	v->1	
makt,	 ->2	
makt.	B->1	D->2	J->2	
maktb	a->2	e->2	
maktd	e->1	i->1	
makte	n->6	r->2	
maktf	ö->1	
makth	a->1	å->1	
maktk	o->1	
maktl	ö->3	
maktm	e->2	i->1	
makäm	n->1	
mal b	i->2	
mal e	f->1	l->1	
mal f	ö->1	
mal p	l->1	
mal s	ä->1	
mala 	e->2	g->1	l->1	m->1	r->1	
malay	a->1	
malis	e->3	t->1	
malit	e->1	
malt 	7->1	i->2	s->2	
malt.	D->1	O->1	V->1	
malte	s->3	
man "	e->1	
man E	U->1	
man F	o->1	
man I	m->2	
man R	o->1	
man a	 ->1	b->1	l->7	n->12	t->12	v->2	
man b	a->3	e->11	l->3	o->4	r->1	ä->1	ö->8	
man d	e->10	i->1	o->1	r->1	ä->8	å->3	ö->1	
man e	f->1	m->1	n->7	r->4	
man f	a->4	i->1	o->3	r->3	u->2	ä->1	ö->16	
man g	a->1	e->4	i->1	o->1	r->3	å->2	ö->8	
man h	a->27	i->2	o->2	u->1	ä->5	å->1	ö->2	
man i	 ->30	f->1	n->57	
man j	a->1	u->2	ä->2	
man k	a->21	n->1	o->9	r->4	u->4	ä->1	
man l	a->1	i->1	y->2	ä->10	å->1	ö->1	
man m	e->13	i->1	o->1	y->1	å->19	ö->1	
man n	a->4	o->1	u->9	ä->1	
man o	c->17	m->5	v->1	
man p	a->1	l->2	o->1	r->2	å->8	
man r	a->1	e->9	i->3	ö->1	
man s	a->6	e->11	i->6	j->1	k->44	l->3	n->1	o->1	t->4	v->1	ä->8	å->1	
man t	a->12	i->13	r->2	v->1	y->1	ä->3	
man u	n->7	p->6	r->1	t->3	
man v	a->5	e->9	i->19	r->1	ä->4	
man y	t->1	
man ä	g->2	n->3	r->8	v->2	
man å	 ->2	r->1	s->1	t->2	
man ö	v->7	
man! 	A->5	B->2	D->33	E->5	F->12	G->2	H->1	I->10	J->74	K->5	L->6	M->5	N->5	O->2	P->4	R->4	S->9	T->8	U->4	V->17	Ä->7	Å->3	Ö->1	
man!A	m->1	
man!D	e->2	
man!E	f->1	n->1	
man!J	a->6	
man!M	i->1	
man!S	a->1	
man!T	a->1	i->1	
man!U	n->1	
man!V	i->2	
man, 	a->9	b->2	d->8	e->4	f->21	h->39	i->3	j->3	k->31	m->16	n->4	p->4	r->1	s->7	t->2	u->2	v->4	ä->11	
man.D	e->1	
man.H	u->1	
man.K	o->1	
man.M	e->1	
man.S	l->1	
man: 	n->1	
mana 	E->1	T->1	d->4	e->1	f->1	k->1	m->1	p->2	s->1	
manad	e->2	
manar	 ->31	,->1	
manas	 ->4	
manat	 ->3	
manbi	n->1	
manbl	a->2	
manbo	e->1	
manbr	o->1	
manbu	n->1	
manda	t->23	
mande	 ->70	,->2	.->4	t->4	
mandi	e->1	
mandr	a->1	
manen	t->8	
maner	.->1	
manfa	l->2	t->12	
manfö	r->1	
mang 	a->1	f->2	h->2	i->1	m->1	n->1	o->1	s->1	u->1	
mang,	 ->1	
mang.	E->1	H->1	J->1	O->1	
mange	n->1	r->2	t->1	
manha	n->47	
manhä	n->1	
manhå	l->53	
manif	e->1	
manin	g->28	
manis	m->1	t->2	
manit	e->1	ä->1	
manjä	m->1	
manka	l->9	
manko	m->2	p->1	
manla	g->1	
manli	g->1	
manlä	n->1	
mann 	o->1	ä->1	
mann,	 ->1	
mann-	g->1	
manna	l->1	r->1	
manne	n->24	
manni	n->2	
mano 	P->2	
mans 	a->3	b->1	f->2	g->1	i->2	m->19	s->1	t->1	v->1	ä->1	
mans,	 ->3	
mans.	L->1	
mans;	 ->1	
mansa	t->3	
mansk	o->9	
mansl	a->5	u->2	
mansm	ä->1	
manst	r->1	ä->5	
mansv	a->1	
mansä	t->5	
mantr	a->3	ä->35	
manöv	r->1	
mapla	n->1	
mar B	r->2	
mar P	o->1	
mar R	o->1	
mar a	t->1	v->1	
mar e	f->1	l->1	
mar f	o->1	r->1	ö->3	
mar i	 ->6	n->1	
mar k	a->1	o->1	
mar n	a->1	u->1	ä->1	
mar o	c->4	m->2	s->3	
mar p	e->1	å->1	
mar s	e->1	i->2	o->2	
mar t	i->1	
mar u	t->1	
mar ö	v->2	
mar! 	F->1	
mar, 	a->3	f->1	i->1	m->1	n->1	o->4	s->1	u->1	v->1	
mar.B	a->1	
mar.H	e->1	
mar.J	a->2	
marbe	t->88	
mare 	2->1	a->3	b->9	f->3	i->1	k->1	m->3	o->3	p->4	s->3	t->3	v->2	ä->2	
mare,	 ->4	
mare.	D->1	H->1	N->1	V->1	Ä->1	
maren	 ->25	,->4	.->5	;->1	s->2	
margi	n->6	
marit	i->3	
mark 	-->1	b->1	e->2	h->1	i->2	k->2	l->1	m->1	o->4	p->1	s->4	t->2	v->1	
mark,	 ->3	
mark.	D->2	F->1	J->1	
marka	n->3	
marke	n->1	r->7	t->1	
markn	a->187	
marko	l->1	
marks	 ->2	
marle	d->1	
marna	 ->20	,->2	.->3	s->1	
mars 	1->1	2->1	i->1	m->1	o->1	
mars,	 ->3	
mars.	N->1	V->1	
marsc	h->1	
mas a	v->2	
mas b	l->1	
mas f	ö->1	
mas o	c->1	
mas p	å->3	
mas r	e->1	
mas s	j->1	å->1	
mas u	n->1	
mas ö	v->1	
mas, 	h->1	
maske	r->2	
maski	n->6	
masku	s->1	
masoc	h->1	
massa	 ->1	k->1	r->2	v->1	
massi	v->3	
massm	e->3	
mast 	a->1	
mast,	 ->1	
maste	 ->11	r->1	
masto	d->1	
mat a	l->1	r->1	
mat e	x->1	
mat f	r->1	ö->1	
mat s	o->1	ä->1	
mat u	r->6	
mat v	i->1	
mat.D	ä->1	
match	a->1	e->1	
matem	a->1	
mater	 ->1	i->27	
matet	 ->4	,->2	.->1	
matfö	r->4	
mati,	 ->1	
matik	,->1	e->4	
matio	n->72	
matis	e->1	k->37	
mativ	t->2	
matny	t->1	
matpe	n->1	
matpr	o->1	
mats 	a->2	
matta	 ->1	.->1	n->1	
mattn	i->1	
matum	 ->1	
mavta	l->3	
maxbe	l->1	
maxim	a->5	e->2	
mb ha	d->1	
mb.An	s->1	
mbads	 ->1	
mbala	m->1	
mband	 ->45	e->2	
mbar 	m->1	
mbara	 ->1	
mbard	e->1	
mbarg	o->1	
mbass	a->1	
mbatt	a->1	e->1	
mbeds	 ->1	
mben 	i->1	
mbeni	 ->2	.->1	
mber 	1->14	a->1	d->1	e->1	f->2	h->1	i->2	l->3	m->2	o->2	r->1	s->1	
mber,	 ->9	
mber.	 ->1	D->1	E->1	J->1	N->1	S->1	
mberv	e->1	
mbesö	r->2	
mbete	 ->4	.->1	
mbets	m->2	r->1	
mbett	s->2	
mbexp	l->1	
mbina	t->1	
mbiti	o->14	ö->12	
mblem	 ->1	
mblic	k->5	
mbnin	g->1	
mbol 	f->2	
mboli	s->7	
mbord	 ->1	
mbrot	t->2	
mbryo	s->1	
mbud 	e->1	r->1	
mbuds	m->10	
mbula	n->1	
mburg	 ->3	,->3	.->1	a->1	
mbus 	ä->1	
mbygd	.->1	
mbärl	i->4	
md at	t->1	
md hö	n->1	
md in	t->1	
md om	 ->1	
md ti	d->1	l->1	
md vi	l->1	
md, e	n->1	
md, h	a->1	
mda a	g->1	
mda m	o->1	
mda o	c->1	
mda r	e->1	
mda v	i->1	
mda å	t->3	
mda, 	e->1	
mde T	r->1	
mde i	 ->1	
mde m	a->1	e->1	
mde s	i->1	
mde.D	e->1	
mdefi	n->1	
mden 	ä->1	
mdes 	s->1	
mdhet	.->1	
mdiri	g->1	
mdriv	a->5	s->1	
mdöme	.->1	s->1	
me eg	e->1	
me få	r->1	
me fö	r->5	
me ko	m->1	
me oc	h->2	
me om	 ->1	
me so	m->4	
me åt	 ->2	
me, d	e->1	
me-fa	l->1	
me.Ko	m->1	
med "	a->2	e->1	
med -	 ->1	
med 1	2->1	3->2	4->1	6->1	9->1	
med 2	 ->2	0->2	4->1	7->2	8->1	
med 3	0->1	6->1	
med 5	 ->1	
med 8	0->1	
med A	.->1	m->2	
med B	S->1	a->1	
med D	a->2	
med E	-->1	D->1	U->1	r->4	u->12	
med F	r->4	
med G	A->1	
med H	a->4	
med I	n->1	s->2	
med J	ö->1	
med K	o->2	
med L	e->1	i->2	
med M	a->3	i->1	
med O	L->1	s->1	
med P	a->1	
med R	y->1	
med S	a->1	y->4	
med T	h->1	u->2	
med U	S->4	
med V	a->1	e->1	
med a	d->1	l->34	n->26	r->12	t->106	u->2	v->14	
med b	a->2	e->7	i->5	r->7	u->1	å->1	
med d	a->3	e->233	i->8	r->2	u->2	y->2	
med e	f->2	k->1	l->1	n->85	r->13	t->28	u->2	x->4	
med f	a->4	e->1	i->1	l->3	o->3	r->30	u->9	å->1	ö->37	
med g	a->1	e->6	i->1	l->2	o->5	r->4	
med h	a->3	e->3	j->24	o->1	u->5	ä->13	å->1	ö->2	
med i	 ->15	f->1	m->1	n->23	
med j	o->1	u->1	ä->1	
med k	a->5	i->1	l->1	n->1	o->31	r->7	u->1	v->9	ä->1	ö->1	
med l	a->2	e->2	i->8	ö->2	
med m	a->6	e->13	i->28	o->5	y->5	å->7	ö->4	
med n	a->13	e->3	u->3	y->4	ä->1	å->7	ö->7	
med o	c->10	f->1	j->1	l->2	m->20	r->6	s->8	
med p	a->13	e->5	l->1	o->3	r->8	s->1	u->2	å->17	
med r	a->1	e->19	i->2	ä->10	å->5	ö->1	
med s	.->1	a->9	e->1	i->26	j->1	k->7	l->2	m->1	n->1	o->6	p->5	t->36	u->2	v->2	y->2	ä->9	å->11	
med t	.->1	a->37	e->2	i->19	o->1	r->6	u->2	v->5	y->1	ä->1	
med u	n->6	p->6	r->1	t->17	
med v	a->13	e->6	i->16	ä->1	å->16	
med y	r->1	t->4	
med Ö	V->1	s->1	
med ä	n->4	r->5	
med å	r->2	t->4	
med ö	k->1	m->1	p->1	s->1	v->11	
med, 	a->1	d->2	e->1	g->1	m->2	n->1	o->3	p->1	s->1	v->1	
med.D	e->3	
med.F	ö->1	
med.V	i->2	
medan	 ->20	s->3	
medar	b->2	
medbe	s->15	
medbo	r->168	
medbr	o->1	
medde	l->59	
medel	 ->54	,->12	.->9	?->1	b->18	l->4	p->2	s->116	t->1	
medfi	n->2	
medfö	r->20	
medge	 ->3	r->9	s->5	t->1	
medgi	v->2	
medgö	r->2	
medhj	ä->1	
media	 ->5	l->1	s->1	t->1	
medic	i->1	
medie	r->5	
medin	f->1	
medkä	n->5	
medla	 ->2	r->1	
medle	m->334	n->12	t->1	
medli	d->2	n->2	
medve	r->19	t->42	
megap	r->1	
meka.	D->1	
mekan	i->10	
mell 	d->1	
mella	 ->4	n->207	
melle	r->67	
melli	 ->1	
mellt	 ->10	,->1	
mels 	i->1	
melse	 ->27	.->4	n->4	r->109	v->1	
men (	F->1	
men -	 ->3	
men A	m->1	
men C	a->1	
men E	u->1	
men F	ö->1	
men I	M->1	
men K	a->2	
men L	e->1	
men a	l->3	n->1	r->1	t->12	v->6	
men b	a->2	e->3	i->1	l->1	o->1	r->1	u->1	å->1	
men d	e->91	i->1	ä->4	å->1	
men e	f->3	g->1	n->8	t->1	
men f	a->1	e->1	o->1	r->4	ö->68	
men g	e->2	
men h	a->5	ä->1	
men i	 ->21	n->18	
men j	a->39	u->1	
men k	a->2	o->4	
men l	å->1	
men m	a->4	e->11	i->1	o->1	y->2	å->2	ö->3	
men n	a->2	i->3	u->4	ä->2	
men o	c->40	l->1	m->5	r->1	t->1	u->1	
men p	o->1	å->3	
men r	a->2	ä->1	å->1	ö->1	
men s	a->5	k->5	o->18	t->1	ä->1	å->3	
men t	a->1	e->1	i->5	r->2	v->1	y->3	
men u	n->4	
men v	a->2	e->1	i->41	ä->2	
men ä	n->2	r->4	v->9	
men ö	k->2	
men, 	W->1	a->1	d->2	e->2	f->4	h->1	i->2	m->2	o->2	s->6	v->1	ä->2	
men.D	e->5	
men.F	ö->1	
men.H	e->1	
men.J	a->5	
men.L	e->1	
men.M	e->1	
men.O	c->1	
men.U	p->1	
men.V	å->1	
men; 	f->1	ä->1	
men?V	i->1	
menad	e->2	
menan	d->2	
menar	 ->25	,->1	.->1	
menas	 ->2	
menda	t->33	
mende	r->12	
mener	g->3	
menet	 ->2	
menin	g->53	
menis	t->2	
mens 	a->2	e->1	f->2	k->1	o->1	r->1	u->1	ä->1	
mensa	m->196	
mensb	e->2	
mensi	o->13	
mensk	a->194	
ment 	-->2	1->1	a->4	b->2	e->1	f->34	g->2	h->8	i->15	k->4	l->1	m->7	o->18	p->1	s->33	t->7	u->2	v->3	ä->5	ö->3	
ment,	 ->21	
ment.	 ->1	D->2	E->1	F->2	H->1	I->4	J->4	L->1	M->1	N->1	P->1	
menta	 ->1	l->1	r->50	t->4	
mente	n->24	r->55	t->478	
mentf	r->6	
mentk	a->1	
mento	r->1	
mentp	o->2	
mentr	e->1	
ments	 ->2	b->1	f->1	k->6	l->28	u->2	
mentt	i->1	
mentv	a->1	ä->1	
mentä	r->2	
mer -	 ->4	
mer 2	 ->1	7->1	
mer 6	0->1	
mer B	S->1	r->1	
mer E	k->1	u->3	
mer G	r->1	
mer I	s->3	
mer J	ö->2	
mer N	a->1	
mer S	y->1	
mer T	u->1	
mer a	b->1	l->10	m->1	n->4	r->2	t->400	v->15	
mer b	e->4	o->3	y->1	ä->1	
mer d	e->50	i->1	j->3	o->2	r->1	y->1	ä->1	å->2	
mer e	f->5	k->1	l->5	m->2	n->6	t->3	x->1	
mer f	a->1	i->1	l->1	r->22	y->1	å->1	ö->24	
mer g	e->5	i->1	l->1	ä->1	
mer h	a->1	e->4	i->1	u->1	ä->3	ö->1	
mer i	 ->20	f->2	l->1	n->25	
mer j	a->11	u->4	
mer k	a->1	o->22	r->3	ä->2	
mer l	e->1	i->2	ä->2	å->4	ö->1	
mer m	a->7	e->17	i->2	y->2	ä->1	å->1	
mer n	a->2	i->9	ä->1	å->3	
mer o	a->1	c->65	f->1	m->16	s->1	
mer p	a->2	e->2	o->3	r->3	å->13	
mer r	a->4	e->2	å->1	
mer s	a->1	e->1	i->2	j->5	k->3	n->1	o->11	p->2	t->6	y->5	ä->4	å->5	
mer t	i->8	o->1	r->2	v->5	y->1	
mer u	n->3	p->1	t->7	
mer v	a->1	e->4	i->39	ä->3	å->2	
mer ä	n->35	r->1	v->6	
mer å	r->1	t->1	
mer ö	p->3	v->3	
mer!"	D->1	O->1	
mer, 	d->2	e->2	h->3	i->1	m->2	s->3	t->1	u->1	
mer. 	D->1	T->1	
mer.B	e->1	
mer.D	e->7	å->1	
mer.F	ö->1	
mer.H	e->1	
mer.I	 ->2	
mer.J	a->1	
mer.K	o->1	
mer.M	e->1	
mer.O	m->1	
mer.S	o->1	
mer.T	i->1	
mer.V	a->2	i->3	å->1	
mera 	E->4	I->1	a->2	b->1	c->1	d->3	e->3	f->2	i->2	k->1	m->1	o->5	p->4	s->4	t->1	u->1	v->2	ä->1	
merad	e->7	
meran	d->1	
merar	 ->4	
meras	 ->5	
meray	,->1	
merfo	r->22	
merge	r->1	
merik	a->17	
merin	g->18	
merit	e->1	
merna	 ->17	,->4	.->1	
merpa	r->1	
mers 	e->1	
mersa	m->1	
mersi	e->7	
mervä	r->5	
mes, 	j->1	
mesgi	l->1	
mest 	a->6	b->3	d->4	e->1	f->3	g->2	k->2	l->4	m->1	o->1	p->1	r->2	s->3	t->2	u->2	v->1	ä->1	
mesta	 ->1	,->2	d->2	
meste	r->4	
met "	K->2	
met (	i->1	
met -	 ->4	
met A	l->2	
met K	u->2	
met L	e->1	
met S	a->1	
met a	t->1	v->3	
met b	e->1	l->1	o->1	ö->2	
met e	l->1	n->1	r->2	
met f	i->1	r->1	ö->27	
met g	e->3	ä->1	
met h	a->1	i->1	o->1	ö->1	
met i	 ->6	n->4	
met k	o->2	
met l	i->1	ö->1	
met m	e->22	å->2	ö->1	
met n	ä->1	
met o	c->4	m->1	
met p	å->4	
met s	a->1	k->5	o->5	t->2	å->1	
met t	i->3	
met u	t->1	
met v	a->2	e->1	
met ä	r->19	
met) 	(->1	C->1	
met).	H->1	
met, 	E->1	d->3	f->1	i->1	k->1	s->4	u->1	v->2	ä->1	
met. 	a->1	
met.1	9->1	
met.B	e->1	
met.D	e->4	
met.E	t->1	
met.H	u->1	ä->1	
met.I	 ->3	
met.J	a->6	
met.M	e->4	
met.N	i->1	
met.O	c->1	
met.P	r->1	
met.V	i->2	
met: 	J->1	
met?K	ä->1	
metal	l->11	
meter	 ->4	n->1	
metod	 ->13	e->16	
metra	r->1	
mets 	e->1	o->1	r->1	
meuro	p->4	
mexis	t->2	
mfart	.->1	
mfatt	a->75	n->8	
mfina	n->1	
mflyt	t->1	
mform	u->3	
mfors	k->1	
mfund	e->5	
mfäll	d->1	
mfång	e->1	s->1	
mför 	E->1	a->73	b->1	d->5	e->4	f->1	h->1	l->1	m->3	o->10	r->1	s->2	t->1	v->2	ä->1	ö->1	
mföra	 ->71	,->1	l->1	n->46	s->24	
mförb	a->11	
mförd	a->1	e->14	r->27	
mföre	l->2	
mförh	a->2	
mförk	l->1	
mförs	 ->9	,->1	.->4	l->2	t->7	
mfört	 ->14	s->16	
mger 	a->1	
mgick	 ->2	
mgiva	n->1	
mgivn	i->1	
mgrip	a->4	
mgäng	e->1	
mgå e	n->1	
mgå i	 ->1	
mgå.F	ö->1	
mgåen	d->1	
mgång	 ->11	"->1	,->3	.->3	a->7	e->4	s->14	
mgår 	a->3	d->6	e->1	n->1	o->2	r->1	s->1	
mgår.	V->1	
mgått	 ->3	
mhet 	a->2	b->1	d->3	e->1	f->6	g->1	h->1	i->4	m->2	o->5	p->9	r->1	s->7	t->1	u->2	v->3	ä->4	å->5	
mhet,	 ->6	
mhet.	D->1	F->1	H->1	J->1	M->1	P->1	V->1	
mhet?	V->1	
mhete	n->18	r->3	
mhets	a->1	b->2	g->2	o->1	t->1	
mhuld	a->1	
mhäll	e->42	s->7	
mhärd	a->1	
mhäva	 ->2	s->1	
mhäve	r->1	
mhåll	a->10	e->3	i->3	s->1	
mhöge	r->14	
mhöll	 ->1	s->1	
mi - 	C->1	
mi at	t->1	
mi me	d->5	
mi oc	h->12	
mi är	 ->1	
mi, l	a->1	
mi, m	e->1	
mi, v	i->1	
mi.De	n->1	t->1	
mi.Fö	r->1	
mi? O	c->1	
mibes	t->2	
midda	g->13	
midig	 ->2	a->1	
midis	k->1	
mier 	o->1	
mier,	 ->1	
mier.	A->1	
miern	a->5	
mifin	a->1	
mig a	l->3	n->1	r->1	t->29	v->5	
mig b	a->6	e->2	ö->1	
mig d	e->4	o->1	ä->3	
mig e	m->1	n->2	r->1	t->2	
mig f	i->1	r->1	u->1	ö->10	
mig g	e->1	r->1	ä->1	ö->1	
mig h	a->3	e->2	
mig i	 ->10	n->5	
mig k	l->1	n->1	o->1	
mig l	i->1	ä->1	
mig m	e->3	o->1	y->5	ä->1	
mig n	e->1	u->1	ä->2	å->1	
mig o	b->2	c->12	m->11	
mig p	e->2	å->9	
mig r	i->1	
mig s	a->2	k->1	l->1	o->3	ä->5	
mig t	a->2	i->6	
mig u	n->4	t->1	
mig v	a->6	e->1	i->4	ä->1	
mig y	t->1	
mig ä	n->2	r->5	v->1	
mig å	 ->1	t->5	
mig ö	v->2	
mig!"	.->1	
mig, 	a->1	e->2	h->4	m->2	n->2	o->1	p->1	s->1	v->1	
mig.D	e->1	
mig.E	r->1	
mig.J	a->3	
mig: 	h->1	
mig?V	a->1	
miga,	 ->1	
mighe	t->2	
migra	n->2	t->8	
migre	r->1	
migt 	m->1	
miinn	e->1	
mik e	l->1	
mik o	c->1	
mikal	i->5	
mikap	i->1	
mikon	t->1	
mikra	v->2	
mikro	f->1	k->2	s->1	
milda	s->1	
mildr	a->3	
milia	-->1	
milis	 ->1	
milit	a->2	ä->6	
milj 	L->1	
milja	r->15	
milje	-->1	f->1	j->3	r->8	å->1	
miljo	n->63	
miljö	 ->8	!->1	,->11	-->2	.->6	a->4	b->4	d->2	e->4	f->10	i->1	k->26	l->1	m->14	n->39	o->5	p->14	r->3	s->24	u->1	v->9	
mille	n->7	
milst	o->1	
milän	g->1	
milön	e->1	
min -	 ->1	
min a	n->1	v->1	
min b	a->1	e->2	i->1	r->1	
min d	e->3	j->2	r->1	
min e	g->3	r->2	
min f	r->9	ö->5	
min g	l->2	r->21	
min i	 ->1	n->2	
min k	a->2	o->24	ä->1	
min m	a->1	e->18	
min o	c->12	r->1	
min p	e->1	l->2	o->1	r->1	
min r	e->3	ö->5	
min s	o->4	t->2	y->1	
min t	i->1	r->1	u->3	
min u	p->13	t->2	
min v	a->1	ä->1	
min å	s->9	
min ö	n->2	
min, 	e->1	m->1	u->1	
min.C	e->1	
min.D	e->1	
min.L	å->1	
min.M	e->1	
min.V	i->1	
mina 	a->1	b->1	d->27	e->1	f->2	g->5	i->2	k->20	o->1	r->1	s->2	t->4	u->1	ä->2	ö->2	
minal	i->3	p->1	
minan	s->1	
minar	i->1	
minat	i->2	
minde	 ->1	
mindr	e->52	
minel	l->3	
miner	a->16	i->28	
ming 	b->1	i->1	p->1	t->1	
ming"	,->1	
ming)	 ->2	.->1	
minim	a->1	e->1	i->19	o->1	u->5	
minir	e->1	
minis	t->95	
miniv	å->1	
minna	 ->21	s->2	
minne	 ->4	,->3	.->1	n->1	r->8	s->2	t->2	
minns	 ->6	
minor	i->22	m->2	
mins 	a->1	k->1	t->1	
minsk	a->47	n->16	
minst	 ->25	,->1	a->5	o->27	
minus	 ->3	g->2	
minut	 ->3	.->3	e->10	
minär	a->3	
mipar	a->1	
mirak	e->1	
miref	o->2	
mireg	l->3	
mis-f	ö->1	
mis-n	o->1	
mis.F	ö->1	
misk 	a->1	b->2	e->1	f->3	g->2	h->2	j->1	k->7	m->1	o->12	p->7	r->1	s->3	t->2	u->3	v->1	
misk.	D->1	
miska	 ->143	.->1	:->1	
miskt	 ->26	.->2	
mism 	h->1	p->1	ä->1	
misme	n->2	
miss 	b->1	i->1	m->1	o->1	p->1	s->1	v->1	
miss,	 ->5	
miss.	D->1	E->1	
missa	 ->1	r->1	t->1	
missb	r->10	
misse	n->1	
missf	a->1	o->2	ö->4	
missg	y->7	
missh	u->1	
missi	o->1151	
missk	ö->6	
missl	y->18	ö->1	
missn	ö->3	
missr	e->2	
misst	a->15	e->1	o->1	r->3	ä->4	
missu	p->2	
miste	 ->1	r->3	
misti	s->11	
mistl	i->1	
misty	r->4	
misär	 ->1	e->1	
mit d	e->1	
mit e	f->2	
mit f	r->7	
mit h	a->1	
mit i	 ->2	
mit m	e->3	y->2	
mit n	i->1	å->1	
mit t	i->6	
mit u	n->1	p->2	t->1	
mit v	i->1	
mit ö	v->6	
mit, 	b->1	f->1	m->1	
mit.M	o->1	
mit.P	a->1	
mita 	i->1	
mitet	 ->3	,->1	.->2	e->1	
mitis	k->1	m->2	
mitiv	a->1	
mitni	n->1	
mitra	k->5	
mits 	a->1	p->1	
mitt 	a->5	b->1	d->2	e->7	f->8	g->1	h->4	i->3	k->1	l->11	p->3	r->1	s->7	t->8	u->2	y->1	ä->3	
mitta	t->1	
mitte	n->2	
mitté	 ->10	e->4	f->2	n->41	s->2	
mium 	o->2	
mium,	 ->1	
mix.D	e->1	
mixen	 ->1	
miärm	i->10	
miåld	e->1	
mja a	n->2	
mja d	e->4	
mja e	n->7	t->1	
mja f	ö->3	
mja g	e->1	r->1	
mja h	å->1	
mja i	n->1	
mja k	u->1	v->2	ö->1	
mja l	i->2	
mja p	a->1	
mja s	a->1	t->1	y->2	
mja v	a->1	
mja y	r->1	
mja å	t->2	
mja.K	o->1	
mjand	e->17	
mjar 	e->2	k->1	p->1	r->1	t->1	
mjas,	 ->1	
mjat 	h->1	
mjuka	 ->1	
mjukn	i->2	
mka i	h->1	
mkar 	m->1	s->1	
mkast	a->1	
mkat 	s->1	
mkat,	 ->1	
mkomm	e->5	i->5	
mkrin	g->15	
mla U	C->1	
mla b	e->2	i->5	
mla d	e->1	
mla f	a->1	o->3	ö->2	
mla h	a->1	
mla i	n->5	
mla k	o->4	v->1	
mla l	ö->1	
mla m	a->2	
mla o	c->1	
mla r	e->1	
mla s	k->2	p->1	y->1	ä->1	
mla t	i->1	
mla u	p->1	
mlade	 ->2	
mlagd	a->3	
mlagt	 ->5	s->4	
mland	 ->1	,->1	.->1	
mlar 	p->1	u->1	
mlarf	o->1	
mlas 	e->1	
mlast	n->1	
mlat 	d->1	f->1	s->1	
mlats	 ->2	
mlen,	 ->1	
mlevn	a->1	
mlig 	d->1	h->1	i->1	k->2	
mlig.	V->1	
mliga	 ->18	
mlige	n->48	
mligg	a->1	
mligh	e->17	å->2	
mligt	 ->19	,->1	.->1	
mlik 	p->1	
mlikh	e->12	
mling	 ->9	,->4	.->2	a->2	e->5	s->37	
mloka	l->2	
mlägg	a->4	e->2	s->2	
mländ	e->1	
mläsn	i->2	
mläst	a->1	
mläxo	r->1	
mlösa	 ->1	,->1	
mlösh	e->3	
mm av	 ->1	
mma -	 ->1	
mma 1	6->1	
mma E	u->1	
mma a	m->1	n->2	r->3	t->15	v->1	
mma b	e->4	i->1	o->4	r->1	
mma d	a->1	e->16	r->1	
mma e	n->3	r->1	t->3	u->2	
mma f	a->1	i->1	r->9	ö->12	
mma g	r->1	ä->2	
mma h	a->1	i->2	o->1	ä->3	å->1	
mma i	 ->10	.->2	f->2	g->1	h->14	n->15	v->1	
mma j	o->5	
mma k	a->2	o->4	r->5	u->2	ä->1	
mma l	a->2	i->1	ä->1	å->2	ö->1	
mma m	a->1	e->17	i->1	o->1	ä->1	å->5	ö->2	
mma n	a->1	i->1	ä->4	å->3	
mma o	c->3	m->5	r->3	
mma p	a->1	e->2	o->5	r->5	u->1	å->7	
mma r	e->9	i->4	o->1	ä->2	
mma s	a->13	k->3	l->1	n->1	o->9	t->54	y->2	ä->17	å->1	
mma t	e->1	i->12	y->1	
mma u	n->1	p->1	t->11	
mma v	a->5	i->4	ä->1	å->1	
mma ä	r->3	
mma å	r->1	s->1	t->2	
mma ö	v->8	
mma, 	a->1	d->3	f->1	o->1	u->1	
mma.H	e->1	
mma.J	a->3	
mma.O	m->1	
mma: 	a->1	u->1	
mmad 	o->1	
mmade	 ->3	s->1	
mmal 	b->2	e->1	p->1	
mman 	d->3	f->1	i->2	m->10	n->1	o->1	t->1	ä->1	
mman,	 ->1	
mman.	M->1	
mmanb	i->1	l->2	o->1	r->1	u->1	
mmand	e->68	r->1	
mmanf	a->14	ö->1	
mmanh	a->47	ä->1	å->53	
mmanj	ä->1	
mmank	a->9	o->3	
mmanl	a->1	ä->1	
mmans	 ->31	,->3	.->1	;->1	a->3	l->7	m->1	t->5	ä->5	
mmant	r->35	
mmapl	a->1	
mmar 	e->2	f->1	i->3	k->2	n->2	o->4	p->1	s->1	t->1	u->1	
mmar!	 ->1	
mmar,	 ->8	
mmar.	J->1	
mmare	 ->21	,->3	.->3	n->37	
mmarl	e->1	
mmarn	a->3	
mmas 	a->1	o->1	p->1	r->1	u->1	ö->1	
mmas,	 ->1	
mmat 	a->1	e->1	f->1	v->1	
mmate	r->1	
mmats	 ->1	
mme e	g->1	
mme f	å->1	ö->5	
mme k	o->1	
mme o	c->2	m->1	
mme s	o->4	
mme å	t->2	
mme, 	d->1	
mmels	e->143	
mmen 	(->1	K->2	L->1	b->3	e->1	f->7	h->3	k->1	m->5	u->1	
mmen,	 ->6	
mmen.	D->4	H->1	J->2	L->1	M->1	V->1	
mmen;	 ->1	
mmend	a->33	e->12	
mment	a->24	e->13	
mmer 	-->4	2->2	6->1	B->1	E->4	G->1	I->3	S->1	T->1	a->410	b->5	d->47	e->11	f->25	g->5	h->8	i->39	j->15	k->12	l->1	m->21	n->14	o->26	p->7	r->3	s->22	t->11	u->8	v->42	ä->7	å->2	ö->2	
mmer,	 ->6	
mmer.	 ->1	D->1	I->1	J->1	V->2	
mmerf	o->22	
mmers	 ->1	a->1	i->7	
mmet 	"->2	(->1	-->1	A->2	K->2	L->1	S->1	b->1	e->4	f->12	g->2	h->2	i->1	k->2	m->1	o->5	s->10	u->1	v->1	ä->4	
mmet)	 ->2	
mmet,	 ->6	
mmet.	 ->1	1->1	D->2	I->1	J->4	M->2	O->1	
mmet:	 ->1	
mmets	 ->2	
mmiga	,->1	
mmigh	e->2	
mmigr	a->7	
mmigt	 ->1	
mmipa	r->1	
mmiss	i->1150	
mmit 	d->1	e->2	f->7	h->1	i->2	m->5	n->2	t->6	u->4	v->1	ö->6	
mmit,	 ->3	
mmit.	M->1	P->1	
mmits	 ->2	
mmitt	é->59	
mmon 	l->1	
mmor 	a->1	b->1	o->1	p->3	s->1	u->1	
mmor,	 ->1	
mmor.	V->1	
mmun.	D->1	
mmuna	l->3	
mmune	r->10	
mmuni	c->2	k->16	s->1	t->1	
mmöbl	e->1	
mn Ko	s->1	
mn by	t->1	
mn i 	E->1	
mn ka	n->1	
mn me	d->1	
mn må	s->2	
mn oc	h->1	
mn på	 ->1	
mn so	m->1	
mn sp	e->1	
mn sv	e->1	
mn, f	ö->1	
mn, m	e->1	
mn, u	t->1	
mn.De	 ->1	n->1	
mn.Me	n->1	
mn.Vi	t->1	
mna A	l->1	
mna L	i->1	
mna a	t->4	
mna b	i->1	
mna d	e->8	i->1	
mna e	t->4	u->2	x->1	
mna f	ö->5	
mna g	a->1	
mna h	a->2	o->1	u->1	ä->1	
mna i	 ->3	n->5	
mna k	o->1	
mna m	i->1	å->1	
mna n	å->1	
mna o	b->1	c->1	
mna p	r->1	å->1	
mna r	å->3	
mna s	i->1	k->2	n->1	o->1	t->1	y->1	
mna t	a->1	i->1	o->1	r->1	v->1	
mna u	t->3	
mna v	i->2	
mna, 	n->1	o->1	
mna.T	r->1	
mnad 	e->1	
mnade	 ->9	
mnand	e->4	
mnar 	a->1	d->14	e->1	f->1	h->1	i->7	j->6	k->2	m->3	o->6	r->2	s->5	u->3	v->8	å->1	
mnar.	M->1	O->1	U->1	
mnare	 ->1	.->2	n->1	
mnarn	a->6	
mnas 	a->2	d->1	f->1	i->3	o->1	p->1	t->3	
mnas,	 ->2	
mnat 	3->1	b->3	e->1	i->4	m->1	o->1	s->1	v->1	
mnats	 ->3	,->1	.->1	
mnavg	i->2	
mnbes	t->1	
mnda 	a->2	h->1	i->2	o->1	u->1	
mndas	 ->1	
mnde 	a->2	d->3	j->1	k->2	o->2	t->1	
mnde,	 ->4	
mnde.	D->1	K->1	
mndes	 ->1	
mne h	a->1	
mne i	 ->1	
mne s	o->1	
mne.D	e->2	
mne: 	N->1	
mnen 	a->1	h->1	i->1	n->1	o->3	s->3	v->2	
mnen,	 ->2	
mnen.	D->3	E->1	N->1	V->1	
mnena	 ->1	
mner 	-->1	d->1	j->1	n->1	
mner.	J->1	
mnet 	"->1	f->1	p->1	u->1	
mnet.	D->1	M->1	
mning	 ->30	,->6	.->6	:->1	a->11	e->25	s->5	
mnins	p->1	
mnkon	t->2	
mns a	l->1	
mns e	n->1	
mns f	ö->1	
mns h	ä->1	
mns i	 ->1	
mns m	ö->1	
mns o	c->1	
mns u	t->1	
mns.D	e->1	
mnt b	ö->1	
mnt e	x->1	
mnt f	ö->1	
mnt g	ä->1	
mnt i	 ->1	
mnt k	a->1	
mnt l	i->1	
mnt n	å->1	
mnt p	u->1	
mnt, 	a->1	i->1	
mnt.D	e->2	
mnts 	o->1	ä->1	
mnts,	 ->2	
mnts.	D->1	J->1	
mnupp	r->4	
mnvik	t->1	
mnvär	d->1	
mo, H	e->1	
mo, d	e->1	
mobil	i->7	
moco,	 ->1	
mod a	t->1	
mod e	n->1	
mod f	ö->1	
mod i	 ->1	
mod m	e->1	
mod s	o->1	
mod ä	r->1	
model	l->12	
moder	a->1	n->37	s->2	
modet	 ->6	
modif	i->3	
modig	a->3	t->1	
modli	g->12	
mofob	i->1	
mogen	 ->1	a->1	t->1	
moget	 ->1	
mogra	f->3	
moko 	C->5	
mokra	t->137	
moln 	o->1	
momen	t->5	
mområ	d->3	
momsp	l->1	
mon l	a->1	
monbe	h->1	
monet	a->1	ä->6	
moni 	o->1	
monis	e->13	k->4	
monit	o->1	
monnä	e->1	
monok	u->3	
monop	o->17	
monst	e->1	r->6	
monte	r->12	
mor a	v->1	
mor b	l->1	
mor o	c->1	
mor p	å->3	
mor s	o->1	
mor u	p->1	
mor, 	s->1	
mor.V	i->1	
moral	 ->1	e->1	i->5	
mord 	i->1	o->1	s->1	
mord,	 ->1	
mord.	U->1	
mordb	r->1	
morde	n->8	
mordi	s->1	
mordn	a->18	i->20	
morga	n->2	
morgo	n->37	
morse	 ->3	,->1	.->2	
morum	,->1	
mos O	z->1	
mosex	u->1	
mosor	,->1	
mot -	 ->1	e->1	
mot 1	3->1	
mot 5	 ->1	
mot A	i->1	
mot D	a->1	
mot E	U->2	u->7	
mot F	r->1	ö->2	
mot G	r->1	
mot H	a->3	
mot I	s->1	
mot J	o->3	
mot L	a->1	
mot M	o->1	
mot R	a->2	
mot S	o->1	
mot T	i->1	o->1	
mot U	N->1	
mot W	u->1	
mot a	i->1	l->7	n->4	r->2	t->12	v->9	
mot b	a->14	e->5	r->1	å->1	
mot d	e->56	i->2	o->2	
mot e	k->1	n->13	r->3	t->7	x->2	
mot f	o->1	r->7	ö->6	
mot g	e->1	l->1	
mot h	a->4	e->1	u->2	ä->2	
mot i	 ->3	d->1	n->6	
mot k	a->1	l->1	o->5	ö->1	
mot l	e->1	o->1	
mot m	a->4	e->5	i->1	ä->1	
mot n	a->3	ä->3	å->1	
mot o	e->1	l->3	s->3	
mot p	e->1	o->1	r->4	u->1	
mot r	a->2	e->3	å->4	
mot s	a->1	e->1	i->3	j->1	k->4	l->2	o->5	p->1	t->4	u->2	v->1	ä->1	
mot t	a->2	e->1	v->1	
mot u	n->2	p->1	
mot v	a->4	e->2	i->5	ä->1	å->4	
mot y	t->1	
mot Ö	s->3	
mot ä	n->1	r->1	
mot å	t->1	
mot ö	k->2	v->4	
mot! 	D->2	J->2	N->1	S->1	V->1	
mot, 	Z->1	a->5	d->1	h->2	o->1	s->2	t->1	u->1	ä->3	
mot. 	7->1	
mot.F	r->2	
mot.V	i->1	
motar	b->1	
moten	 ->22	.->2	s->2	
motgå	n->1	
motio	n->1	
motiv	 ->2	a->1	e->18	
motor	 ->1	.->2	c->4	i->2	
motpa	r->4	
motsa	t->23	
motst	r->1	y->3	å->12	
motsv	a->17	
motsä	g->8	t->9	
motta	g->16	r->1	
motve	r->4	
motvi	k->1	l->1	
motåt	g->3	
mouti	e->1	
mp Jö	r->1	
mp at	t->2	
mp fö	r->2	
mp i 	b->1	f->1	k->1	
mp me	l->1	
mp mo	t->4	
mp sj	ö->1	
mp.De	 ->1	
mpa -	 ->1	
mpa a	l->1	n->1	r->5	
mpa b	e->3	
mpa d	a->1	e->9	i->2	
mpa e	l->1	n->1	x->2	
mpa f	r->2	ö->10	
mpa g	e->2	l->1	
mpa i	 ->1	
mpa k	o->2	r->3	
mpa m	o->1	
mpa n	a->1	
mpa o	c->1	l->1	
mpa p	e->1	l->1	o->1	r->2	
mpa r	e->2	
mpa s	i->1	k->2	t->2	u->1	
mpa t	e->1	
mpa u	n->1	r->1	
mpa å	t->1	
mpad 	b->1	k->1	
mpagn	e->1	
mpake	t->1	
mpand	e->4	
mpanj	 ->3	.->1	e->2	
mpar 	d->3	e->1	f->3	m->2	o->2	ö->1	
mpar.	A->1	
mpas 	a->7	b->1	d->1	e->1	f->4	g->2	i->4	k->3	o->1	p->5	r->1	s->3	v->1	
mpas,	 ->1	
mpas.	-->1	D->4	K->1	P->1	V->1	
mpas:	 ->1	
mpass	i->1	
mpat 	f->1	m->1	t->1	
mpati	 ->4	e->1	s->3	
mpats	 ->4	.->1	
mpel 	-->2	B->1	N->1	R->1	a->2	b->2	d->1	e->1	f->10	g->2	h->6	i->5	n->2	o->4	p->20	r->1	s->7	t->1	v->1	ä->2	
mpel,	 ->5	
mpel.	J->1	M->1	V->1	
mpel:	 ->3	
mpelv	i->28	
mpen 	f->2	m->11	o->1	
mpen,	 ->1	
mpen.	H->1	
mpens	a->3	e->7	
mpera	 ->1	t->5	
mperi	o->3	
mpete	n->11	
mpic 	B->1	
mpisk	a->1	
mplan	e->8	t->1	
mplar	i->2	
mplem	e->11	
mplen	 ->3	
mplet	 ->3	t->14	
mplex	 ->1	.->1	a->1	t->1	
mplic	e->12	
mplig	 ->7	,->1	.->1	a->19	h->3	t->29	
mplim	a->3	e->1	
mplin	g->1	
mpnin	g->85	
mpone	n->4	r->3	
mpopu	l->1	
mpor,	 ->1	
mport	.->1	e->4	f->1	
mporä	r->2	
mproc	e->10	
mprog	r->15	
mproj	e->1	
mprom	i->22	
mpröv	a->6	n->2	
mpson	 ->1	
mptom	 ->1	
mpuls	 ->2	e->4	
mpunk	t->1	
mpåle	n->1	
mra e	u->1	
mra i	 ->1	
mra k	o->1	
mrad 	m->1	s->1	ö->5	
mrade	 ->3	.->1	
mrand	e->1	
mrapp	o->2	
mrar 	o->2	v->1	
mras 	n->1	
mras.	 ->1	
mrat 	S->1	o->1	
mre b	å->1	
mre f	r->1	ö->1	
mre h	a->1	
mre l	ä->1	
mre s	t->1	
mrest	e->1	
mring	a->1	
mrum 	f->1	
mrum,	 ->1	
mrund	a->1	
mrätt	 ->1	
mråd 	i->1	o->1	s->1	
mråd,	 ->1	
mråd.	L->1	
mråda	 ->2	
mråde	 ->57	,->14	.->23	:->1	;->1	?->1	n->130	t->90	
mråds	r->1	
mröst	n->57	
ms Bl	o->1	
ms an	s->2	
ms ef	t->2	
ms fö	r->1	
ms i 	d->1	
ms sä	k->1	
ms tu	r->1	
ms ut	i->1	
ms va	r->1	
ms- o	c->3	
ms-, 	u->1	
msa d	e->2	
msa u	t->1	
msan 	t->1	
msan.	V->1	
msar 	e->1	
msavt	a->2	
msbet	a->2	
msbro	t->1	
msesi	d->5	
msfrå	g->3	
msful	l->1	
msgrä	n->1	
mshav	e->1	
mshem	 ->1	
mside	s->1	
msign	a->2	
msk k	l->1	
mska 	r->2	s->1	
mskan	 ->1	
mskap	 ->1	e->1	
mskas	t->1	
mskin	l->1	
mskju	t->1	
mskri	d->1	
mskyd	d->4	
mslag	 ->2	s->1	
mslan	d->9	
mslut	 ->3	
mslän	d->27	
msnit	t->11	
msoll	m->1	
msorg	 ->8	s->1	
mspar	l->1	
mspli	k->1	
mspän	n->1	
msreg	e->1	
msrät	t->1	
msråd	 ->1	,->1	
mssta	r->1	t->283	
mst I	n->1	
mst a	n->1	r->1	
mst d	e->2	
mst e	n->1	t->1	
mst f	ö->1	
mst g	e->1	ö->1	
mst i	 ->1	n->5	
mst k	o->2	u->1	
mst l	o->3	
mst m	e->1	
mst o	c->1	m->2	v->1	
mst p	e->3	o->1	r->1	
mst s	k->1	
mst t	a->2	
mst u	t->3	
mst v	a->1	i->6	
mst ö	n->1	
mst.F	ö->1	
msta 	b->1	h->2	m->2	o->2	p->2	r->1	s->3	
mstad	t->1	
msteg	 ->22	,->2	.->2	e->6	
msten	 ->2	
mster	 ->2	,->2	.->1	d->39	n->1	
mstfö	r->1	
msthä	l->1	
mstkä	l->1	
mstol	 ->6	.->2	a->25	e->44	s->9	
mstra	r->1	
mstri	d->2	n->2	
mstru	k->10	
mstäl	l->35	
mstäm	m->4	p->1	
mstän	d->34	
mstå 	s->1	
mståe	n->5	
mstår	 ->1	
mstöt	a->1	
msvep	 ->1	
msvät	s->1	
msyn 	-->1	o->1	
msyn,	 ->1	
msyra	 ->3	
msätt	a->6	e->1	n->1	
msåtg	ä->1	
mt Au	s->1	
mt Ga	r->1	
mt He	b->1	
mt Wa	f->1	
mt al	i->1	
mt an	g->1	t->1	
mt ar	b->1	
mt as	y->1	
mt at	t->14	
mt av	 ->3	
mt ba	s->1	
mt be	s->2	v->1	
mt bi	l->1	
mt bo	r->1	
mt bö	r->1	
mt de	t->3	
mt ek	o->3	
mt en	 ->2	
mt er	a->1	
mt et	t->3	
mt eu	r->2	
mt fa	l->1	
mt fo	r->1	
mt fr	ä->1	å->2	
mt fö	l->2	r->7	
mt ha	n->1	
mt hå	r->3	
mt i 	a->1	e->1	f->1	
mt in	b->1	f->1	
mt jä	r->1	
mt ko	a->1	m->2	
mt ku	l->1	
mt kv	a->1	
mt lu	f->1	
mt lä	g->2	
mt me	d->1	
mt mi	n->1	
mt mo	t->1	
mt my	c->1	
mt må	s->2	
mt ne	d->1	
mt oc	h->5	
mt om	 ->7	r->3	
mt pa	r->2	
mt po	l->1	
mt på	 ->1	
mt ra	d->1	
mt re	g->1	k->1	s->1	
mt ry	k->1	
mt rä	t->2	
mt sa	m->1	
mt si	g->2	n->2	
mt sk	a->1	
mt st	r->3	y->1	ö->2	
mt sy	s->1	
mt ta	c->6	
mt ti	l->4	
mt un	d->2	
mt up	p->2	
mt ut	f->1	i->1	s->1	t->1	ö->1	
mt va	k->1	r->1	
mt vi	k->1	
mt vä	l->1	
mt yt	t->1	
mt än	d->1	
mt äv	e->2	
mt åt	 ->1	
mt ök	a->1	
mt öv	e->2	
mt, f	u->1	ö->1	
mt, g	r->1	
mt, v	a->1	
mt, ä	r->1	v->1	
mt.De	t->1	
mt.På	 ->1	
mt.Un	d->1	
mt.År	e->1	
mta s	i->1	y->1	
mta u	p->1	
mtaga	n->3	
mtagi	t->1	
mtagn	i->1	
mtal 	i->2	m->2	
mtala	d->1	r->1	
mtale	n->8	t->1	
mtals	p->1	r->1	
mtand	e->1	
mtank	a->1	
mtar 	u->1	
mtas 	i->1	
mtat 	r->1	
mte F	o->1	
mte b	e->1	
mte d	e->1	
mte h	a->1	
mte k	v->1	
mte p	e->1	u->1	
mte r	a->6	
mte v	å->1	
mtede	l->2	
mtid 	b->1	e->1	f->4	s->1	
mtid,	 ->3	
mtid.	.->1	D->2	M->1	N->1	T->1	
mtid:	 ->1	
mtida	 ->22	
mtide	n->64	
mtidi	g->67	
mtids	d->1	f->1	i->1	o->1	
mtiel	f->1	
mtio 	å->1	
mtioe	l->1	
mtion	,->1	.->1	
mtlig	a->25	
mtnin	g->1	
mton 	m->2	o->1	p->1	s->1	
mträd	a->2	
mts a	v->2	
mts i	 ->1	
mtsam	,->1	
mtvin	g->2	
mtyck	e->6	
mtänk	t->1	
mtåli	g->1	
muggl	i->1	
mula 	ö->1	
mulan	s->4	
mulat	i->1	o->2	
muler	a->20	i->6	
mull,	 ->1	
multi	e->3	l->1	n->5	
mum -	 ->1	
mum a	v->1	
mum m	i->1	
mum p	å->1	
mun.D	e->1	
munal	a->2	p->1	
muner	 ->7	n->2	s->1	
munic	e->2	
munik	a->16	
munis	m->1	
munit	e->1	
muntl	i->8	
muntr	a->21	
murar	 ->1	
mus e	n->1	
mus-b	e->1	
musik	 ->2	e->2	
musse	l->2	
mussl	a->1	
mutfo	r->1	
mutor	 ->1	
mutsa	r->1	t->1	
mutsi	g->1	
mvand	l->5	
mverk	a->3	s->1	
mvete	n->1	
mvets	s->1	
mvikt	;->1	e->1	
mvill	k->3	
mvist	,->1	
mväg 	f->1	
mväge	n->1	
mvälv	a->1	n->3	
mvänd	 ->3	a->1	
mvänt	 ->1	
mvärd	a->1	
mväxl	a->1	
mycke	n->2	t->450	
myggo	r->1	
myllr	a->1	
mynda	r->1	
myndi	g->161	
mynna	 ->1	r->1	
mytis	k->1	
mán, 	a->1	
mädel	s->1	
mäkta	 ->1	
mäkti	g->2	
mäla 	d->1	v->1	
mälan	 ->1	
mälda	 ->1	
mäler	.->1	
mälni	n->12	
mäls 	m->1	t->1	
mält 	s->1	
mältn	i->1	
män a	c->1	t->1	
män d	e->2	
män e	l->1	t->1	
män f	e->1	r->1	ö->2	
män g	e->1	i->2	
män h	a->1	
män i	 ->4	n->1	
män l	ä->1	
män n	ä->1	
män o	c->11	m->2	
män p	o->1	å->2	
män r	a->2	
män s	k->2	o->9	å->1	
män t	i->4	
män u	t->2	
män å	k->6	
män, 	e->1	
män.I	n->1	
män.J	a->1	
män.T	y->1	
mändr	i->3	
mängd	 ->14	e->8	
mängi	l->1	
mänhe	t->47	
mänie	n->1	
männa	 ->39	
männe	 ->1	n->28	
männi	s->93	
männy	t->2	
mäns 	f->1	p->1	s->2	
mänsk	l->42	
mänt 	a->2	g->1	h->1	i->3	k->1	m->3	p->1	s->2	t->1	u->1	
mänt,	 ->1	
märka	 ->4	
märkb	a->3	
märke	 ->7	l->5	n->2	r->4	t->1	
märkl	i->4	
märkn	i->13	
märks	 ->1	a->53	
märkt	 ->14	.->1	a->17	
märre	 ->1	
märta	r->1	
märts	a->1	
mässi	g->31	
mästa	r->2	
mäta 	d->1	s->1	
mätar	e->1	
mätas	 ->1	
mäter	 ->1	
mätig	t->1	
mätta	 ->1	
mätte	 ->1	s->1	
må Eu	r->1	
må an	m->1	
må be	f->1	
må bl	o->1	
må ek	o->1	
må fa	m->1	
må fr	å->1	
må fö	r->2	
må ha	 ->1	
må he	t->1	
må lä	n->2	
må me	d->2	
må mä	n->1	
må mö	j->1	
må oc	h->33	
må pl	a->1	
må rå	d->1	
må sp	r->1	
må st	a->2	e->1	u->1	
må va	r->1	
må åt	g->1	
må, m	e->1	
må, s	å->1	
må.De	n->1	
måend	e->2	
måför	e->6	
måga 	a->11	b->1	g->1	i->3	o->1	s->2	
måga,	 ->2	
måga.	O->2	
mågan	 ->5	,->3	
mågrä	l->1	
måhän	d->5	
mål (	B->1	
mål 1	 ->2	,->2	-->11	.->1	
mål 2	 ->5	,->1	-->3	.->1	
mål 5	b->2	
mål a	t->2	v->1	
mål b	e->2	
mål e	n->1	
mål f	i->1	ö->19	
mål g	å->1	
mål h	e->1	i->1	
mål i	 ->5	
mål j	a->1	
mål l	i->1	
mål n	å->1	
mål o	c->5	m->3	
mål p	å->2	
mål r	ö->1	
mål s	k->1	o->13	ä->1	
mål t	i->1	
mål u	p->2	
mål ä	r->4	
mål, 	R->1	f->2	g->1	h->1	m->2	n->1	o->1	p->1	s->5	u->1	
mål-2	-->1	
mål.B	ä->1	
mål.D	e->2	ä->1	
mål.E	t->1	
mål.F	r->1	
mål.H	e->2	
mål.I	 ->2	
mål.J	a->1	
mål.K	u->1	
mål.M	a->1	e->1	
mål.N	ä->2	
mål.Ä	v->1	
mål: 	a->1	
målar	f->1	
målen	 ->12	.->2	s->1	
målet	 ->21	,->2	.->5	
målig	a->1	
målin	r->4	
målme	d->1	
målsd	o->1	
målse	n->2	
målss	i->1	
målsä	t->17	
mån b	i->1	
mån d	e->3	r->1	ä->1	
mån f	ö->11	
mån h	a->1	
mån l	i->1	
mån o	m->1	
mån s	a->1	å->1	
mån, 	f->1	
måna 	o->3	
månad	 ->7	,->2	.->3	e->58	s->1	
månda	g->3	
månde	.->1	
måner	 ->1	.->1	
många	 ->137	,->2	.->2	
mångf	a->15	u->1	ä->1	
mångs	i->3	
månin	g->4	
månsp	a->1	
mår.H	e->1	
mår.L	a->1	
mårig	t->1	
mårsp	e->1	r->1	
måska	l->1	
måste	 ->693	,->3	
måt i	 ->5	
måt m	e->2	o->1	
måt o	c->2	
måt p	å->1	
måt v	e->1	
måt, 	i->1	m->2	
måt.D	a->1	e->1	ä->1	
måt.F	r->1	
måt.H	e->1	
måt.J	a->1	
måt.V	a->1	
måtgä	r->1	
mått 	a->1	
mått.	D->1	
måttf	u->1	
måtto	 ->2	
mé oc	h->2	
mé pe	r->1	
méavt	a->1	
mékon	v->1	
mén o	c->1	
mén.W	o->1	
més R	u->1	
möble	r->2	
möda 	o->2	s->1	
mödos	a->1	
mödra	r->1	
mögel	m->1	
mögna	 ->1	
möjli	g->307	
mönst	e->2	
mör s	o->1	
mör v	i->1	
mörda	d->2	n->1	r->1	t->1	
mörk 	d->1	
mörkl	ä->1	
mösso	r->1	
möta 	d->7	e->1	m->1	v->1	
möte 	d->1	i->4	k->1	m->4	o->1	p->1	s->1	
möten	 ->2	a->2	
möter	 ->40	!->14	,->7	.->1	n->24	s->1	
mötes	 ->1	.->1	g->3	
mötet	 ->19	.->2	
möts 	a->1	m->1	
mötte	s->1	
möver	 ->1	,->1	
n "Eu	r->1	
n "Lo	t->1	
n "Ti	b->2	
n "de	n->1	
n "dö	d->1	
n "en	 ->1	
n "eu	r->2	
n "he	r->1	
n "no	r->1	
n "re	s->2	
n "sp	e->1	
n "ut	v->1	
n "åt	e->1	
n (14	0->2	
n (19	9->1	
n (A5	-->5	
n (B5	-->2	
n (CE	N->2	
n (EI	F->1	
n (FU	F->1	
n (H-	0->21	
n (IM	O->1	
n (KO	M->1	
n (el	l->1	
n (fo	r->1	
n (fö	r->2	
n (in	f->1	
n (ma	i->1	
n (oc	h->1	
n (så	s->1	
n , b	o->1	
n - "	d->1	
n - '	V->1	
n - 2	,->1	
n - 6	 ->1	
n - A	l->1	
n - R	i->1	
n - a	l->1	t->3	
n - b	e->1	ö->1	
n - d	e->9	
n - e	f->1	k->1	l->1	n->1	t->1	x->1	
n - f	r->1	ö->2	
n - h	a->3	u->1	ä->1	
n - i	 ->2	n->1	
n - j	a->2	
n - l	i->2	
n - m	e->2	å->1	
n - n	å->1	
n - o	c->8	
n - s	e->1	k->1	o->4	
n - t	r->1	ä->1	
n - u	t->2	
n - v	a->1	e->1	i->1	
n - Ö	s->1	
n - ä	v->3	
n - ö	v->1	
n 1 j	a->5	u->1	
n 1 m	a->2	
n 1 o	c->2	
n 1 p	r->2	
n 1 s	e->1	
n 1, 	4->1	
n 10 	j->1	p->1	
n 100	 ->4	
n 105	 ->1	
n 11 	j->2	
n 12/	9->3	
n 124	4->2	
n 126	0->1	
n 13 	f->1	j->1	o->1	
n 13,	 ->1	
n 14 	f->5	o->1	s->1	
n 15 	o->1	s->1	
n 150	 ->1	
n 16 	o->1	r->1	
n 17 	d->1	m->1	o->1	
n 17,	 ->1	
n 18 	d->1	m->1	n->3	
n 19 	m->1	
n 191	7->1	
n 194	5->1	
n 196	7->4	9->1	
n 197	7->1	
n 198	2->1	6->1	9->1	
n 199	0->1	1->2	2->1	3->5	4->2	5->4	6->3	7->5	8->3	9->4	
n 2 d	e->1	
n 2 o	c->1	
n 2, 	1->1	
n 20 	å->1	
n 200	0->16	
n 21 	j->1	s->1	
n 23 	d->1	
n 24 	o->1	
n 26 	n->1	o->1	p->1	
n 28 	j->1	
n 29,	 ->1	
n 3 f	e->1	
n 3 j	a->1	
n 3 m	a->1	
n 3 o	k->1	
n 3, 	7->1	
n 3,8	 ->1	
n 30 	j->1	o->1	p->1	
n 31 	j->1	m->1	o->1	
n 34.	1->1	
n 38 	o->1	
n 39,	 ->1	
n 4 e	n->1	
n 4 j	u->2	
n 4, 	1->2	
n 5 0	0->2	
n 5 o	k->1	
n 50-	t->1	
n 520	 ->1	
n 57,	5->1	
n 6 d	e->1	
n 7 d	e->1	
n 7 o	c->1	
n 79/	4->1	
n 8 o	c->2	
n 89 	t->1	
n 9 d	e->1	
n 9 f	e->1	
n 90 	p->1	
n 95 	t->1	
n ABB	 ->1	
n ABC	 ->1	
n ADR	)->1	
n Act	.->1	
n Afr	i->1	
n Alb	a->1	
n Alt	e->2	
n Amo	k->1	
n Ams	t->5	
n Ann	a->1	
n Ari	 ->1	
n Ata	t->2	
n Aut	o->1	
n BSE	-->1	
n Bar	a->2	
n Bas	k->1	
n Bel	g->1	
n Ber	g->2	t->1	
n Boe	t->1	
n Bon	d->1	
n Bre	t->1	
n Bro	k->2	
n Bru	n->1	
n Bry	s->1	
n CEN	 ->2	,->1	:->1	
n Can	a->1	
n Cas	a->1	
n Cen	t->1	
n Cha	m->1	
n Cre	s->2	
n Dal	a->1	
n Dam	 ->2	
n Dan	m->1	
n De 	G->1	P->1	g->4	
n Dui	s->1	
n EG-	d->2	k->1	
n EKS	G->1	
n EMU	-->1	
n EU 	s->1	
n EU,	 ->1	
n EU-	m->1	
n EU:	s->2	
n EU?	H->1	
n Eie	c->1	
n En 	a->1	
n Enl	i->2	
n Eri	k->5	t->1	
n Eur	o->50	
n FEO	 ->1	
n FMI	 ->1	
n FN,	 ->1	
n Flo	r->4	
n Fol	k->1	
n Fon	t->1	
n Fra	n->2	
n För	e->2	
n GUE	/->1	
n Gal	i->1	
n Gar	g->1	
n Gaz	a->1	
n Gol	a->1	
n Gor	s->1	
n Gra	ç->1	
n Gre	k->1	
n Gru	p->1	
n Göt	e->1	
n Hai	d->2	
n Har	 ->2	
n Hel	s->2	
n Hul	t->23	
n I -	 ->1	
n I o	c->1	
n IMO	:->1	
n IRA	 ->1	
n IX,	 ->1	
n Imb	e->2	
n Ind	i->1	
n Int	e->2	
n Isa	b->2	
n Isr	a->12	
n Jac	o->1	q->1	
n Jap	a->1	
n Jor	d->1	
n Jug	o->1	
n Jun	k->1	
n Kal	e->2	
n Kar	l->2	t->1	
n Kin	a->3	n->1	
n Koc	h->4	
n Kom	m->1	
n Kor	e->1	
n Kos	o->1	
n Kyo	t->2	
n Köl	n->1	
n Köp	e->1	
n Lan	g->3	
n Lea	d->1	
n Lis	s->1	
n Loi	r->1	
n Loy	o->1	
n Mar	s->1	
n Min	u->1	
n Nat	i->3	o->2	
n Nie	l->1	
n Noi	r->1	
n OSS	E->1	
n PPE	-->2	
n PR-	e->1	
n PSE	)->1	
n Pal	e->2	
n Par	i->1	
n Pla	t->1	
n Pol	e->1	
n Por	t->4	
n Pro	d->6	v->1	
n Ran	d->2	
n Red	i->2	
n Rot	t->1	
n Rov	e->2	
n SPÖ	 ->1	
n SS 	o->1	
n Sam	m->3	
n Sch	e->1	u->1	
n Seb	a->1	
n Sha	r->2	
n Sol	a->1	
n Syd	k->1	
n Syr	i->4	
n São	 ->1	
n Tam	m->4	
n Ter	r->1	
n The	a->1	
n Tot	a->1	
n Tys	k->4	
n UNI	F->1	
n USA	.->1	
n Uni	o->2	
n VII	I->2	
n Val	d->3	
n Vel	z->1	
n Ven	d->1	
n Viv	i->1	
n Wal	e->1	
n Wie	l->3	n->1	
n Wog	a->18	
n Wur	t->1	
n XXV	I->1	
n a p	r->1	
n abs	o->3	u->1	
n acc	e->15	
n ade	k->1	
n adm	i->5	
n adr	i->1	
n adv	o->1	
n age	r->3	
n agr	a->1	
n akt	i->2	u->9	ö->1	
n alb	a->2	
n ald	r->4	
n all	 ->1	a->9	d->3	e->2	i->2	m->22	r->1	s->2	t->20	v->3	
n amb	i->2	
n ame	r->3	
n an 	p->1	
n ana	 ->1	l->10	
n anb	u->1	
n and	a->6	e->2	r->65	
n ang	e->3	r->2	å->6	
n ani	n->3	
n anl	e->22	ä->1	ö->1	
n anm	ä->5	
n ann	a->40	
n ano	r->2	
n anp	a->1	
n ans	e->17	j->2	k->1	l->3	p->1	t->4	v->15	å->2	ö->2	
n ant	a->6	i->5	o->2	
n anv	i->1	ä->16	
n app	l->2	
n ara	b->2	
n arb	e->22	
n ark	i->1	
n art	e->1	i->4	
n asp	e->7	
n asy	l->1	
n att	 ->426	,->1	:->1	i->1	
n auk	t->2	
n aut	o->1	
n av 	-->1	1->1	2->1	A->1	B->1	E->13	G->1	K->5	L->1	O->2	S->1	W->1	a->22	b->16	c->2	d->100	e->26	f->50	g->9	h->3	i->4	j->4	k->29	l->10	m->22	n->4	o->13	p->22	r->13	s->35	t->9	u->18	v->17	Ö->2	ä->1	å->7	ö->4	
n av.	E->1	J->1	
n avb	r->7	
n avd	e->1	
n avf	a->3	ö->3	
n avg	e->2	i->2	j->1	å->1	ö->9	
n avi	s->2	
n avl	e->2	ä->1	
n avs	e->10	i->6	k->3	l->22	p->2	t->2	
n avt	a->1	
n avv	i->3	ä->2	
n axe	l->1	
n bad	a->1	
n bak	g->3	o->1	
n bal	a->8	
n ban	a->1	b->1	k->1	t->1	
n bar	a->23	
n bea	k->6	r->1	
n bed	r->2	ö->12	
n bef	a->1	i->6	o->9	ä->1	
n beg	r->12	ä->13	
n beh	a->3	o->1	å->2	ö->18	
n bek	l->5	r->9	ä->1	
n bel	a->4	g->4	
n bem	ä->3	ö->3	
n ben	e->1	
n ber	 ->2	e->7	i->1	o->3	ä->4	ö->3	
n bes	e->1	k->5	l->5	p->2	t->18	v->5	y->1	
n bet	a->8	o->4	r->12	t->1	v->1	y->14	ä->2	
n beu	n->1	
n bev	a->1	i->5	
n bib	e->1	
n bid	r->13	
n bil	 ->6	,->1	.->1	a->3	d->4	e->1	i->4	s->2	t->1	
n bin	d->1	
n bio	l->2	
n bit	t->2	
n bla	n->8	
n ble	k->1	v->3	
n bli	 ->8	r->14	v->1	x->1	
n blo	c->1	m->1	t->1	
n boe	n->1	
n bok	 ->3	
n bom	b->1	
n bon	d->2	
n bor	d->13	t->4	
n bos	n->1	ä->1	
n bot	a->2	t->2	
n bra	 ->11	n->3	
n bre	d->6	t->1	
n bri	s->10	t->4	
n bro	 ->1	k->1	m->1	r->1	t->3	
n bru	n->1	
n brä	n->2	
n bud	d->1	g->12	
n byg	g->3	
n byr	å->6	
n byt	a->1	t->1	
n bär	 ->4	a->1	
n bäs	t->6	
n bät	t->17	
n båd	a->1	e->2	
n bör	 ->38	j->18	
n cen	t->10	
n cer	t->1	
n cha	n->6	
n che	c->1	f->1	
n cho	c->1	
n con	d->1	
n cor	p->1	
n cos	t->4	
n dag	 ->7	.->1	e->4	l->1	o->7	s->2	
n dam	 ->1	
n dan	s->7	
n de 	1->1	a->4	b->4	d->3	e->7	f->4	g->1	h->2	i->6	k->4	m->6	n->7	o->16	p->1	s->6	t->5	u->4	v->4	ö->1	
n dea	d->1	
n deb	a->30	
n dec	e->8	
n def	i->6	
n deg	e->1	
n del	 ->55	,->2	.->1	a->5	e->5	l->1	s->1	t->3	v->2	
n dem	 ->4	.->1	o->16	
n den	 ->87	.->1	n->15	
n dep	a->1	
n der	 ->8	a->3	
n des	s->19	
n det	 ->162	,->2	.->1	a->4	t->26	
n dia	l->7	
n dik	t->2	
n dir	e->8	
n dis	k->17	
n dit	 ->1	
n div	e->1	
n dju	p->7	
n djä	r->1	
n doc	k->3	
n dog	m->1	
n dok	u->2	
n dom	 ->2	a->1	i->1	s->5	
n dra	 ->5	b->3	r->1	
n dri	v->2	
n dro	p->1	
n dru	c->1	n->2	
n dry	g->1	
n drö	j->2	
n dub	b->1	
n dum	h->1	
n dun	a->1	
n dyk	a->1	
n dyn	a->1	
n där	 ->38	,->1	.->1	e->5	f->5	i->1	m->5	p->1	
n då 	E->2	b->2	f->1	i->1	k->2	o->1	p->2	s->3	v->2	
n dål	i->1	
n dåv	a->1	
n död	f->1	s->1	
n döl	j->2	
n döm	a->1	d->1	
n döp	a->1	e->1	t->1	
n dör	 ->1	r->2	
n eff	e->24	
n eft	e->31	
n ege	n->22	
n egn	a->4	
n ej 	a->2	
n eko	l->5	n->50	
n ele	f->1	k->2	
n ell	e->36	
n elo	g->2	
n eme	l->6	
n emi	g->1	
n en 	a->6	b->5	c->1	d->3	e->3	f->7	g->29	h->3	i->4	j->1	k->4	l->5	m->9	n->3	o->4	p->4	r->2	s->13	t->9	u->2	v->2	ä->1	ö->2	
n ena	 ->11	d->1	s->2	
n enb	a->5	
n end	a->31	
n ene	r->4	
n eng	a->2	e->6	
n enh	e->13	ä->4	
n enk	e->2	l->2	
n enl	i->10	
n eno	r->9	
n ens	i->4	k->7	t->1	
n ent	u->1	
n env	i->1	
n epo	k->1	
n er 	p->1	v->1	
n er,	 ->1	
n era	 ->1	
n erb	j->3	
n erf	a->2	
n erh	ö->2	
n eri	n->1	
n erk	ä->6	
n ers	ä->3	
n ert	 ->2	
n etn	i->3	
n ett	 ->52	
n eur	o->145	
n eve	n->4	
n ex 	a->1	
n exa	k->1	m->2	
n exe	m->1	
n exi	s->5	
n exk	l->1	
n exp	a->1	e->6	l->1	o->2	
n ext	e->2	r->5	
n fak	t->7	
n fal	l->4	
n fan	n->1	t->1	
n far	a->3	l->2	t->4	
n fas	c->1	t->11	
n fat	t->9	
n fed	e->2	
n fel	 ->1	b->1	s->1	
n fem	 ->4	t->3	
n fic	k->3	
n fil	o->1	
n fin	 ->1	a->4	l->1	n->32	s->1	
n fjo	r->1	
n fjä	r->6	
n fla	g->3	
n fle	r->5	x->3	
n fli	t->1	
n flo	d->1	
n fly	g->1	
n fok	u->1	
n fol	k->2	
n fon	d->4	
n for	m->8	s->2	t->23	
n fra	m->35	n->12	
n fre	d->8	s->1	
n fri	 ->2	,->1	a->10	
n fro	d->2	
n fru	,->1	k->3	
n fry	s->1	
n frä	m->4	
n frå	g->82	n->77	
n ful	l->12	
n fun	d->3	g->5	k->4	n->1	
n fus	i->1	
n fyl	l->1	
n fyr	a->2	t->1	
n fys	i->2	
n fäl	l->1	
n fär	d->1	
n fäs	t->4	
n få 	d->3	e->6	f->2	k->1	l->1	m->1	n->1	s->2	t->2	v->1	
n få,	 ->1	
n fån	g->1	
n får	 ->24	
n fås	 ->1	
n fåt	t->1	
n föd	e->2	
n föl	j->6	l->2	
n fön	s->1	
n för	 ->464	,->1	a->5	b->19	d->15	e->66	f->4	g->1	h->9	k->12	l->7	m->5	n->11	o->7	p->2	r->14	s->103	t->8	u->12	v->13	ä->9	
n gam	l->7	m->1	
n gan	s->7	
n gar	a->20	
n gav	 ->1	
n ge 	d->3	e->5	g->1	i->1	j->1	o->2	p->1	u->2	
n ged	i->1	
n gem	e->100	
n gen	a->1	e->3	o->44	t->3	
n geo	s->1	
n ger	 ->6	
n ges	 ->2	
n get	t->2	
n gic	k->2	
n gig	a->2	
n gil	t->2	
n giv	a->1	e->2	
n gjo	r->14	
n gla	d->1	
n gle	s->1	
n glo	b->3	
n glä	d->9	
n gnu	t->2	
n god	 ->6	a->7	k->11	t->11	
n gra	d->4	n->10	v->1	
n gre	k->5	
n gri	p->1	
n gru	n->19	p->37	v->1	
n grä	n->3	
n grö	n->1	
n gum	m->1	
n gyn	n->1	
n gäl	l->26	
n gär	n->1	
n gå 	f->2	i->3	o->1	s->1	u->1	
n gån	g->56	
n går	 ->9	,->1	
n gåt	t->1	
n gör	 ->18	a->29	s->4	
n ha 	d->1	e->2	h->1	k->1	m->1	s->2	t->1	u->1	ä->1	
n had	e->17	
n haf	t->7	
n hal	v->8	
n ham	m->1	n->3	
n han	 ->5	d->18	s->2	t->1	
n har	 ->312	,->2	.->1	:->1	?->1	m->4	
n hav	e->1	
n heb	r->1	
n hej	d->2	
n hel	 ->11	a->5	h->12	l->3	t->12	
n hem	b->1	s->2	v->1	
n her	r->1	
n hin	d->2	
n his	t->3	
n hit	t->8	
n hjä	l->9	r->1	
n hon	 ->1	
n hop	p->10	
n hor	d->1	
n hos	 ->10	
n hot	a->4	e->1	f->1	
n hun	d->2	
n hur	 ->8	
n huv	u->7	
n hyp	o->1	
n hys	e->1	
n häl	s->1	
n häm	n->2	
n hän	d->5	f->1	g->1	s->6	v->9	
n här	 ->77	.->1	l->1	r->1	
n häv	d->6	
n hål	l->17	
n hår	d->4	
n hög	 ->5	a->4	e->3	n->1	r->4	s->7	t->2	
n höj	d->3	n->1	
n hör	 ->4	.->1	
n i A	B->1	f->1	m->2	v->1	
n i B	N->1	e->2	i->1	o->1	r->4	
n i C	e->1	u->1	
n i D	D->1	u->1	
n i E	U->3	u->31	
n i F	o->1	r->1	ö->3	
n i G	a->1	r->2	u->1	
n i H	a->1	e->2	
n i I	C->1	r->2	s->1	t->1	
n i K	a->2	o->10	y->1	
n i L	a->2	e->1	i->1	o->2	u->3	
n i M	a->1	e->7	
n i N	e->1	o->1	
n i O	m->1	
n i P	a->1	
n i R	a->1	y->1	
n i S	a->1	e->2	k->1	r->1	t->5	y->2	
n i T	a->1	h->2	i->2	u->2	y->2	
n i V	a->1	ä->1	
n i W	a->2	
n i a	l->11	n->5	r->4	v->1	
n i b	e->7	i->2	r->1	u->1	å->1	
n i c	e->2	
n i d	a->20	e->83	i->2	o->1	
n i e	f->1	n->14	r->3	t->9	u->1	
n i f	a->2	e->1	l->2	o->12	r->30	ö->11	
n i g	e->1	l->1	r->1	å->5	
n i h	a->5	e->3	i->1	
n i i	c->1	n->3	
n i j	u->2	
n i k	a->1	n->1	o->5	v->2	
n i l	a->3	i->1	j->2	y->1	å->1	
n i m	a->1	e->9	i->7	o->6	å->7	
n i n	ä->1	
n i o	k->1	l->1	m->5	
n i p	a->4	e->2	l->3	o->1	r->6	
n i r	a->1	e->5	i->2	å->6	
n i s	a->7	e->3	i->21	j->6	l->4	t->11	y->1	ä->1	å->2	
n i t	a->1	o->2	r->1	v->1	
n i u	n->11	r->1	t->7	
n i v	a->7	e->1	i->5	ä->2	å->11	
n i z	o->1	
n i Ö	s->14	
n i ä	n->1	r->1	
n i å	r->2	t->1	
n i ö	v->1	
n i, 	u->1	
n ibl	a->1	
n ick	e->4	
n ide	n->4	o->2	
n idé	 ->3	n->1	
n ifr	å->3	
n ign	o->1	
n ihä	r->1	
n ihå	g->1	
n ill	a->1	e->1	o->1	
n imp	u->1	
n in 	i->1	
n inb	e->3	j->1	
n inc	i->1	
n ind	e->1	i->2	u->4	
n ine	f->2	
n inf	o->16	r->1	ö->16	
n ing	e->1	r->1	å->5	
n inh	e->1	ä->2	
n ini	t->1	
n ink	l->1	ö->1	
n inl	e->8	ä->1	
n inn	a->6	e->22	o->1	
n ino	m->50	
n inr	e->62	i->6	ä->2	
n ins	a->3	e->4	i->2	k->2	l->1	t->17	
n int	e->240	o->1	r->7	y->2	
n inv	e->3	ä->1	å->1	
n ira	k->1	
n irl	ä->2	
n isr	a->11	
n ist	ä->1	
n ita	l->5	
n jag	 ->126	,->2	.->1	a->1	
n jak	t->2	
n jan	u->1	
n ju 	i->1	o->1	u->1	ä->1	
n jub	l->1	
n jul	 ->1	i->1	
n jun	i->1	
n jur	i->7	
n jus	t->15	
n jäm	f->3	l->2	n->1	s->1	v->1	
n kab	a->1	
n kal	l->5	
n kam	,->1	m->1	p->3	r->1	
n kan	 ->132	,->1	s->10	
n kap	a->1	
n kar	r->1	t->1	
n kas	k->1	t->1	
n kat	a->15	o->2	
n ked	j->1	
n kel	t->1	
n kin	e->1	
n kl.	 ->11	1->1	
n kla	g->2	r->14	s->3	
n kli	m->1	
n kna	p->3	
n koa	l->4	
n kol	l->29	o->1	
n kom	 ->7	b->1	m->238	p->12	
n kon	c->4	f->6	k->30	s->24	t->20	v->1	
n kop	i->1	p->2	
n kor	r->1	t->4	
n kos	t->13	
n kra	f->11	
n kri	n->2	s->2	t->8	
n krä	n->5	v->15	
n krö	n->1	
n kul	t->11	
n kun	d->6	n->10	s->2	
n kur	s->1	
n kva	l->3	n->1	
n kvi	n->4	
n kvo	t->6	
n kyl	a->1	
n käl	l->3	
n kän	n->5	s->11	
n kär	a->1	n->1	
n kön	e->3	
n kör	a->1	
n lad	e->3	
n lag	s->12	t->7	
n lan	d->1	
n lar	m->1	
n law	.->1	
n led	a->16	e->4	
n leg	a->1	i->1	
n lev	a->2	
n lib	e->4	
n lid	e->1	
n lig	g->9	
n lik	a->3	n->3	r->2	s->1	t->1	v->1	
n lin	b->1	d->2	j->2	
n lit	a->1	e->10	
n liv	s->4	
n log	i->2	
n lok	a->8	
n lov	a->1	o->1	v->1	
n luc	k->1	
n lyc	k->8	
n lyd	e->1	
n lys	a->2	s->2	
n läg	e->1	g->16	r->4	
n läm	n->4	p->3	
n län	d->7	g->4	
n lär	a->2	
n läs	a->1	e->4	
n lät	t->4	
n låg	 ->1	a->1	t->1	
n lån	g->20	
n låt	 ->1	a->1	e->1	
n löj	e->1	
n lök	m->1	
n lön	s->1	
n löp	e->1	
n lös	a->5	n->15	
n m.m	.->1	
n mag	e->1	n->1	
n maj	 ->1	o->5	
n mak	t->5	
n mal	t->1	
n man	 ->47	
n mar	g->2	k->15	
n mas	k->2	o->1	s->3	
n max	i->2	
n med	 ->133	a->2	b->5	d->3	e->3	f->8	g->2	i->1	k->2	l->55	v->2	
n mel	l->41	
n men	 ->8	,->1	a->1	i->21	
n mer	 ->19	.->1	a->3	v->1	
n mes	t->2	
n met	o->5	
n mil	d->1	i->1	j->15	s->1	
n min	 ->7	d->6	i->9	o->3	s->16	u->2	
n mis	s->11	t->1	ä->1	
n mit	t->1	
n mod	e->14	
n mon	e->2	o->1	
n mor	a->1	g->1	
n mot	 ->34	i->2	s->7	t->3	v->1	å->1	
n mul	t->1	
n mun	t->3	
n myc	k->69	
n myn	d->12	
n män	g->9	n->4	s->2	
n mär	k->3	
n mät	a->2	
n må 	h->2	
n måh	ä->1	
n mål	 ->1	e->1	m->1	
n mån	 ->4	,->1	a->4	g->5	
n mås	t->139	
n möj	l->21	
n mör	d->1	k->1	
n möt	a->2	e->1	t->1	
n nat	i->20	t->1	u->15	
n ned	e->4	g->1	m->1	s->1	
n neg	a->5	
n neu	t->1	
n ni 	b->2	d->1	f->1	h->2	o->1	s->4	v->2	
n nio	n->1	
n niv	å->3	
n nog	g->1	
n nol	l->1	
n nom	i->2	
n nor	d->2	m->3	
n not	e->5	
n nu 	b->1	g->3	h->3	i->1	k->2	l->1	m->3	n->1	o->1	s->6	t->2	u->1	v->2	ä->1	
n nu,	 ->1	
n num	e->1	
n nuv	a->16	
n ny 	b->1	e->1	f->3	i->1	k->5	l->1	m->1	o->1	p->1	r->1	s->5	t->1	u->1	v->2	
n nya	 ->37	s->1	
n nyc	k->2	
n nye	 ->1	
n nyh	e->1	
n nyl	i->5	
n nyn	a->1	
n nys	s->4	
n nyt	t->8	
n näm	l->2	n->13	
n när	 ->32	a->3	h->1	m->5	v->1	
n näs	t->2	
n nå 	d->1	e->1	f->1	
n nåb	a->2	
n någ	o->30	r->6	
n nöd	s->1	v->14	
n nöj	a->1	
n nöt	.->1	
n oac	c->2	
n oan	s->2	
n oav	b->1	s->1	
n oba	l->1	
n obe	r->21	
n obl	i->5	
n och	 ->582	,->3	
n ock	s->96	u->1	
n oeg	e->1	
n oen	i->1	
n oer	h->2	
n ofa	n->1	
n off	e->25	i->1	
n oft	a->2	
n ofö	r->5	
n ohä	m->1	
n okl	a->2	
n oko	n->1	
n okä	n->2	
n oli	k->8	
n olj	a->1	e->1	
n oly	c->7	
n om 	"->1	-->1	1->1	3->1	4->1	A->1	B->1	C->1	E->6	K->3	M->2	T->2	a->33	b->10	c->1	d->72	e->21	f->22	g->3	h->13	i->15	j->16	k->26	l->8	m->13	n->4	o->4	p->4	r->20	s->23	t->9	u->3	v->28	Ö->1	å->2	ö->4	
n om"	.->1	
n om,	 ->4	
n om.	J->1	N->1	
n omI	.->1	
n omb	e->1	
n omd	e->1	
n ome	d->5	
n omf	a->13	o->1	
n omi	s->1	
n omm	ö->1	
n omo	r->1	
n omp	l->1	r->4	
n omr	ö->7	
n oms	o->1	t->2	v->1	ä->1	
n omv	a->1	ä->5	
n omö	j->4	
n ond	 ->1	
n one	-->1	
n onö	d->2	
n ope	r->2	
n opp	o->2	
n opt	i->2	
n ord	 ->1	e->4	f->2	l->1	n->10	v->1	
n org	a->7	
n ori	e->1	
n ork	a->1	
n orm	 ->1	
n oro	 ->19	a->4	n->1	v->1	
n ors	a->3	
n ort	,->1	
n orä	t->1	
n oss	 ->6	
n ota	c->1	
n oti	l->2	
n otj	ä->1	
n oum	b->2	
n oun	d->1	
n ova	n->2	
n ovi	l->3	
n oän	d->1	
n oön	s->1	
n oöv	e->2	
n p.g	.->1	
n pal	e->4	
n par	a->3	l->27	t->4	
n pas	s->2	
n ped	o->1	
n pek	a->2	
n pel	a->2	
n pen	n->1	
n per	 ->4	f->2	i->8	m->3	s->10	
n pet	i->1	
n pla	c->1	n->13	t->8	
n pli	k->1	
n plu	r->1	
n plö	t->2	
n poe	t->1	
n pol	e->2	i->55	
n poo	l->1	
n por	s->1	t->4	
n pos	i->15	
n pot	e->1	
n poä	n->2	
n pra	k->1	t->1	
n pre	c->3	l->1	m->1	s->9	
n pri	n->3	o->3	s->1	v->5	
n pro	b->3	c->6	d->13	f->2	g->2	p->1	t->1	v->2	
n pun	k->28	
n pur	i->1	
n pyr	a->1	
n på 	3->2	B->3	E->1	I->1	R->1	V->1	a->23	b->2	d->59	e->36	f->11	g->15	h->5	i->1	k->9	l->5	m->10	n->8	o->4	p->1	r->8	s->10	t->9	u->3	v->4	ä->1	å->3	ö->3	
n på:	 ->1	
n på?	.->1	
n påb	ö->1	
n påf	r->1	
n påg	i->1	å->4	
n påm	i->3	
n påp	e->6	
n pås	k->1	t->5	
n påt	a->2	
n påv	e->5	
n rad	 ->18	e->1	i->4	
n ram	 ->3	,->1	
n rap	p->11	
n ras	a->2	i->1	
n rat	i->1	
n rea	g->2	k->1	l->1	
n red	a->22	o->5	u->1	
n ree	l->3	
n ref	l->1	o->17	
n reg	e->31	i->33	l->2	
n rek	o->5	
n rel	a->2	e->1	i->2	
n rem	i->1	
n ren	 ->3	t->5	
n rep	u->1	
n res	e->1	o->16	p->12	t->1	u->9	
n rev	i->9	
n rig	h->1	
n rik	a->1	e->1	l->1	t->17	
n rim	l->3	
n ris	k->17	
n rol	l->11	
n ros	 ->1	
n run	d->1	t->1	
n rus	a->1	
n rys	k->1	
n räc	k->2	
n räd	d->2	s->2	
n räk	n->7	
n rät	a->1	t->47	
n råd	e->24	g->2	
n råg	a->1	
n réf	é->1	
n röd	a->1	g->1	
n rör	 ->2	a->3	
n rös	t->17	
n sad	e->17	
n sag	t->9	
n sak	 ->10	,->1	.->1	:->1	e->3	k->1	n->5	
n sam	a->1	e->1	h->2	m->16	o->8	s->1	t->18	
n san	n->5	
n sat	e->1	s->5	t->2	
n sce	n->1	
n sco	r->1	
n se 	a->1	e->1	f->1	h->1	i->1	o->1	t->4	u->1	v->1	
n sed	a->10	
n seg	 ->1	l->1	
n sek	t->2	
n sen	a->12	
n sep	a->1	
n ser	 ->11	b->7	i->1	
n set	t->2	
n sex	m->1	
n sif	f->1	
n sig	 ->9	n->3	
n sin	 ->4	a->6	e->1	
n sis	t->20	
n sit	t->5	u->18	
n sju	k->1	n->3	t->1	
n sjä	l->18	t->11	
n ska	d->4	f->1	l->162	m->4	n->3	p->14	r->1	t->2	
n ske	 ->2	r->3	
n ski	c->1	l->8	
n skj	u->3	
n sko	g->2	
n skr	i->7	o->2	ä->2	
n sku	g->1	l->71	
n sky	d->2	l->6	n->1	
n skä	r->3	
n skö	r->1	t->3	
n sla	g->4	
n slo	g->1	
n slu	m->5	t->17	
n slå	r->1	
n smi	d->1	
n smu	l->1	
n smä	d->1	r->1	
n små	 ->1	
n sna	b->6	r->15	
n sne	d->2	
n so 	f->1	
n soc	i->41	
n sol	i->6	
n som	 ->347	,->5	m->1	
n sor	t->6	
n spa	n->3	r->1	
n spe	c->10	g->1	l->7	t->1	
n spl	i->2	
n spo	n->1	
n spr	i->2	å->1	
n spä	r->1	
n sri	l->1	
n sta	b->3	d->10	n->3	r->16	t->24	
n sti	g->2	l->1	m->2	
n sto	p->3	r->54	
n str	a->11	i->8	u->18	ä->5	ö->1	
n stu	n->7	
n sty	r->4	
n stä	d->2	l->11	m->5	n->6	r->2	
n stå	n->9	r->15	
n stö	d->16	l->1	r->26	t->1	
n sub	s->2	
n suc	c->2	
n sum	m->1	
n sun	d->2	
n sup	r->1	
n suv	e->1	
n sva	g->2	r->4	
n sve	n->1	p->1	
n svå	r->3	
n syf	t->3	
n sym	b->3	
n syn	d->1	n->2	p->2	t->1	v->3	
n syr	i->4	
n sys	s->2	t->4	
n säg	a->15	e->9	s->1	
n säk	e->9	
n säl	l->2	
n sär	b->1	s->16	
n sät	t->5	
n så 	a->6	b->3	d->1	f->1	g->3	h->1	j->1	k->3	l->6	p->2	r->2	s->8	u->2	ä->3	ö->1	
n så,	 ->1	
n så:	 ->1	
n såd	a->47	
n såg	 ->1	
n såh	ä->1	
n sål	e->2	
n sån	g->1	
n sås	o->4	
n såv	ä->1	
n söd	r->2	
n sök	e->1	
n t.e	x->1	
n ta 	e->1	f->1	h->2	i->1	l->1	m->1	n->1	o->1	p->1	s->2	t->1	u->3	
n tac	k->10	
n tag	i->7	
n tal	a->28	m->1	
n tan	k->2	
n tap	p->1	
n tar	 ->10	
n tas	 ->4	k->1	
n tec	k->2	
n tek	n->9	
n ten	d->1	
n ter	a->1	r->3	
n tex	t->2	
n tib	e->4	
n tid	 ->10	e->1	i->19	n->1	p->2	s->10	
n til	l->316	
n tim	m->1	
n tio	 ->1	
n tit	t->6	
n tjä	n->8	
n tog	 ->4	
n tol	k->2	
n tom	 ->1	
n ton	 ->1	v->1	
n top	p->2	
n tot	a->11	
n tra	d->3	g->3	n->1	
n tre	 ->3	d->30	k->1	v->2	
n tro	 ->1	r->5	t->5	v->1	
n trä	d->2	f->1	t->1	
n trö	g->1	
n tuf	f->1	
n tun	g->5	
n tur	 ->5	,->1	k->3	
n tve	k->16	t->3	
n tvi	n->5	v->17	
n tvä	r->5	
n två	 ->7	
n tyc	k->5	
n tyd	l->15	
n tyg	e->1	
n tyn	a->1	g->2	
n typ	 ->4	e->1	
n tys	k->9	t->3	
n tyv	ä->6	
n tän	k->9	
n täv	l->1	
n und	a->3	e->72	r->1	v->3	
n ung	 ->1	
n uni	o->14	v->1	
n upp	b->3	d->1	e->4	f->29	g->12	h->2	l->1	m->14	n->11	r->9	s->14	t->4	v->2	
n ur 	E->1	b->1	d->1	e->1	s->1	
n urm	i->1	
n urs	p->4	ä->2	
n urv	a->1	
n ut,	 ->1	
n uta	n->18	
n utb	i->4	r->1	u->1	
n ute	s->3	
n utf	a->1	o->3	r->2	ö->6	
n utg	a->1	å->3	ö->9	
n uti	f->1	
n utj	ä->1	
n utk	o->1	
n utl	a->1	o->2	
n utm	a->5	ä->2	
n utn	y->6	
n utp	l->1	
n utr	e->1	ä->1	
n uts	a->1	e->1	k->18	t->6	ä->1	å->3	
n utt	a->9	j->2	r->5	
n utv	e->15	i->17	ä->2	
n utö	v->5	
n vad	 ->16	
n val	d->5	k->2	l->1	t->2	
n van	 ->3	h->1	l->2	
n var	 ->26	a->43	e->2	f->1	i->3	j->3	k->1	m->2	n->1	s->3	t->2	
n vat	t->1	
n vec	k->3	
n ved	e->2	
n vek	h->1	
n vem	 ->2	
n ver	i->1	k->40	
n vet	 ->7	e->11	t->2	
n vi 	a->9	b->15	d->2	e->1	f->10	g->3	h->12	i->15	k->11	l->2	m->16	o->2	r->2	s->12	t->2	u->4	v->5	y->1	ä->8	å->1	
n vi,	 ->1	
n vi.	V->1	
n vic	e->1	
n vid	 ->41	a->4	t->15	
n vif	t->1	
n vik	t->59	
n vil	j->10	k->4	l->42	
n vin	n->1	s->1	
n vis	a->19	s->32	u->1	
n vit	b->5	
n vol	u->1	
n vor	e->3	
n vri	d->1	
n vun	n->1	
n väc	k->2	
n väd	j->2	
n väg	 ->1	e->1	r->5	
n väl	 ->6	,->1	d->1	j->1	k->3	m->1	u->1	
n vän	 ->1	d->6	s->3	t->7	
n vär	d->5	l->2	s->1	
n väs	e->6	
n väv	n->1	
n väx	a->5	e->1	l->1	
n våg	e->1	
n vål	d->4	
n vår	 ->3	a->7	t->3	
n wal	e->1	
n web	b->1	
n ytt	e->7	r->1	
n zig	e->2	
n Öst	e->3	
n äga	 ->1	r->2	
n äge	r->1	
n ägn	a->4	
n ägt	 ->1	
n äls	k->1	
n än 	a->1	d->2	e->2	h->1	l->1	m->1	p->1	v->1	ä->1	
n änd	r->27	å->4	
n änn	u->10	
n änt	l->1	
n är 	-->1	E->1	P->1	a->33	b->31	d->39	e->34	f->25	g->5	h->6	i->18	j->4	k->7	l->8	m->14	n->9	o->10	p->4	r->4	s->18	t->5	u->5	v->12	y->1	ä->2	å->1	ö->4	
n är,	 ->3	
n är.	D->1	H->1	J->1	k->1	
n är:	 ->2	
n ära	n->1	
n ärl	i->1	
n äve	n->32	
n å a	n->1	
n å d	e->3	
n å e	n->4	
n åbe	r->1	
n åkl	a->8	
n åla	g->1	
n åld	e->2	
n ålä	g->1	
n år 	1->2	2->5	a->1	t->1	
n årl	i->1	
n åsi	k->22	
n åst	a->5	
n åsy	f->1	
n åt 	a->1	d->2	e->1	n->1	s->1	t->1	
n åta	r->1	
n åte	r->23	
n åtf	ö->3	
n åtg	ä->11	
n åtm	i->3	
n åts	k->1	
n ått	o->1	
n öde	s->1	
n öka	 ->2	.->1	d->14	r->5	t->1	
n ökn	i->9	
n öm 	t->1	
n öns	k->9	
n öpp	e->7	n->1	
n öre	g->1	
n öst	e->18	
n öve	r->74	
n övn	i->2	
n övr	i->4	
n! Al	l->2	
n! At	t->1	
n! Av	 ->1	f->1	
n! Be	s->1	t->1	
n! Da	g->1	
n! De	 ->1	n->4	t->25	
n! Dä	r->1	
n! Dí	e->1	
n! EU	 ->1	
n! En	d->1	
n! Er	t->1	
n! Eu	r->3	
n! Fr	a->1	u->1	å->1	
n! Få	r->1	
n! Fö	r->8	
n! Gr	u->2	
n! He	r->1	
n! I 	b->2	d->4	e->2	l->1	
n! In	t->1	
n! Ja	g->75	
n! Ko	m->4	n->1	
n! Li	k->1	
n! Lå	t->5	
n! Ma	n->1	
n! Mi	n->5	
n! Ni	 ->1	
n! Nu	 ->1	
n! Nä	r->4	
n! Ol	j->1	
n! Om	 ->1	
n! Pa	r->1	
n! Pr	i->1	
n! På	 ->1	s->1	
n! Re	g->1	
n! Ro	t->1	
n! Rå	d->2	
n! Sc	h->1	
n! Se	d->3	
n! Sk	u->1	
n! So	m->3	
n! St	r->1	
n! Ta	c->1	
n! Th	e->1	
n! Ti	l->4	
n! To	r->1	
n! Tr	o->1	
n! Un	d->2	
n! Ut	s->2	
n! Va	d->2	r->1	
n! Vi	 ->11	d->1	
n! Vå	r->2	
n! Än	n->1	
n! Äv	e->6	
n! Å 	P->1	k->1	s->1	
n! Ös	t->1	
n!Ams	t->1	
n!Den	 ->1	
n!Det	 ->2	
n!Eft	e->1	
n!En 	v->1	
n!Her	r->1	
n!Jag	 ->6	
n!Min	a->1	
n!När	 ->2	
n!Rös	t->1	
n!San	n->1	
n!Tac	k->1	
n!Til	l->1	
n!Und	e->1	
n!Vi 	h->1	ä->1	
n" al	d->1	
n" at	t->1	
n" et	c->1	
n" ge	m->1	
n" i 	A->1	
n" oc	h->1	
n" på	 ->1	
n" so	m->1	
n", "	s->1	
n", d	e->1	
n", o	c->1	
n", s	o->2	
n".De	 ->1	t->2	
n".Or	d->1	
n".Rå	d->1	
n) (K	O->2	
n) (S	E->1	
n) fö	r->1	
n) ha	r->1	
n) zo	n->1	
n)(Pa	r->2	
n), o	c->1	
n).De	 ->1	t->1	
n).He	r->1	
n)Jag	 ->1	
n)Näs	t->1	
n, "o	v->1	
n, 1 	p->1	
n, 10	,->1	
n, 15	,->1	
n, 19	9->1	
n, 50	0->1	
n, 8,	 ->1	
n, Am	o->2	
n, BN	I->1	
n, Be	l->1	r->2	
n, Br	e->1	
n, Cu	x->1	
n, Du	b->1	
n, Eu	r->2	
n, IV	 ->1	
n, Ir	l->1	
n, Jo	r->1	
n, Ka	r->1	z->1	
n, Ko	c->1	r->1	
n, Lo	m->1	r->1	
n, Ne	d->1	
n, Ol	y->1	
n, Pa	l->3	
n, Pe	i->1	
n, Ra	p->1	
n, Ro	t->1	
n, Sh	a->1	
n, Sl	o->1	
n, Sv	e->1	
n, To	t->1	
n, Ty	s->1	
n, Uz	b->1	
n, V 	-->1	
n, Vl	a->1	
n, Wi	e->1	
n, al	l->4	
n, an	g->2	n->1	s->4	
n, ar	b->1	
n, at	t->20	
n, av	 ->3	
n, ba	n->1	r->2	
n, be	h->1	
n, bl	.->2	a->3	i->1	
n, bo	r->1	
n, br	i->1	
n, bä	s->2	
n, bå	d->3	
n, bö	r->5	
n, de	 ->2	l->1	m->2	n->13	s->4	t->22	
n, du	 ->1	
n, dv	s->6	
n, dä	r->14	
n, då	 ->3	
n, dö	l->1	
n, ef	t->19	
n, ek	o->1	
n, el	l->5	
n, en	 ->12	l->4	
n, et	a->1	c->1	t->9	
n, ex	a->1	
n, fa	c->1	s->1	
n, fi	c->2	n->1	
n, fl	y->1	
n, fr	a->2	i->1	u->25	ä->3	å->4	
n, få	r->3	t->1	
n, fö	d->1	r->54	
n, ga	n->1	
n, ge	n->5	
n, gj	o->2	
n, gr	u->1	
n, ha	m->1	n->1	r->12	
n, he	l->1	r->56	
n, ho	s->1	
n, hä	n->1	
n, hö	j->1	
n, i 	T->1	b->1	d->4	e->6	f->2	k->1	s->6	
n, ig	å->1	
n, in	f->1	k->2	n->4	o->5	s->1	t->16	
n, ja	 ->1	g->7	
n, ju	 ->1	s->3	
n, ka	m->1	n->5	
n, ko	l->9	m->6	n->1	r->2	s->1	
n, kr	ä->2	
n, ku	n->1	
n, kv	i->1	
n, kä	n->1	r->26	
n, li	k->5	
n, lä	m->2	
n, lå	t->1	
n, ma	n->2	
n, me	d->13	n->42	
n, mi	l->2	n->17	
n, mu	l->1	
n, mä	n->1	
n, må	s->7	
n, na	t->1	
n, nu	 ->1	
n, nä	m->4	r->19	
n, nå	g->5	
n, oc	h->118	
n, of	f->1	
n, om	 ->15	
n, os	v->1	
n, pa	r->4	
n, pr	e->1	i->1	
n, pu	b->1	
n, på	 ->10	m->1	
n, ra	s->1	
n, rä	t->1	
n, rå	d->4	
n, sa	d->1	k->1	m->8	n->1	
n, se	k->1	
n, sk	a->5	o->1	r->1	u->6	
n, sl	u->2	
n, sn	a->2	
n, so	l->1	m->78	
n, st	a->1	r->1	y->1	
n, sä	r->6	
n, så	 ->17	g->1	s->2	v->4	
n, t.	e->3	
n, ta	c->3	r->1	
n, ti	l->12	o->1	
n, tr	o->5	
n, tv	i->1	ä->1	å->1	
n, ty	 ->3	v->1	
n, un	d->2	
n, up	p->2	
n, ut	a->26	i->1	o->1	s->1	t->2	
n, va	d->1	r->9	
n, ve	r->1	
n, vi	 ->6	d->3	l->36	
n, vo	n->1	
n, vä	l->1	r->1	
n, yt	t->1	
n, Îl	e->1	
n, äg	a->1	
n, än	 ->1	d->1	
n, är	 ->18	a->9	
n, äv	e->14	
n, åt	m->1	
n, öp	p->1	
n- oc	h->4	
n-Cla	u->1	
n-Har	r->1	
n-Kee	s->1	
n-SS:	s->1	
n-gru	p->1	
n-råd	e->3	
n. De	r->1	t->6	
n. Dä	r->1	
n. Fo	g->1	
n. Ha	n->1	
n. Hä	r->1	
n. I 	r->1	
n. In	i->1	
n. Ja	g->3	
n. Lå	t->1	
n. Me	n->3	
n. Nä	s->1	
n. Oc	h->3	
n. Rå	d->1	
n. Vi	 ->2	
n." Ä	r->1	
n.(EL	)->1	
n.(IT	)->1	
n.(Li	v->1	
n.(Pa	r->2	
n.) H	e->1	
n.) T	a->1	
n.).H	e->1	
n.)An	d->1	
n.)Be	t->4	
n.)Fr	u->3	
n.)Ge	m->1	
n.)He	r->1	
n.. (	E->6	F->3	
n.. D	e->1	
n..(E	N->1	S->1	
n..(N	L->1	
n..He	r->1	
n.14 	e->1	
n.15 	m->1	
n.All	a->6	m->1	t->4	
n.And	r->1	
n.Ann	a->1	
n.Arb	e->1	
n.Art	i->1	
n.Att	 ->4	
n.Av 	4->1	b->1	d->3	v->1	
n.Avs	a->1	l->1	
n.Bed	r->1	
n.Bet	r->2	
n.Bil	t->1	
n.Bri	s->1	
n.Bry	s->1	
n.Cen	t->1	
n.Cun	h->1	
n.DEB	A->1	
n.De 	d->1	f->1	g->1	h->4	k->5	n->1	o->1	r->1	s->5	u->1	
n.Den	 ->38	n->10	
n.Des	s->10	
n.Det	 ->143	,->1	t->32	
n.Där	 ->2	a->1	f->23	m->2	
n.Då 	d->1	k->1	ä->1	
n.EU 	m->1	ä->1	
n.Eff	e->1	
n.Eft	e->3	
n.Eme	l->1	
n.En 	a->3	d->1	f->1	m->1	s->3	
n.End	a->2	
n.Enl	i->6	
n.Er 	a->1	
n.Eri	k->1	
n.Ett	 ->10	
n.Eur	o->5	
n.Eve	n->1	
n.FEO	 ->1	
n.Fak	t->1	
n.Far	l->1	
n.Fin	n->1	
n.Fle	r->1	
n.For	s->1	
n.Fru	 ->5	
n.Frå	g->4	
n.Fyr	t->1	
n.Föl	j->2	
n.För	 ->29	b->1	e->2	h->1	s->6	u->3	v->1	
n.Gen	o->1	
n.Gol	a->1	
n.Gäl	l->1	
n.Gå 	h->1	
n.Had	e->1	
n.Han	 ->5	
n.Har	 ->2	
n.Hel	a->1	
n.Her	r->56	
n.Hit	 ->1	t->1	
n.Hon	 ->2	
n.Hur	 ->5	
n.Här	 ->6	m->1	
n.I E	u->1	
n.I T	y->1	
n.I a	v->2	
n.I d	a->4	e->10	
n.I e	g->1	n->3	t->1	
n.I f	r->1	
n.I m	i->2	o->1	
n.I r	a->1	å->1	
n.I s	i->1	j->1	t->3	y->1	å->1	
n.I v	e->1	
n.Ill	e->1	
n.Ing	a->1	e->1	
n.Ino	m->1	
n.Inr	ä->1	
n.Ins	a->1	
n.Int	e->2	
n.Ja,	 ->1	
n.Jac	k->1	
n.Jag	 ->133	
n.Jor	d->1	
n.Jus	t->2	
n.Kan	 ->5	
n.Koc	h->1	
n.Kom	m->20	
n.Kon	k->3	
n.Kor	t->1	
n.Kra	v->1	
n.Kul	t->1	
n.Kva	n->1	
n.Led	a->1	
n.Lik	s->1	
n.Liv	s->1	
n.Lån	g->1	
n.Låt	 ->10	
n.Man	 ->6	
n.Mar	k->1	
n.Max	i->1	
n.Med	 ->2	a->1	l->2	
n.Men	 ->35	
n.Min	 ->5	a->1	
n.Mit	t->1	
n.Mot	 ->4	
n.Myn	d->1	
n.Män	n->1	
n.Mär	k->1	
n.Mån	g->1	
n.Möj	l->1	
n.Nat	u->2	
n.Ni 	b->1	h->1	l->1	m->1	s->4	
n.Nie	l->1	
n.Nu 	a->2	f->1	ä->1	
n.Nyl	i->1	
n.När	 ->9	
n.Och	 ->10	
n.Ock	s->1	
n.Om 	S->1	b->1	d->2	g->1	k->2	m->1	n->1	r->1	s->1	t->2	v->5	
n.Ord	e->1	f->3	
n.Ors	a->1	
n.Oz 	h->1	
n.Par	l->4	
n.Per	s->1	
n.Pla	n->1	
n.Pre	c->1	
n.Pro	d->2	
n.På 	d->3	m->1	o->1	s->2	v->2	
n.Ref	o->1	
n.Ren	t->1	
n.Rik	a->1	
n.Rot	h->1	
n.Rät	t->1	
n.Råd	e->4	
n.Sam	h->1	m->2	t->2	
n.San	n->2	
n.Sch	r->1	
n.Sed	a->3	
n.Set	t->1	
n.Sis	t->2	
n.Sit	u->1	
n.Ska	l->1	
n.Sku	l->1	
n.Slu	t->11	
n.Sna	b->1	
n.Soc	i->1	
n.Som	 ->9	l->1	
n.Sta	t->1	
n.Stå	l->1	
n.Stö	d->1	r->1	
n.Sub	v->1	
n.Syf	t->2	
n.Säk	e->1	
n.Sär	s->2	
n.Så 	d->1	l->1	s->1	v->4	
n.Sål	e->1	
n.Tac	k->5	
n.The	a->1	
n.Thy	s->1	
n.Tid	i->1	
n.Til	l->5	
n.Tor	v->2	
n.Tro	t->3	
n.Tvä	r->1	
n.Ty 	s->1	v->1	
n.Tyv	ä->3	
n.Und	a->2	e->6	
n.Uni	o->2	
n.Upp	g->1	
n.Uta	n->1	
n.Uti	f->1	
n.Uts	k->1	
n.Utv	e->1	
n.Vad	 ->13	
n.Val	e->1	
n.Van	l->1	
n.Var	 ->1	j->1	
n.Vet	e->1	
n.Vi 	a->8	b->6	d->1	f->1	g->1	h->11	i->2	j->1	k->9	l->1	m->14	o->1	s->9	t->5	u->1	v->9	ä->5	
n.Vid	 ->4	
n.Vil	k->4	l->1	
n.Vis	s->2	
n.Vit	b->2	
n.Vår	 ->2	a->2	t->1	
n.Wor	l->1	
n.Än 	e->1	
n.Änd	r->1	å->1	
n.Ära	d->2	
n.Äve	n->4	
n.Å E	D->1	
n.Å a	n->1	
n.Å e	n->1	
n.Ögo	n->2	
n.Öve	r->1	
n/Nor	d->2	
n/år)	?->1	
n/år,	 ->1	
n: "d	e->1	
n: At	t->1	
n: De	 ->1	t->1	
n: Er	i->1	
n: Ha	m->1	
n: Ja	g->2	
n: Ko	m->3	
n: Re	v->1	
n: Tå	g->1	
n: Va	d->1	
n: Vi	 ->1	
n: at	t->1	
n: de	f->1	t->1	
n: dä	r->1	
n: en	 ->1	
n: fo	r->1	
n: fö	r->2	
n: i 	F->1	
n: in	s->1	
n: ja	g->1	
n: me	d->2	
n: nä	r->2	
n: va	d->1	r->2	
n: vi	 ->2	
n:För	 ->1	
n; Ja	v->1	
n; av	 ->1	
n; de	n->2	s->2	t->5	
n; dä	r->1	
n; en	l->1	
n; fi	s->1	
n; fö	r->1	
n; in	f->1	
n; me	n->1	
n; oc	h->1	
n; pu	n->1	
n; sa	m->1	
n; sk	o->1	
n; vi	 ->1	
n; än	n->1	
n? 21	 ->1	
n? De	n->1	
n? In	t->1	
n?. (	E->1	
n?Ans	e->1	
n?Den	 ->3	
n?Des	s->1	
n?Det	 ->4	
n?Eft	e->1	
n?Fol	k->1	
n?Fru	 ->2	
n?För	 ->1	s->1	
n?Her	r->3	
n?Hur	 ->1	
n?I d	a->1	
n?Ja,	 ->1	
n?Jag	 ->3	
n?Kan	 ->2	s->1	
n?Kom	m->2	
n?När	 ->1	
n?Om 	i->1	
n?Par	l->1	
n?Sed	a->1	
n?Vad	 ->1	
n?Vem	 ->1	
n?Vet	s->1	
n?Vi 	b->1	f->1	m->1	ä->1	
n?Vil	k->4	
n?Är 	d->2	h->1	i->1	
n?Äve	n->1	
nFråg	a->1	o->2	
nHerr	 ->2	
nI de	n->1	
nJag 	f->2	
nNäst	a->7	
na (K	O->1	
na - 	d->3	e->1	f->4	h->1	i->2	j->1	l->1	m->2	o->1	p->2	r->1	s->2	t->1	u->1	
na 1 	o->2	
na 12	3->1	
na 13	3->1	
na 16	 ->1	
na 33	 ->1	
na 6 	o->1	
na 81	 ->3	.->1	
na 85	 ->3	
na 87	,->1	
na Al	i->1	
na Az	o->1	
na B 	o->1	
na El	l->1	
na Eu	r->1	
na IX	 ->1	
na Li	b->1	
na Mo	u->1	
na Pr	o->1	
na Te	r->1	x->1	
na Tu	r->2	
na ab	s->1	
na ad	m->1	
na af	f->1	
na ak	t->2	
na al	l->2	
na am	b->2	
na an	d->6	g->2	m->1	o->1	s->13	v->7	
na ar	b->4	t->3	
na as	p->1	
na at	t->67	
na av	 ->47	d->1	g->1	l->1	s->6	t->2	
na ba	k->5	r->3	
na be	a->1	d->2	f->4	g->4	h->2	k->2	m->1	s->10	t->7	v->4	
na bi	d->3	l->9	s->1	
na bl	a->1	i->11	
na bo	m->1	r->5	
na br	i->2	o->1	å->1	
na bu	d->5	
na by	g->4	r->1	
na bä	r->1	
na bö	r->7	
na ca	n->1	
na ce	n->1	r->1	
na da	g->3	m->38	t->1	
na de	 ->13	b->25	l->9	m->4	n->6	s->4	t->11	
na di	a->2	f->3	m->1	p->1	r->3	s->1	
na do	k->1	m->2	
na dr	a->6	i->2	
na dy	n->1	
na dä	r->12	
na då	 ->3	
na dö	m->1	r->1	
na ef	f->2	t->4	
na eg	n->15	
na ek	o->5	
na el	l->18	
na em	e->4	
na en	 ->15	d->1	h->3	l->3	v->1	
na er	 ->3	f->1	s->1	
na et	a->2	c->1	t->7	
na eu	r->4	
na ex	e->1	p->2	
na fa	k->2	l->3	m->2	n->1	r->5	s->1	t->1	
na fe	m->1	
na fi	n->7	
na fo	g->1	r->11	
na fr	a->8	i->3	u->3	å->97	
na fu	n->4	
na få	 ->6	n->1	r->13	
na fö	l->4	r->206	
na ga	l->1	m->3	n->1	r->3	v->1	
na ge	 ->7	m->13	n->15	r->2	s->1	
na gi	l->1	v->1	
na gj	o->3	
na gl	ä->1	
na go	d->1	
na gr	a->8	e->1	u->8	ä->1	ö->1	
na gä	l->5	
na gå	 ->2	n->4	r->2	
na gö	r->16	
na ha	 ->1	d->2	m->1	n->6	p->1	r->45	
na he	l->5	m->1	
na hi	n->1	
na hj	ä->2	
na ho	n->3	s->3	
na hu	r->3	v->1	
na hy	s->1	
na hä	n->5	r->5	v->2	
na hå	l->5	v->1	
na hö	g->2	r->3	
na i 	A->2	B->1	C->4	E->38	F->1	I->1	K->2	L->1	M->1	P->2	R->1	T->5	U->1	a->5	b->2	d->43	e->13	f->9	g->5	h->3	i->2	j->1	k->6	m->10	o->3	p->3	r->2	s->7	u->4	v->11	Ö->6	ä->1	
na ib	l->1	
na id	é->2	
na if	r->1	
na ig	e->1	n->1	
na ik	a->1	
na in	 ->2	f->10	h->1	i->2	k->3	l->2	n->5	o->12	r->1	s->9	t->29	v->1	
na jo	b->1	r->1	
na ju	r->2	
na jä	m->1	
na ka	m->23	n->14	t->3	
na kl	a->2	i->1	
na kn	a->1	
na ko	d->2	l->19	m->34	n->19	p->1	r->3	s->3	
na kr	a->1	i->2	ä->2	
na ku	l->1	n->6	
na kv	a->6	o->1	
na kä	l->1	n->6	r->4	
na la	d->1	g->2	n->1	r->1	
na le	d->3	v->3	
na li	b->1	g->2	k->1	t->2	v->1	
na lj	u->1	
na lo	k->2	
na lu	c->1	
na ly	c->1	
na lä	g->2	m->3	n->2	r->1	
na lå	n->1	t->1	
na lö	f->1	p->1	s->9	
na ma	j->1	n->3	r->4	t->1	
na me	d->56	l->19	n->2	s->2	t->1	
na mi	g->1	l->4	n->3	s->1	
na mo	d->2	t->4	
na mu	n->2	
na my	c->6	n->4	
na mä	k->1	n->1	r->1	
na må	l->5	n->1	s->18	
na mö	j->5	t->1	
na na	t->6	
na ne	d->1	g->1	
na no	g->1	r->1	
na nr	 ->2	
na ny	 ->1	a->2	l->1	
na nä	r->8	s->1	
na nå	 ->2	g->5	
na ob	e->1	
na oc	h->163	k->7	
na of	f->1	
na oj	ä->1	
na ol	i->1	j->1	y->2	
na om	 ->64	,->4	f->3	r->1	s->3	
na op	e->1	i->1	
na or	d->5	g->4	o->4	s->1	t->1	
na os	s->9	
na pa	r->9	s->1	
na pe	n->2	r->3	s->1	
na pl	a->3	
na po	l->7	s->1	
na pr	a->2	e->4	i->10	o->18	ö->1	
na pu	m->1	n->9	
na på	 ->37	,->1	:->1	g->1	v->1	
na ra	d->1	m->1	p->6	
na re	d->5	f->14	g->32	l->2	s->23	v->2	
na ri	k->8	
na ro	l->2	
na rä	d->2	k->1	t->8	
na rå	d->4	t->1	
na rö	r->2	s->3	t->2	
na sa	k->1	m->6	t->1	
na se	 ->3	d->2	k->6	n->2	r->4	s->1	t->1	x->1	
na si	d->14	f->4	g->10	n->2	t->12	
na sj	u->2	ä->8	
na sk	a->41	i->3	r->2	u->10	y->1	ö->2	
na sl	a->1	u->7	ä->1	å->1	
na sm	u->1	å->1	
na sn	a->2	e->1	
na so	c->3	l->1	m->60	
na sp	a->1	e->7	o->1	r->1	å->1	
na st	a->9	o->2	r->4	u->3	y->2	ä->6	å->10	ö->10	
na su	m->1	v->1	
na sv	a->3	
na sy	f->1	n->5	s->2	
na sä	g->4	k->2	n->1	r->2	t->3	
na så	 ->4	g->1	s->1	v->1	
na sö	n->1	r->1	
na t.	o->1	
na ta	 ->7	c->3	l->3	n->3	r->3	s->1	
na te	k->1	r->1	x->6	
na ti	d->4	l->56	t->1	
na tj	ä->2	
na to	g->3	r->1	t->2	
na tr	a->1	e->3	i->1	o->1	ä->1	
na tv	i->2	å->4	
na ty	d->1	n->1	p->12	
na tä	n->3	
na ul	t->1	
na un	d->15	i->2	
na up	p->36	
na ur	 ->1	s->1	
na ut	 ->3	a->6	f->3	g->5	l->2	m->2	n->2	s->3	v->14	
na va	c->1	d->1	g->1	l->2	r->18	
na ve	c->4	n->1	r->4	t->2	
na vi	d->12	k->8	l->14	r->1	s->9	t->3	
na vo	n->1	
na vä	g->5	l->1	n->1	r->4	x->1	
na vå	g->1	r->5	
na yr	k->2	
na yt	t->2	
na äm	n->1	
na än	 ->3	d->10	n->3	t->1	
na är	 ->49	.->1	a->1	
na äv	e->2	
na åk	l->1	
na år	e->2	l->1	s->1	
na ås	a->1	i->1	t->1	
na åt	.->1	a->4	e->5	g->10	
na öd	e->2	
na ög	a->1	o->1	
na ök	a->2	n->1	
na ön	s->2	
na öp	p->1	
na ös	t->1	
na öv	e->11	
na!De	t->1	
na!He	r->1	
na!Om	 ->1	
na".D	e->1	
na".K	i->1	
na"in	d->1	
na, B	r->1	
na, S	a->1	
na, a	l->2	r->2	t->5	v->3	
na, b	a->1	e->1	i->1	å->1	
na, d	e->15	v->1	ä->4	å->1	
na, e	f->3	k->1	l->2	n->5	r->1	t->1	
na, f	o->1	r->4	ö->5	
na, g	e->1	
na, h	a->4	e->3	u->2	
na, i	 ->13	n->5	
na, j	a->1	u->2	
na, k	a->2	o->1	
na, l	i->3	ä->1	å->1	
na, m	e->21	i->3	å->1	
na, n	e->1	ä->4	å->3	
na, o	c->31	m->4	r->1	
na, p	å->1	
na, r	e->3	
na, s	a->3	k->1	l->1	o->21	t->2	ä->1	å->12	ö->1	
na, t	a->1	i->5	j->1	o->1	r->3	u->1	
na, u	n->2	t->7	
na, v	a->2	e->1	i->14	o->1	
na, ä	r->1	v->1	
na, ö	v->1	
na-Is	r->1	
na. D	e->1	ä->1	å->1	
na. H	å->1	
na. J	a->1	
na. K	o->1	ä->1	
na. S	o->1	
na. V	a->1	
na. Å	t->1	
na.(T	a->1	
na.)B	e->1	
na.- 	(->2	
na..(	I->1	
na.Al	l->6	
na.Am	s->1	
na.Av	 ->2	
na.Be	s->2	
na.De	 ->5	n->12	s->4	t->40	
na.Do	c->1	
na.Dä	r->6	
na.Ef	t->3	
na.Em	e->1	
na.En	k->1	
na.Et	t->5	
na.Eu	r->3	
na.Fa	c->2	
na.Fr	å->1	
na.Fö	l->1	r->12	
na.Ge	m->1	
na.Gi	v->1	
na.Ha	n->1	
na.He	r->5	
na.Hu	l->1	r->2	
na.Hä	r->2	
na.I 	E->1	b->1	d->3	e->1	l->2	m->1	p->1	t->1	ö->1	
na.Ib	l->1	
na.In	g->1	o->1	t->1	
na.Ja	g->29	
na.Ju	s->2	
na.Ka	f->1	n->1	
na.Ko	m->6	n->2	
na.Li	k->1	v->1	
na.Lå	t->2	
na.Ma	n->1	
na.Me	d->4	n->9	
na.Mi	n->5	
na.Na	t->1	
na.Ni	 ->2	
na.Nu	 ->1	
na.Nä	r->3	
na.Oc	h->1	
na.Om	 ->5	
na.Or	d->1	
na.Pr	e->1	
na.På	 ->4	
na.Re	s->1	
na.Se	d->1	
na.Sk	y->1	
na.Sl	u->3	
na.So	m->3	
na.St	ö->1	
na.Sy	f->1	
na.Så	 ->1	n->1	
na.Ta	c->1	d->1	
na.Ti	l->1	
na.Tr	o->2	
na.Un	d->2	
na.Up	p->1	
na.Ur	 ->1	
na.Ut	a->1	b->1	d->1	n->1	
na.Va	d->3	r->1	
na.Ve	r->1	
na.Vi	 ->29	l->1	s->2	
na.Vä	r->1	s->1	
na.Vå	r->1	
na.Än	 ->1	d->1	
na.Är	 ->1	
na.Äv	e->2	
na.Å 	a->1	
na/Eu	r->1	
na/sa	m->1	
na: F	ö->1	
na: m	a->1	
na: v	i->1	
na; j	a->2	
na; l	o->1	
na; o	c->1	
na; p	u->1	
na?Et	t->1	
na?Ha	r->1	
na?Hu	r->1	
na?I 	F->1	
na?Ja	g->1	
na?Jo	,->1	
na?Ma	n->1	
na?På	 ->1	
na?Sv	a->1	
na?Va	d->2	
na?Vi	 ->1	l->1	
na?Är	 ->1	
naHer	r->1	
nabb 	h->1	o->2	v->1	
nabba	 ->10	r->11	s->3	
nabbt	 ->34	,->3	.->6	
nabbv	a->1	
nabis	e->1	
nacka	t->2	
nackd	e->8	
nad -	 ->1	
nad a	n->1	t->1	v->5	
nad b	e->2	
nad d	å->1	
nad e	f->1	l->1	
nad f	r->2	ö->6	
nad h	a->1	
nad i	 ->6	n->2	
nad j	u->1	
nad k	a->2	o->2	
nad m	e->4	å->2	
nad n	å->1	
nad o	c->2	m->2	
nad r	o->1	ä->1	
nad s	e->1	k->1	o->5	
nad t	i->1	
nad u	r->1	t->2	
nad ö	v->1	
nad, 	"->1	e->1	h->1	i->1	m->2	o->1	s->1	t->1	u->1	ä->1	
nad.D	e->2	
nad.E	u->1	
nad.H	e->2	
nad.J	a->2	
nad.P	a->1	
nad: 	e->1	
nad; 	d->1	
nad?H	e->1	
nad?V	i->1	
nada,	 ->2	
nade 	N->1	a->2	b->6	d->3	e->2	f->3	i->1	j->2	k->17	m->2	n->2	o->2	p->2	r->5	s->4	t->1	u->1	v->2	ä->3	å->2	ö->1	
nade,	 ->1	
nade.	J->1	P->1	T->1	
naden	 ->83	)->3	,->29	.->30	s->19	
nader	 ->57	,->10	.->16	n->79	s->3	
nades	 ->8	.->1	
nads-	 ->1	i->2	n->1	
nads/	i->1	
nadsa	k->1	n->3	r->1	
nadsb	e->4	
nadsd	o->1	
nadse	f->4	k->14	
nadsf	r->4	ö->1	
nadsi	n->3	
nadsk	r->1	
nadsl	i->1	å->1	
nadsm	y->1	ö->1	
nadsn	i->1	
nadso	r->1	
nadsp	r->5	
nadss	t->3	
nadst	i->1	
nadsu	p->1	
nadsv	e->1	i->2	
nafly	k->1	
nafrå	g->1	
nagav	 ->3	
nage 	p->1	
nagel	,->1	
nager	 ->1	
naget	t->1	
nagiv	a->2	i->1	
naiva	 ->1	
naivi	t->1	
nakis	 ->1	!->1	
nakna	,->1	
nakry	.->1	
nal C	o->1	
nal d	e->1	
nal f	r->2	ö->2	
nal i	 ->1	n->2	
nal m	å->1	
nal o	c->1	m->3	r->1	
nal p	l->1	
nal r	a->1	
nal s	o->3	
nal t	i->2	
nal u	t->2	
nal v	a->1	e->1	
nal, 	e->1	n->1	r->1	
nal-s	o->2	
nal. 	J->1	
nal.D	e->1	
nal.F	r->1	
nal.P	e->1	
nal.S	å->1	
nal.V	i->1	
nala 	a->1	e->2	k->1	l->1	m->7	o->14	r->1	s->10	u->9	
nalag	e->1	
nalek	o->4	
nalen	 ->2	
naler	 ->7	,->1	.->2	n->1	
nalfa	b->1	
nalfö	r->3	
nalis	e->21	m->2	t->7	
nalit	e->8	
nalli	b->1	
nalpa	r->1	
nalpo	l->40	
nalpr	o->1	
nalre	s->3	
nalrä	k->1	
nalso	c->1	
nalst	a->3	ö->2	
nalsy	s->1	
nalt 	s->1	
nalut	b->1	
nalve	r->1	
nalys	 ->26	,->4	.->5	?->2	e->21	
namba	l->1	
namik	 ->1	
namis	k->4	
namma	t->4	
namn 	K->1	b->1	k->1	m->1	o->1	s->2	
namn,	 ->2	
namn.	M->1	V->1	
namne	t->2	
namnu	p->4	
nan E	G->1	K->1	u->1	
nan a	m->1	n->1	r->1	
nan b	e->2	l->1	
nan c	e->1	
nan d	a->1	e->9	ä->1	
nan e	k->1	t->1	
nan f	r->2	ö->1	
nan g	r->1	
nan h	a->1	
nan i	 ->5	n->1	
nan j	a->2	u->1	
nan k	o->1	
nan m	a->2	e->4	y->1	å->1	
nan n	i->1	
nan o	c->1	m->1	r->1	
nan p	o->1	
nan r	e->1	i->1	å->1	
nan s	a->3	i->2	k->1	t->2	y->1	
nan t	r->1	
nan v	i->16	
nan å	r->1	s->1	
nan, 	a->1	d->1	f->1	v->1	
nan.L	å->1	
nande	 ->47	,->4	.->6	;->1	?->1	f->1	n->2	t->5	
naner	n->1	
nans 	m->1	o->1	
nansd	e->1	
nanse	r->2	
nansi	e->78	ä->1	
nansl	å->1	
nansm	i->1	
nanst	a->2	
nansv	a->1	
nant 	o->1	
napp 	h->1	
nappa	 ->2	s->9	
nappn	i->1	
nappt	 ->5	
napro	c->2	
nar C	e->1	
nar E	u->1	
nar R	E->1	
nar a	b->1	l->5	t->11	
nar b	e->3	r->1	
nar d	e->24	o->1	r->1	ä->12	ö->1	
nar e	k->1	n->2	r->3	t->3	
nar f	i->1	r->1	ö->4	
nar h	a->1	e->2	j->1	
nar i	 ->15	g->1	n->3	
nar j	a->15	u->3	
nar k	a->2	l->1	o->12	r->1	
nar l	ä->1	
nar m	a->2	e->15	i->2	o->1	y->1	
nar n	i->1	ä->2	å->1	
nar o	c->8	l->1	m->3	r->5	s->5	
nar p	a->2	
nar r	ä->1	å->2	ö->1	
nar s	i->6	k->7	t->2	ä->1	å->1	
nar t	i->7	
nar u	p->1	t->4	
nar v	a->3	e->1	i->12	å->1	
nar Ö	V->1	
nar ä	n->1	r->1	
nar å	t->2	
nar ö	n->1	
nar, 	e->1	m->1	o->1	p->1	s->1	t->1	v->1	
nar..	 ->1	
nar.D	e->4	
nar.H	e->2	
nar.M	a->1	
nar.O	m->1	
nar.S	t->1	å->1	
nar.U	t->1	
nar.V	i->1	
nar: 	o->1	
narar	e->24	
naras	t->13	
narbe	t->1	
nard 	K->1	
nare 	b->1	d->3	e->2	f->4	g->1	h->2	i->4	k->2	o->1	p->1	r->1	s->3	t->5	ä->1	å->4	
nare,	 ->5	
nare.	D->2	I->1	M->1	S->1	
narel	ä->1	
naren	 ->3	,->1	s->1	
narep	r->1	
narie	r->1	
nario	 ->1	r->1	t->2	
nariu	m->1	
narko	m->1	t->6	
narli	k->1	
narna	 ->9	,->1	.->5	s->2	
nars 	b->1	f->1	h->2	i->3	k->5	m->1	s->3	t->1	ä->1	
nars,	 ->1	
narsa	m->4	
nart 	-->1	a->2	d->1	h->1	k->3	m->2	s->15	v->1	
nart.	J->1	
naråd	a->1	
nas E	u->7	
nas S	j->2	
nas a	g->1	l->1	n->16	r->5	t->3	v->10	x->1	
nas b	e->3	l->1	ä->1	
nas c	e->1	
nas d	e->3	i->1	u->1	ä->4	
nas e	f->1	g->2	k->2	l->1	n->9	t->4	
nas f	a->1	l->1	r->3	u->1	ö->24	
nas g	a->1	e->3	r->1	
nas h	a->1	ä->3	å->1	
nas i	 ->6	d->1	n->16	r->1	
nas j	u->1	ä->1	
nas k	a->4	l->1	o->5	r->3	u->1	v->3	ä->1	ö->1	
nas l	a->4	e->3	i->1	ä->1	
nas m	a->2	e->8	i->1	ö->4	
nas n	a->5	i->1	u->1	ä->1	å->5	
nas o	c->19	f->3	i->2	m->3	r->3	
nas p	a->2	e->2	l->2	o->2	r->4	å->3	
nas r	e->5	o->2	ä->7	ö->1	
nas s	a->5	i->5	k->3	l->1	o->4	p->3	t->5	u->4	v->1	ä->2	å->1	
nas t	i->10	j->1	r->2	u->1	v->1	y->1	
nas u	n->1	p->1	t->4	
nas v	a->3	e->1	i->1	ä->4	
nas y	r->1	
nas ä	n->1	r->1	
nas å	l->2	r->1	t->1	
nas ö	p->1	v->1	
nas!E	u->1	
nas, 	a->1	b->1	e->1	h->1	o->3	s->2	u->1	
nas. 	D->1	
nas.D	e->3	
nas.E	n->1	
nas.J	a->1	
nas.K	o->1	
nas.M	e->1	
nas.V	i->1	
nas.Å	t->1	
nast 	a->1	i->2	k->2	l->1	m->1	o->1	u->2	v->2	å->1	
nast?	V->1	
naste	 ->63	
nastå	e->2	
nat -	 ->1	
nat 3	9->1	
nat E	u->1	
nat I	t->1	
nat K	i->1	
nat a	l->1	n->1	v->1	
nat b	a->1	e->4	i->1	l->1	ö->1	
nat d	e->3	i->2	r->1	ö->1	
nat e	f->1	n->2	
nat f	a->7	o->1	r->1	å->1	ö->6	
nat g	e->2	ö->3	
nat h	a->1	å->1	
nat i	 ->6	c->2	f->1	n->5	
nat j	a->1	
nat k	o->9	
nat l	a->2	e->1	ä->1	
nat m	e->2	i->1	y->1	å->1	
nat o	c->6	m->1	r->1	
nat p	r->2	å->4	
nat r	å->1	ö->2	
nat s	a->1	i->2	j->1	k->2	t->1	y->1	ä->5	å->1	ö->1	
nat t	a->3	i->10	
nat u	n->2	p->2	t->3	
nat v	a->1	i->4	ä->1	
nat ä	m->1	n->12	
nat å	r->3	
nat ö	k->1	
nat, 	e->1	h->1	v->1	ä->1	
nat. 	H->1	
nat.D	e->1	
nat.G	e->1	
nat.J	a->1	
nat.K	o->1	
nat.Ä	n->1	
naten	,->1	
natio	n->271	
nativ	 ->7	.->1	;->1	a->2	t->1	
nats 	e->1	f->2	i->2	p->1	t->3	ä->1	å->1	
nats,	 ->2	
nats.	D->1	E->1	
natt 	o->1	
natte	n->2	
natur	 ->3	,->2	-->1	.->3	a->1	e->8	k->13	l->87	n->1	o->1	v->1	
nauer	 ->1	
navgi	f->2	
navis	k->1	
navta	l->3	
nazis	m->8	t->8	
nbana	 ->1	
nbar 	s->1	
nbar.	D->1	F->1	
nbara	.->1	
nbarl	i->12	
nbarn	 ->1	
nbart	 ->49	,->1	.->1	
nbegr	i->12	
nbeha	n->1	
nber 	m->1	v->1	
nberg	 ->3	
nbest	ä->1	
nbetä	n->5	
nbila	r->8	
nbind	a->1	
nbjud	a->2	e->1	n->3	
nbjöd	 ->1	
nblan	d->16	
nblic	k->16	
nboen	d->1	
nbok 	o->1	
nboke	n->1	
nbrot	t->1	
nbryt	a->1	
nbuds	f->2	i->2	
nbul 	f->1	
nbund	e->1	
nburg	 ->1	,->1	h->1	
nbygg	d->1	
nc då	 ->1	
nc, d	v->1	
nca, 	o->1	
ncas 	s->1	
nce, 	D->1	
nce..	.->1	
ncent	r->31	
ncept	 ->2	.->2	e->3	
ncer!	D->1	
ncer,	 ->1	
ncera	t->1	
ncerb	ö->1	
ncern	e->2	
nchen	.->1	
nchez	 ->1	
nchti	d->1	
ncide	n->1	
ncil 	-->1	
ncip 	a->3	e->3	f->1	i->7	o->4	r->1	s->5	ä->4	
ncip,	 ->3	
ncip.	J->1	S->1	V->2	
ncipe	n->102	r->48	s->1	
ncipi	e->8	
ncips	k->1	
ncis 	W->1	a->1	
ncist	 ->1	
ncita	m->8	
nckhe	e->14	
nd (e	f->1	
nd (k	o->1	
nd (r	å->1	
nd - 	E->1	d->1	m->1	Ö->1	
nd 80	 ->1	
nd EU	-->1	
nd LT	C->1	
nd La	n->3	
nd Sv	e->1	
nd Ti	b->1	
nd ac	q->1	
nd al	l->4	
nd an	d->2	n->18	s->2	
nd at	t->11	
nd av	 ->80	
nd be	d->1	h->1	r->2	v->3	
nd bi	b->1	
nd by	g->1	
nd bå	d->1	
nd ci	r->1	
nd de	 ->7	f->1	m->2	n->5	s->1	t->1	
nd dä	r->5	
nd ef	f->1	
nd el	l->3	
nd en	 ->9	
nd er	 ->1	t->1	
nd fi	n->1	
nd fo	r->1	
nd fr	å->6	
nd fy	r->1	
nd fö	l->1	r->25	
nd ge	m->1	n->1	r->1	
nd go	d->1	
nd gr	u->1	
nd ha	n->4	r->9	
nd i 	E->1	a->1	d->2	e->4	f->2	k->1	r->2	s->4	t->1	u->1	v->1	
nd in	o->1	t->4	
nd iv	ä->1	
nd ju	s->1	
nd ka	n->1	
nd ko	m->2	n->2	
nd kv	i->3	
nd kä	n->1	
nd la	d->1	
nd lä	g->1	n->1	
nd me	d->50	l->3	r->1	t->1	
nd mi	n->3	
nd my	c->1	
nd må	n->1	s->2	
nd ny	l->1	
nd nä	m->1	r->4	
nd nö	d->1	
nd oc	h->25	k->1	
nd om	 ->14	f->1	
nd os	s->6	
nd pa	l->1	
nd på	 ->4	f->1	
nd re	g->1	n->1	
nd se	 ->1	d->5	
nd si	g->1	
nd sj	ä->1	
nd sk	a->1	u->3	
nd sm	ä->1	
nd so	c->1	m->24	
nd st	a->2	r->2	ö->1	
nd sy	m->1	
nd sä	g->4	
nd så	 ->2	
nd t.	o->1	
nd ta	l->1	
nd ti	l->11	
nd tv	å->1	
nd un	d->4	
nd up	p->1	
nd ut	a->2	v->1	
nd va	r->4	
nd ve	r->2	
nd vi	 ->1	l->1	s->2	
nd vä	r->1	
nd vå	r->1	
nd än	d->1	
nd är	 ->17	
nd åt	 ->1	
nd öv	e->1	
nd! L	i->1	
nd! N	i->1	
nd), 	o->1	
nd, 5	6->1	
nd, D	a->1	
nd, E	C->1	
nd, F	i->1	
nd, I	t->2	
nd, N	o->1	
nd, S	p->2	
nd, b	ö->1	
nd, d	v->1	ä->2	å->1	
nd, f	ö->3	
nd, h	a->1	y->1	
nd, k	a->1	r->1	
nd, l	ä->1	
nd, m	e->4	i->1	
nd, n	å->1	
nd, o	c->7	
nd, p	å->1	
nd, r	e->1	ä->1	
nd, s	k->1	o->3	ä->1	å->1	
nd, t	o->1	
nd, u	n->2	
nd, v	i->2	
nd- (	P->1	
nd. V	i->1	
nd.An	d->1	
nd.At	t->1	
nd.De	n->2	t->6	
nd.Di	r->2	
nd.Em	e->1	
nd.Fr	å->1	
nd.Ge	n->1	
nd.He	r->1	
nd.I 	k->1	s->1	
nd.In	f->1	i->1	n->1	
nd.Ir	l->1	
nd.Ja	g->7	
nd.Ko	m->1	n->1	
nd.Lå	t->1	
nd.Me	n->1	
nd.Mi	t->1	
nd.Ni	 ->1	
nd.Nu	 ->1	
nd.Nä	r->1	
nd.Om	 ->2	
nd.På	 ->1	
nd.So	m->1	
nd.Up	p->1	
nd.Va	r->1	
nd.Vi	 ->2	
nd.Å 	a->1	
nd? H	a->1	
nd?. 	(->1	
nd?Fö	r->1	
nd?Ja	g->1	
nda -	 ->1	
nda 1	2->1	
nda 2	0->1	
nda E	U->1	r->1	
nda a	l->3	n->2	r->1	t->4	v->8	
nda b	a->2	e->1	
nda c	h->1	
nda d	e->19	o->1	r->1	
nda e	l->2	n->6	r->1	u->1	
nda f	i->1	r->3	ö->14	
nda g	i->1	r->1	
nda h	a->2	y->1	
nda i	 ->5	g->2	n->6	
nda j	a->2	o->2	
nda k	o->1	
nda l	a->2	o->1	u->1	
nda m	a->2	e->4	o->1	y->1	å->1	
nda n	e->1	i->1	ö->1	
nda o	c->1	m->3	r->2	s->1	
nda p	a->2	e->2	o->1	r->4	u->1	å->2	
nda r	e->3	i->1	y->1	ö->1	
nda s	a->1	e->4	i->9	k->2	o->9	t->5	u->1	ä->5	
nda t	e->1	i->4	
nda u	n->1	p->1	t->1	
nda v	e->1	i->2	ä->1	
nda ä	n->2	r->2	
nda ö	a->1	r->1	
nda, 	f->1	k->1	s->3	v->2	
nda.B	e->1	
nda.D	e->2	å->1	
nda.F	r->1	ö->1	
nda.H	e->1	
nda.I	 ->1	
nda.K	ä->1	
nda.M	i->1	
nda.N	i->1	ä->1	
nda.R	u->1	
nda.V	i->2	
nda?D	e->1	
ndabo	c->2	
ndad 	a->1	i->1	p->3	r->1	
ndade	 ->8	,->1	.->1	s->1	
ndag 	o->1	
ndage	n->2	
ndags	 ->1	.->1	
ndahå	l->43	
ndair	e->1	
ndal!	H->1	
ndal,	 ->1	
ndala	n->1	
ndale	r->5	
ndalö	s->1	
ndama	f->1	
ndame	n->1	
ndamå	l->13	
ndan 	b->1	e->1	f->1	i->5	k->1	m->2	o->1	p->1	v->1	
ndan,	 ->2	
ndan.	D->1	
ndanb	e->2	
ndand	e->17	r->1	
ndanf	l->1	
ndanh	å->1	
ndanm	a->1	
ndano	r->1	
ndanr	ö->6	
ndant	a->39	
ndar 	e->1	h->1	i->2	m->2	n->1	o->1	s->1	
ndard	 ->6	,->2	.->1	;->1	e->5	i->9	
ndare	 ->7	,->1	n->2	
ndarn	a->4	
ndars	k->1	
ndas 	f->2	i->2	m->1	o->1	p->10	s->1	t->3	
ndas,	 ->1	
ndas.	A->1	H->1	I->1	M->1	V->1	Å->1	
ndast	 ->82	
ndat 	a->3	f->1	h->1	m->1	p->4	s->2	
ndat,	 ->4	
ndate	n->1	t->4	
ndati	o->33	
ndatp	e->9	
ndbar	 ->1	a->3	t->5	
ndbet	ä->1	
ndbul	t->1	
nde "	a->1	k->1	s->1	
nde (	A->29	m->1	
nde -	 ->15	
nde 1	2->1	
nde A	h->1	l->2	
nde B	 ->1	
nde D	u->1	
nde E	U->1	u->3	
nde G	a->3	r->2	
nde I	m->1	
nde J	a->1	
nde K	a->2	o->2	
nde L	a->1	o->1	
nde M	a->3	e->1	
nde N	a->1	
nde O	L->1	
nde P	r->14	
nde R	a->1	o->2	
nde S	a->1	c->2	e->1	
nde a	b->1	d->3	g->1	i->1	l->5	n->16	p->2	r->3	s->2	t->29	v->150	
nde b	a->7	e->38	i->7	l->2	o->1	r->9	y->2	å->1	
nde d	a->4	e->50	i->8	o->2	r->1	ä->3	å->2	
nde e	f->2	j->1	k->5	l->5	n->12	p->1	r->1	t->6	u->5	x->16	
nde f	a->8	e->2	i->12	l->1	o->6	r->46	u->1	ä->1	å->5	ö->98	
nde g	a->2	e->8	i->1	o->1	r->5	ö->2	
nde h	a->20	e->3	i->2	j->1	o->4	u->2	ä->4	å->1	ö->2	
nde i	 ->54	d->1	g->1	n->49	t->1	
nde j	a->2	o->1	ä->1	
nde k	a->9	l->1	n->1	o->35	r->4	u->1	v->5	ä->2	
nde l	a->7	e->2	i->5	o->3	y->1	ä->3	
nde m	a->13	e->28	i->8	o->4	y->7	ä->1	å->12	ö->1	
nde n	e->2	u->1	y->3	ä->5	å->3	
nde o	c->81	f->2	l->3	m->45	n->2	p->1	r->13	s->1	t->1	
nde p	a->12	e->10	o->13	r->28	u->7	å->33	
nde r	a->4	e->41	i->7	o->7	u->2	ä->29	å->3	ö->2	
nde s	a->15	e->5	i->10	k->10	l->1	o->44	p->2	t->21	v->1	y->13	ä->14	å->1	
nde t	a->15	e->4	i->30	j->6	r->6	v->4	
nde u	n->7	p->7	r->1	t->27	
nde v	a->9	e->8	i->12	o->2	r->1	ä->8	å->1	
nde ä	n->7	r->25	v->1	
nde å	 ->1	r->14	s->1	t->24	
nde ö	a->1	k->1	n->1	p->1	v->12	
nde! 	J->5	N->1	
nde!A	l->1	
nde!J	a->1	
nde!N	i->1	
nde",	 ->1	
nde(A	5->1	
nde, 	,->1	D->1	F->1	G->1	L->1	a->4	b->4	d->6	e->4	f->8	h->5	i->10	j->1	k->6	l->1	m->8	n->4	o->15	p->4	s->14	t->5	u->2	v->9	ä->2	
nde. 	D->2	M->1	
nde.-	 ->1	
nde..	 ->1	
nde.A	v->2	
nde.D	e->25	ä->3	
nde.E	f->2	m->1	n->3	
nde.F	P->1	r->1	ö->2	
nde.G	r->1	
nde.H	a->1	e->5	o->1	u->4	
nde.I	 ->2	n->2	
nde.J	a->26	
nde.K	a->2	o->2	
nde.L	i->1	y->1	å->1	
nde.M	a->4	e->7	i->2	
nde.N	i->1	u->1	ä->1	
nde.O	c->1	m->3	
nde.P	a->1	o->1	
nde.S	a->1	c->1	e->1	o->2	t->1	å->1	
nde.T	a->2	i->1	r->1	v->1	
nde.U	n->2	
nde.V	a->2	i->8	
nde.Å	t->1	
nde: 	"->2	A->3	D->2	F->3	G->3	H->1	I->1	J->2	K->3	M->1	N->2	P->1	S->2	T->1	U->1	V->3	b->1	f->1	i->1	t->1	Å->2	
nde; 	d->2	h->1	p->1	
nde?F	ö->1	
nde?H	e->2	
nde?V	i->1	
ndebe	s->1	
ndebu	d->9	
ndebä	n->1	
ndefr	i->1	
ndefö	r->12	
ndehö	j->1	
ndeko	d->8	l->1	
ndekr	i->1	
ndel 	a->3	k->1	o->3	p->2	s->1	t->1	ä->1	
ndel,	 ->4	
ndel.	D->1	E->1	J->1	
ndela	d->1	n->3	r->4	s->1	
ndele	n->1	
ndeln	 ->2	i->1	
ndels	e->43	f->2	h->1	l->1	m->2	o->5	p->4	s->1	v->1	
ndeme	n->5	
ndemi	s->1	
nden 	(->1	,->1	-->2	B->1	G->2	K->5	L->1	P->3	R->1	T->1	a->14	b->7	d->4	e->7	f->36	g->4	h->12	i->12	j->1	k->7	m->11	n->1	o->35	p->5	r->1	s->25	t->13	u->1	v->5	ä->10	å->1	ö->1	
nden"	 ->1	
nden,	 ->43	
nden.	 ->1	A->1	D->10	F->4	H->2	I->2	J->6	K->2	L->1	M->1	P->1	S->1	T->2	V->4	
nden:	 ->2	F->1	
nden;	 ->1	
nden?	N->1	
ndenN	ä->1	
ndena	 ->30	,->3	.->5	;->1	?->1	
ndenb	u->2	
ndens	 ->15	,->2	e->7	
nder 	-->1	1->8	2->2	4->1	E->3	F->2	N->2	a->12	b->15	d->133	e->20	f->38	g->7	h->17	i->22	j->2	k->11	l->2	m->33	n->13	o->25	p->13	r->9	s->63	t->16	u->10	v->19	ä->5	å->11	ö->1	
nder"	 ->1	
nder,	 ->27	
nder.	 ->2	A->1	B->1	D->6	E->2	F->1	H->1	I->4	J->7	K->2	M->2	N->1	R->1	T->1	V->3	Ä->2	
nder?	H->1	Ä->1	
ndera	 ->11	,->1	d->1	n->1	r->19	s->2	t->1	
nderb	a->1	l->2	
nderd	e->4	
ndere	g->3	
nderg	r->4	
nderh	u->2	å->3	
nderk	a->4	u->1	
nderl	a->7	e->2	i->5	ä->19	å->3	
nderm	e->1	i->1	å->1	
ndern	a->132	
ndero	r->4	
nderr	e->2	ä->1	
nders	 ->6	k->3	t->38	å->1	ö->48	
ndert	e->17	
nderu	t->3	
nderv	i->1	
nderä	t->3	
nderö	s->1	
ndes 	-->1	a->3	e->1	f->2	i->2	j->1	p->1	s->1	
ndes,	 ->1	
ndesk	a->113	i->1	y->1	
ndest	a->1	
ndet 	"->1	-->1	E->1	G->1	M->1	P->3	S->1	a->199	b->6	d->4	e->3	f->27	g->4	h->10	i->18	k->5	l->2	m->15	n->2	o->26	p->3	r->3	s->19	t->5	u->5	v->6	ä->9	å->2	ö->1	
ndet)	 ->1	
ndet,	 ->22	
ndet.	-->1	.->1	A->2	B->1	D->10	H->2	I->1	J->5	M->2	P->1	S->3	U->1	V->3	Ö->1	
ndet;	 ->1	
ndet?	V->1	
ndeta	k->1	
ndets	 ->15	
ndeva	l->6	
ndevi	s->2	
ndful	l->1	
ndfäl	l->4	
ndför	d->1	t->1	u->2	
ndgän	g->2	
ndgår	d->2	
ndgåt	t->1	
ndi r	e->1	
ndi s	o->1	
ndi: 	f->1	
ndica	p->1	
ndida	t->14	
ndie,	 ->1	
ndien	 ->4	s->1	
ndier	,->1	
ndig 	d->4	e->1	f->4	g->1	i->2	j->1	m->1	o->4	p->1	r->2	s->1	t->3	
ndig,	 ->2	
ndig.	D->1	M->1	U->1	
ndiga	 ->32	,->2	.->3	r->2	
ndigh	e->210	
ndigt	 ->100	,->8	.->4	?->1	v->7	
ndika	p->4	t->6	
ndina	v->1	
ndire	k->7	
ndis 	B->1	
ndisk	a->1	
ndit 	s->3	
nditi	o->1	
ndivi	d->14	
ndkur	s->1	
ndla 	d->7	f->1	g->1	i->2	m->1	o->7	s->1	u->1	
ndla.	D->1	V->1	
ndlad	 ->1	e->9	
ndlar	 ->115	e->2	n->1	
ndlas	 ->12	,->1	.->1	
ndlat	 ->6	s->1	
ndlig	 ->6	a->7	h->2	t->7	
ndlin	g->186	
ndläg	g->75	
ndlös	a->1	
ndmed	e->3	
ndmän	 ->1	
ndna 	k->1	r->1	s->1	t->1	
ndnin	g->74	
ndo.F	ö->1	
ndom 	o->1	r->1	
ndoml	i->2	
ndomr	å->14	
ndoms	 ->1	
ndon 	b->1	
ndon,	 ->2	
ndon.	O->1	
ndors	a->1	
ndpel	a->1	
ndpri	n->1	
ndpun	k->103	
ndra 	-->1	E->2	R->1	a->20	b->17	d->18	e->12	f->31	g->14	h->12	i->18	k->12	l->16	m->26	n->6	o->26	p->25	r->17	s->46	t->8	u->3	v->13	y->2	ä->7	å->3	ö->1	
ndra,	 ->22	
ndra.	D->2	J->1	N->2	U->1	V->1	
ndra:	 ->4	
ndra;	 ->2	
ndrab	e->5	
ndrad	 ->1	e->20	
ndrag	 ->3	
ndrah	a->1	
ndrak	a->1	
ndran	 ->2	d->2	
ndrar	 ->23	,->1	e->6	n->3	
ndras	 ->17	,->2	.->4	
ndrat	 ->8	a->5	s->8	u->3	
ndre 	a->2	b->3	d->1	e->2	f->6	g->1	h->1	i->1	k->4	l->3	m->1	o->3	p->3	r->1	s->4	t->2	u->5	v->1	ä->8	
ndre.	D->1	
ndre?	V->1	
ndren	 ->3	
ndres	a->2	
ndrin	g->314	
ndrom	e->1	
ndrän	k->2	
nds a	l->1	
nds b	e->3	
nds d	e->2	
nds e	n->1	
nds f	e->1	ö->4	
nds g	r->1	
nds i	 ->1	n->3	
nds l	a->1	
nds m	e->2	y->1	
nds n	y->1	
nds o	b->1	m->1	
nds p	a->1	å->6	
nds r	e->1	
nds v	i->1	
nds å	t->1	
nds, 	s->1	
ndsam	t->4	
ndsan	m->1	
ndsat	s->1	
ndsav	g->3	
ndsbe	h->1	
ndsby	g->43	
ndsde	l->12	
ndsju	k->1	
ndsk 	a->1	k->3	t->1	
ndsk-	b->1	
ndska	 ->18	,->2	n->1	p->1	s->8	
ndsko	g->1	n->4	
ndskt	 ->1	
ndslä	n->2	
ndsme	d->6	
ndsmä	n->3	
ndspl	a->3	
ndspo	l->2	
ndspr	o->3	
ndsre	g->1	p->4	
ndsrö	r->1	
ndssy	s->1	
ndsta	g->2	
ndste	n->1	
ndsvä	g->1	
ndsän	d->1	
ndt f	r->1	
ndt h	a->1	
ndt o	c->1	
ndt s	a->1	
ndt t	a->1	
ndt u	t->1	
ndt, 	f->1	
ndtes	,->1	
ndupp	b->1	r->2	
ndust	r->114	
nduty	p->1	
ndvag	n->1	
ndval	 ->20	a->3	e->1	
ndvat	t->1	
ndvik	a->31	e->3	i->1	l->4	
ndvin	n->2	
ndzio	-->4	
ndärr	ä->1	
ndå A	s->1	
ndå a	n->2	t->6	
ndå b	a->1	e->1	l->2	o->1	
ndå d	å->1	
ndå e	n->5	
ndå f	i->1	r->1	å->1	ö->2	
ndå g	e->1	ö->1	
ndå h	a->2	e->1	
ndå i	 ->1	n->3	
ndå k	a->2	o->1	v->1	
ndå l	a->1	
ndå o	c->1	e->1	
ndå s	k->2	o->1	å->1	
ndå t	a->2	i->1	v->1	
ndå u	n->2	p->2	
ndå v	i->1	
ndå ä	r->2	
ndå, 	n->1	
ndå..	.->1	
ndée,	 ->1	
ndövt	 ->1	
ne Fo	r->1	
ne an	d->1	s->1	
ne at	t->3	
ne av	 ->1	
ne bl	a->1	
ne de	l->1	
ne di	e->1	
ne ek	o->1	
ne fo	r->1	
ne fr	å->2	
ne få	r->1	
ne fö	r->4	
ne gä	l->1	
ne ha	n->1	r->4	
ne hj	ä->1	
ne hö	g->1	
ne i 	F->1	f->2	s->1	
ne in	d->1	l->1	o->1	
ne ja	g->1	
ne je	t->1	
ne ka	n->1	
ne ko	m->1	
ne lo	k->1	
ne nä	r->4	
ne nå	g->1	
ne nö	j->1	
ne oc	h->6	
ne om	 ->2	
ne på	 ->1	,->1	
ne qu	a->2	
ne ry	k->1	
ne so	m->5	
ne så	 ->1	
ne ti	l->2	
ne to	l->1	
ne va	r->1	
ne vi	l->1	
ne är	 ->2	
ne åk	l->1	
ne! N	i->1	
ne, E	r->1	
ne, R	a->1	
ne, d	v->1	ä->1	
ne, g	ö->1	
ne, k	ä->1	
ne, n	ä->1	
ne, t	y->1	
ne, ä	r->1	
ne- o	c->1	
ne-Al	p->1	
ne-Ar	d->1	
ne-Ma	n->1	
ne-st	o->1	
ne.De	t->3	
ne.Ja	g->1	
ne: N	a->1	
nearb	e->1	
nearv	e->1	
nebar	 ->1	
neboe	n->1	
nebär	 ->90	,->1	.->2	a->15	
nebör	d->7	
ned a	v->2	
ned d	e->1	
ned e	n->2	t->1	
ned f	ö->1	
ned i	 ->5	
ned m	i->2	y->1	
ned n	å->1	
ned o	c->1	
ned p	å->2	
ned t	i->1	
ned v	å->1	
ned.E	f->1	
ned.J	a->1	
neder	l->9	
nedgå	n->2	
nedla	g->1	
nedlä	g->4	
nedmo	n->3	
nedom	e->1	
nedra	n->2	
nedru	s->1	
nedsk	r->1	ä->3	
nedst	ä->3	
nedvr	i->12	
nedvä	r->1	
neexe	m->1	
nefat	t->6	
neffe	k->3	
nefit	-->5	
negat	i->26	
nehar	 ->2	
nehav	a->1	
nehål	l->78	
nehöl	l->4	
nej l	å->1	
nej t	i->1	
nej, 	b->1	s->1	
nej.(	A->1	
neka 	a->1	d->2	f->1	
neka,	 ->1	
neka.	M->1	
nekad	 ->1	
nekan	d->2	
nekar	 ->2	
nekas	 ->2	
nelag	 ->1	
neler	n->1	
nelig	h->1	t->1	
nell 	b->1	d->3	e->2	f->5	k->5	m->1	n->7	o->3	p->5	r->8	s->4	t->1	u->1	v->1	å->1	ö->2	
nell,	 ->3	
nell.	D->1	V->1	
nella	 ->197	,->1	
nellt	 ->26	,->2	
neln,	 ->1	
neln.	D->1	
nelse	 ->1	
neltr	a->1	
nelux	,->1	
neman	g->4	
nen "	L->1	
nen (	B->2	I->1	i->1	o->1	s->1	
nen -	 ->7	
nen C	h->1	
nen E	n->2	
nen I	X->1	
nen J	a->1	
nen P	r->1	
nen a	l->3	m->1	n->12	r->1	t->63	v->33	
nen b	a->2	e->19	i->3	l->1	o->4	y->1	ö->6	
nen d	e->3	r->1	ä->5	
nen e	f->1	g->2	l->5	n->7	t->2	
nen f	a->2	e->1	i->2	o->2	r->12	u->3	ä->2	å->6	ö->59	
nen g	e->6	i->1	j->4	l->2	o->3	ä->1	å->1	ö->4	
nen h	a->55	e->1	i->1	o->4	u->1	å->2	
nen i	 ->62	n->26	
nen j	u->1	
nen k	a->25	l->1	o->35	r->3	u->2	ä->2	
nen l	a->3	i->1	ä->5	
nen m	e->12	o->1	y->1	å->21	ö->1	
nen n	o->2	u->7	y->1	ä->3	å->1	
nen o	c->87	f->3	m->29	
nen p	a->1	l->3	r->2	å->22	
nen r	e->12	i->1	ä->4	å->1	
nen s	a->1	e->3	i->4	j->6	k->34	n->2	o->29	t->12	ä->2	å->6	
nen t	a->1	i->16	r->3	v->1	y->2	ä->1	
nen u	n->10	p->4	t->7	
nen v	a->3	e->4	i->16	ä->1	
nen ä	n->7	r->35	v->1	
nen å	l->1	t->2	
nen ö	k->2	v->2	
nen!N	ä->1	
nen".	D->1	
nen)N	ä->1	
nen, 	I->1	a->4	b->2	d->5	e->6	f->11	h->2	i->7	k->1	l->2	m->10	n->2	o->11	p->4	r->2	s->21	t->3	u->4	v->9	ä->5	å->1	
nen. 	D->3	H->1	
nen.(	E->1	
nen.)	A->1	B->4	G->1	
nen..	 ->5	(->1	H->1	
nen.1	5->1	
nen.A	l->2	
nen.B	e->1	i->1	
nen.D	e->28	ä->8	å->1	
nen.E	f->1	n->2	t->3	u->1	
nen.F	r->1	ö->5	
nen.G	e->1	
nen.H	e->10	i->1	
nen.I	 ->4	
nen.J	a->16	
nen.K	o->2	
nen.L	i->1	å->1	
nen.M	a->1	e->2	i->2	y->1	
nen.N	i->1	u->1	y->1	ä->3	
nen.O	c->2	m->2	
nen.P	a->2	e->1	r->1	å->3	
nen.R	å->2	
nen.S	e->1	l->1	å->1	
nen.T	r->1	
nen.U	n->1	t->1	
nen.V	a->2	i->14	
nen.Ä	v->2	
nen: 	K->1	
nen; 	i->1	m->1	o->1	
nen?H	e->1	
nen?K	a->1	
nen?V	i->1	
nen?Ä	r->1	
nenJa	g->2	
nena 	k->1	o->1	
nener	g->8	
nens 	2->1	B->1	E->2	X->1	a->22	b->13	c->1	d->8	e->20	f->43	g->8	h->9	i->26	k->15	l->10	m->20	n->6	o->14	p->15	r->40	s->44	t->17	u->25	v->15	y->4	å->4	ö->5	
nens,	 ->1	
nent 	i->1	k->2	o->3	u->1	
nent,	 ->1	
nent.	E->1	
nenta	 ->2	l->2	
nente	n->1	r->3	
nenti	e->1	
neona	z->1	
neonl	a->1	
nepot	i->5	
ner (	C->2	a->1	
ner -	 ->6	
ner E	M->1	
ner I	-->1	I->3	
ner J	o->1	
ner K	i->1	v->1	
ner [	S->1	
ner a	l->1	n->1	r->4	t->10	v->3	
ner b	a->1	e->2	i->7	r->1	ä->1	
ner d	e->12	o->5	ä->4	å->2	ö->1	
ner e	c->1	f->2	l->4	n->4	u->17	
ner f	a->3	l->1	o->5	r->5	å->1	ö->15	
ner g	e->5	o->1	å->1	ö->1	
ner h	a->6	i->1	ä->2	å->1	
ner i	 ->23	g->1	n->21	r->1	
ner j	a->4	u->1	
ner k	a->4	o->4	u->2	
ner l	i->1	ä->1	
ner m	a->4	e->27	i->6	o->3	ä->5	å->1	
ner n	i->2	u->1	ä->2	
ner o	c->47	m->7	s->13	
ner p	r->1	å->6	
ner r	e->1	ä->1	
ner s	a->2	i->19	j->1	k->3	l->1	n->1	o->45	p->1	t->4	å->3	
ner t	a->1	i->30	o->2	r->1	
ner u	n->3	t->2	
ner v	a->1	i->9	ä->3	
ner ä	n->3	r->4	
ner å	t->1	
ner ö	v->1	
ner")	,->1	
ner, 	a->2	d->2	e->1	f->2	g->1	h->3	i->2	k->1	l->2	m->8	n->1	o->7	p->1	s->9	t->1	u->2	v->5	ä->1	å->1	
ner-p	r->10	
ner. 	E->1	Ä->1	
ner.(	I->1	
ner.-	 ->1	
ner..	 ->1	
ner.A	n->1	
ner.B	e->1	
ner.D	e->11	ä->2	
ner.F	ö->1	
ner.G	e->1	
ner.H	e->1	ä->1	
ner.I	 ->5	n->1	
ner.J	a->11	
ner.K	o->2	
ner.L	i->1	
ner.M	e->2	
ner.N	ä->1	
ner.R	e->1	
ner.S	å->1	
ner.T	i->1	
ner.U	n->1	
ner.V	a->1	i->4	
ner.Ä	r->1	v->1	
ner; 	o->1	
ner?-	 ->1	
ner?H	e->1	
ner?J	a->1	
ner?K	o->1	
ner?V	e->1	
nerNä	s->2	
nera 	E->1	d->4	e->1	h->1	i->2	o->1	p->1	s->3	v->2	
nerad	 ->3	.->2	e->20	
neral	d->17	i->1	s->2	
neran	d->7	
nerar	 ->9	,->1	
neras	 ->8	,->1	.->1	
nerat	 ->3	,->3	i->4	s->1	
nere 	a->1	k->1	
nere.	M->1	
nerel	l->16	
nerer	a->3	
nergi	 ->13	,->2	-->1	.->5	a->7	b->3	c->1	e->4	f->5	i->1	k->39	m->2	n->4	o->2	p->7	s->13	ä->1	å->1	
nerhe	t->46	
nerie	t->1	
nerin	g->63	
nerli	g->14	
nerna	 ->125	,->25	.->28	;->1	s->29	
ners 	a->4	e->1	f->2	i->1	l->1	s->1	u->1	ö->1	
nersh	i->1	
nersk	a->17	
nerst	a->2	
nerös	 ->2	a->1	t->1	
nes a	r->2	t->1	
nes b	a->1	e->1	y->1	
nes e	k->1	n->1	
nes f	r->2	ö->1	
nes i	n->1	
nes k	l->1	o->3	u->1	
nes m	a->1	y->1	
nes o	c->1	r->1	
nes s	t->1	v->1	
nes t	i->1	j->1	
nes u	p->1	
nes v	i->1	
nes, 	s->1	
neser	,->1	n->1	
nesis	k->8	
nesma	n->1	
nesmä	r->1	
nesrö	r->1	
ness 	i->1	
nesta	 ->1	
net "	E->1	
net a	t->1	
net f	ö->4	
net i	n->1	
net m	a->1	
net n	ä->1	
net o	b->1	c->1	
net p	å->2	
net s	k->1	
net t	a->1	
net u	n->1	
net v	i->1	
net ä	r->1	
net, 	a->1	f->1	n->1	o->1	s->1	u->1	
net. 	J->1	
net.D	e->4	
net.F	r->1	
net.I	n->1	
net.J	a->1	
net.M	i->1	
net.N	a->1	
net.O	m->1	
net.V	i->1	
netar	i->1	
netec	k->6	
netis	k->1	
nett 	h->1	
nett.	Ä->1	
nette	t->1	
netär	a->6	
neutr	a->2	
nevån	a->2	
nez a	n->1	
nezue	l->1	
nfall	e->2	
nfatt	a->6	n->6	
nfede	r->1	
nfekt	e->1	i->1	
nfere	n->170	
nfess	i->1	
nfide	n->2	
nfilt	r->1	
nfini	t->1	
nfinn	e->1	
nfisk	e->2	
nflik	t->16	
nflyk	t->1	
nflyt	a->11	e->1	
nford	r->2	
nform	a->72	e->18	
nfras	t->15	
nfred	e->1	
nfria	 ->1	
nfron	t->1	
nfråg	a->3	o->1	
nfärd	i->1	
nför 	-->1	2->1	B->2	D->1	E->4	K->3	S->1	a->6	b->2	d->15	e->19	f->5	h->1	i->4	j->2	k->3	l->1	m->8	o->1	p->5	r->4	s->5	t->2	u->7	v->4	Ö->1	ä->1	
nför,	 ->1	
nför.	D->1	V->1	
nför:	 ->1	
nföra	 ->39	n->23	s->6	
nförd	e->4	
nföre	t->5	
nförl	i->19	
nförs	 ->2	,->1	.->2	t->2	ö->1	
nfört	 ->4	r->3	s->2	
ng (1	9->1	
ng (E	G->1	
ng (a	r->2	
ng (r	e->1	
ng (å	t->1	
ng - 	S->1	d->3	g->1	i->1	m->1	o->3	s->1	
ng -,	 ->1	
ng 17	,->1	
ng 19	9->1	
ng 20	 ->1	0->1	
ng 37	/->1	
ng 60	0->1	
ng 68	5->1	
ng 80	 ->2	
ng De	t->1	
ng Ec	e->1	
ng Eu	r->1	
ng Fä	s->1	
ng IV	 ->2	
ng Ta	d->1	
ng VI	 ->1	
ng aj	o->1	
ng al	d->1	l->3	
ng an	n->5	t->3	
ng ar	b->1	
ng at	t->27	
ng av	 ->326	g->1	l->1	v->1	
ng ba	s->2	
ng be	a->1	k->1	r->1	s->2	t->2	
ng bi	l->1	
ng bl	a->1	i->2	
ng bo	r->1	
ng br	o->1	
ng by	r->1	
ng bö	r->5	
ng de	 ->1	l->1	n->2	s->1	t->4	
ng di	s->1	
ng dy	l->1	
ng dä	r->7	
ng e.	d->1	
ng ef	t->2	
ng el	l->9	
ng en	 ->7	d->1	
ng et	t->7	
ng ex	 ->1	i->1	
ng fi	e->1	n->4	
ng fo	r->1	
ng fr	a->4	ä->1	å->24	
ng fu	n->1	
ng få	r->2	
ng fö	l->1	r->88	
ng ga	r->1	
ng ge	n->8	
ng gj	o->1	
ng gl	ä->1	
ng gr	o->1	
ng gå	r->1	
ng ha	 ->2	d->1	n->3	r->19	
ng he	l->1	
ng ho	s->3	
ng hä	n->1	
ng hå	l->1	
ng i 	"->1	E->9	a->1	b->1	d->15	e->9	f->14	g->1	h->2	j->2	k->2	m->9	o->1	p->2	r->4	s->13	v->2	Ö->2	
ng ia	k->1	
ng in	f->2	g->1	n->5	o->12	r->1	t->11	
ng ir	r->1	
ng ja	g->1	
ng ka	n->7	
ng kn	a->1	
ng ko	m->15	n->3	p->1	
ng kr	ä->2	
ng ku	n->1	
ng le	d->1	
ng li	d->1	g->1	k->1	s->1	t->1	
ng lä	g->1	m->1	
ng lå	t->1	
ng ma	n->4	r->1	
ng me	d->30	l->12	n->3	r->1	
ng mi	g->1	s->1	
ng mo	t->10	
ng må	l->1	s->11	
ng ne	g->1	
ng ni	 ->4	
ng nr	 ->2	
ng nu	 ->1	
ng nä	r->3	
ng nö	d->1	
ng oc	h->149	k->1	
ng of	 ->1	t->1	
ng ol	j->1	
ng om	 ->32	.->1	ö->1	
ng pe	k->1	r->1	
ng pl	a->1	
ng po	l->1	
ng pr	o->4	
ng på	 ->48	,->1	.->2	b->1	v->1	
ng ra	d->1	t->1	
ng re	a->1	s->1	
ng ri	k->1	
ng rä	k->2	t->1	
ng rö	r->1	s->1	
ng sa	d->1	m->2	
ng se	n->1	r->1	
ng si	g->1	k->9	n->1	
ng sk	a->10	u->11	
ng so	m->108	
ng st	r->3	ä->1	å->1	ö->1	
ng sy	s->1	
ng sä	g->4	
ng så	 ->2	d->1	v->1	
ng ta	c->2	g->3	n->1	r->1	
ng ti	d->12	l->62	
ng tr	o->2	ä->1	
ng ty	d->1	v->1	
ng un	d->6	
ng up	p->2	
ng ur	v->1	
ng ut	a->7	k->1	o->1	s->1	t->1	
ng va	d->6	r->3	
ng ve	r->3	
ng vi	 ->7	d->4	l->3	s->2	
ng vo	r->1	
ng vä	g->2	
ng äg	n->1	
ng än	 ->3	d->3	
ng är	 ->38	o->1	
ng äv	e->2	
ng åt	 ->3	e->1	g->1	
ng ök	a->1	
ng öv	e->2	
ng!Ja	g->1	
ng" a	v->1	
ng" o	c->1	
ng", 	m->1	o->1	
ng".J	a->1	
ng".N	ä->1	
ng) i	 ->1	n->1	
ng) o	c->2	
ng).V	i->1	
ng)Nä	s->1	
ng, O	L->1	
ng, a	c->1	t->4	v->1	
ng, b	e->1	l->3	
ng, d	e->7	r->1	v->4	ä->1	
ng, e	f->7	l->1	n->5	t->2	
ng, f	a->1	i->1	o->1	r->5	ö->17	
ng, g	e->1	r->1	
ng, h	a->2	e->1	å->1	
ng, i	 ->8	n->6	
ng, k	a->1	o->3	u->1	
ng, l	e->2	i->1	å->1	
ng, m	a->1	e->14	i->2	o->2	
ng, n	u->2	ä->5	å->1	
ng, o	c->21	m->1	
ng, p	e->1	r->2	å->3	
ng, r	ä->1	å->1	
ng, s	a->3	j->1	k->3	o->12	p->2	t->1	ä->1	å->6	
ng, t	a->2	i->1	r->1	v->1	
ng, u	p->1	t->8	
ng, v	a->3	i->11	
ng, ä	r->2	v->2	
ng, å	t->3	
ng, ö	v->1	
ng-PM	 ->1	
ng. D	e->2	
ng. E	n->1	
ng. M	e->1	
ng. S	k->1	
ng.(A	p->1	
ng.. 	(->2	
ng..(	D->1	
ng.Al	l->3	
ng.An	s->1	
ng.Av	 ->3	s->1	
ng.Da	n->1	
ng.De	 ->6	n->11	s->1	t->48	
ng.Do	k->1	m->1	
ng.Dä	r->6	
ng.Ef	t->1	
ng.En	 ->1	d->1	l->3	
ng.Et	t->1	
ng.Eu	r->1	
ng.Fl	e->1	
ng.Fr	u->3	å->2	
ng.Fö	r->10	
ng.Ge	n->2	
ng.Ha	n->1	
ng.He	r->12	
ng.Hu	r->1	
ng.Hä	r->1	
ng.Hö	g->1	
ng.I 	d->8	e->1	f->1	s->1	v->2	
ng.In	g->2	
ng.Ja	g->32	
ng.Ka	n->1	
ng.Ko	m->6	n->1	s->1	
ng.Li	k->1	
ng.Lå	t->2	
ng.Ma	n->6	
ng.Me	d->1	n->3	
ng.My	n->1	
ng.Må	h->1	l->1	
ng.Na	t->1	
ng.Ni	 ->3	
ng.Nu	 ->2	
ng.Nä	r->2	
ng.Nå	j->1	
ng.Oc	h->7	
ng.Of	t->1	
ng.Om	 ->9	
ng.PP	E->1	
ng.Pa	r->1	
ng.Pr	o->1	
ng.På	 ->2	
ng.Re	f->1	
ng.Sa	m->1	
ng.Se	d->1	
ng.Sl	u->4	
ng.Så	 ->1	
ng.Ta	c->1	
ng.Ti	l->2	
ng.Tr	o->1	
ng.Va	d->1	
ng.Vi	 ->16	l->1	
ng.Vå	r->1	
ng.Är	 ->2	a->1	
ng: e	t->1	
ng: f	ö->1	
ng: i	n->1	
ng:De	t->1	
ng; d	e->1	
ng; e	n->1	
ng; f	ö->2	
ng?De	n->1	t->1	
ng?Hä	r->1	
ng?Ja	g->1	
ng?Ol	i->1	
ng?Ty	c->1	
ng?Är	 ->1	
nga -	 ->1	
nga a	l->1	n->13	r->2	v->21	
nga b	a->1	e->7	l->1	o->1	r->1	u->1	
nga c	e->1	
nga d	a->1	e->4	i->2	o->1	ä->1	å->2	
nga e	f->1	n->1	r->1	x->1	
nga f	a->3	e->1	l->4	r->5	ö->3	
nga g	e->1	o->2	r->2	å->3	
nga h	a->1	ä->1	
nga i	 ->3	c->1	n->1	
nga k	l->1	o->6	v->2	
nga l	a->1	e->1	i->1	
nga m	e->11	i->3	o->1	u->1	ä->3	å->1	ö->1	
nga n	a->1	y->4	ä->1	
nga o	c->4	e->1	k->1	l->3	m->3	s->1	
nga p	a->1	r->1	u->1	
nga r	e->6	å->2	
nga s	a->2	i->4	k->1	m->1	o->5	t->2	v->4	y->1	ä->1	
nga t	a->2	e->1	i->2	j->1	r->1	u->1	y->1	
nga u	n->2	t->2	
nga v	a->1	i->4	ä->2	
nga ä	m->1	n->5	r->1	
nga å	r->9	t->1	
nga ö	s->1	
nga, 	b->1	i->1	l->1	n->1	o->1	
nga.J	a->2	
nga.V	i->1	
ngade	 ->3	s->3	
ngage	m->9	r->9	
ngalu	n->3	
ngand	e->13	
ngar 	(->1	-->3	E->2	R->1	a->39	b->5	d->3	e->2	f->30	g->5	h->8	i->32	k->3	m->15	n->3	o->64	p->14	r->1	s->51	t->16	u->5	v->13	ä->11	å->2	ö->1	
ngar!	M->1	
ngar"	 ->1	
ngar)	.->1	
ngar,	 ->52	
ngar-	 ->1	
ngar.	 ->2	)->1	-->1	.->1	B->2	D->18	E->3	F->6	H->3	I->6	J->11	K->3	L->3	M->1	N->1	O->5	P->1	R->2	T->2	U->1	V->9	Ä->1	
ngar:	 ->7	
ngar;	 ->1	
ngar?	J->1	
ngare	 ->6	,->2	.->1	
ngari	k->15	
ngarn	a->159	
ngars	 ->3	
ngas 	a->2	b->1	e->1	f->1	i->1	k->1	p->1	r->1	t->1	v->1	ö->1	
ngas.	E->1	J->1	
ngast	e->2	
ngat 	l->1	o->1	s->1	
ngats	 ->1	
ngav 	h->1	
ngbro	 ->1	
ngd a	v->1	
ngd b	a->1	r->1	
ngd f	o->1	r->2	ö->2	
ngd i	n->1	
ngd n	i->1	
ngd o	c->2	l->1	t->1	
ngd s	a->1	o->1	
ngd y	t->1	
ngd ä	n->1	
ngd å	t->1	
ngda 	a->1	
ngde 	s->1	v->1	
ngden	 ->5	
ngder	 ->5	
ngdom	 ->1	a->7	s->7	
ngdpu	n->4	
ngdra	g->1	
ngdyr	k->1	
nge E	u->1	
nge a	l->1	n->2	t->1	
nge b	u->1	
nge d	e->4	
nge e	n->1	
nge h	a->2	
nge i	 ->1	n->1	
nge k	o->1	u->1	
nge m	a->1	
nge n	u->1	å->1	
nge o	c->4	r->1	
nge p	e->1	å->3	
nge s	e->5	o->5	ä->1	å->1	
nge t	r->1	
nge u	n->1	
nge v	a->2	e->1	i->2	
nge ä	n->1	
nge å	t->1	
nge, 	s->1	
ngefä	r->10	
ngel 	s->1	
ngeli	l->1	
ngeln	s->2	
ngels	e->1	k->9	m->1	
ngelä	g->22	n->1	
ngema	n->4	
ngen 	-->4	1->2	A->2	B->2	E->1	a->243	b->15	d->6	e->10	f->45	g->12	h->22	i->74	j->3	k->26	l->3	m->38	n->4	o->61	p->23	r->5	s->58	t->35	u->11	v->20	ä->19	ö->2	
ngen"	,->1	
ngen,	 ->80	
ngen.	 ->5	.->1	A->3	D->26	E->4	F->4	G->1	H->8	I->3	J->9	K->1	L->2	M->7	O->1	P->2	S->2	T->4	U->2	V->9	Ä->1	
ngen:	 ->4	
ngen;	 ->2	
ngen?	D->4	F->1	H->1	V->1	
ngenI	 ->1	
ngena	v->3	
ngenb	e->1	
ngenj	ö->2	
ngenk	o->1	
ngeno	m->1	
ngenr	e->1	
ngens	 ->23	,->1	t->1	
ngent	i->22	
ngenä	m->1	
nger 	-->1	2->1	S->1	a->1	b->1	d->2	f->5	h->3	i->2	k->1	l->1	m->1	o->3	p->2	s->13	t->4	u->1	v->3	ä->1	
nger,	 ->5	
nger.	D->1	E->1	N->1	
ngera	 ->20	!->1	,->2	.->6	n->6	r->17	t->4	
nges 	b->1	d->1	i->2	o->1	ä->1	
nges,	 ->2	
nges.	R->1	
ngesf	o->1	
nget 	a->4	b->1	e->1	f->1	g->2	i->4	k->2	m->5	n->1	o->2	s->13	t->5	u->3	v->3	ä->1	ö->1	
nget,	 ->1	
ngetd	e->1	
ngett	 ->1	
ngfal	d->15	
ngflö	d->1	
ngfon	d->1	
ngfor	s->20	
ngfri	s->1	
ngfru	t->1	
ngfun	k->1	
ngfär	d->1	g->1	
nggå 	l->1	
nggås	,->1	
ngigg	j->1	
ngigt	 ->1	
ngilt	i->1	
ngiva	n->2	r->3	
ngive	r->1	
ngivi	t->6	
ngivn	a->1	
ngkör	n->1	
nglew	o->2	
nglig	 ->2	,->1	a->26	e->3	h->1	t->4	
ngmet	a->6	
ngmål	,->1	
ngna 	a->6	å->2	
ngnin	g->44	
ngom 	u->1	ä->2	
ngom.	D->1	
ngpol	i->2	
ngra 	f->1	o->1	
ngran	d->2	
ngre 	a->2	b->1	f->6	g->1	h->1	i->2	k->7	n->2	o->3	p->5	r->1	s->8	t->7	u->1	v->4	ä->5	
ngre,	 ->1	
ngre.	F->1	I->1	M->1	N->1	R->1	V->1	
ngred	i->2	
ngrem	s->1	
ngrep	 ->1	p->10	
ngres	s->1	u->1	
ngrin	g->1	
ngrip	a->12	e->3	s->1	
ngrod	d->1	
ngrän	s->1	
ngs b	r->1	
ngs d	i->1	
ngs e	n->1	
ngs h	ä->1	
ngs k	u->1	
ngs p	o->1	
ngs s	k->3	
ngs v	i->1	
ngs- 	f->1	o->11	
ngsak	t->3	
ngsal	t->1	
ngsam	m->3	t->3	
ngsan	f->1	l->4	s->2	
ngsar	b->5	t->2	
ngsav	g->1	t->5	
ngsba	r->2	
ngsbe	d->1	h->1	l->1	s->3	t->1	v->4	
ngsbi	d->2	l->7	s->2	
ngsbo	l->2	r->1	
ngsce	n->5	
ngsch	e->8	
ngsdi	r->2	
ngsdo	k->1	
ngsdr	a->1	
ngsen	h->1	
ngser	b->1	
ngset	a->1	
ngsfa	k->1	r->2	s->4	
ngsfe	l->2	
ngsfi	e->30	n->1	
ngsfl	y->1	
ngsfo	n->21	r->1	
ngsfr	ä->2	å->13	
ngsfu	l->10	n->1	
ngsfö	r->232	
ngsgr	a->3	u->3	
ngsha	n->1	
ngsho	t->1	
ngsid	i->3	k->1	
ngsik	t->7	
ngsin	d->4	f->1	i->1	s->4	
ngska	p->1	
ngskl	a->2	i->1	
ngsko	a->2	m->24	n->134	r->2	s->8	
ngskr	a->13	i->1	
ngsku	r->1	
ngskv	o->1	
ngsla	g->1	n->1	
ngsli	g->1	n->2	s->47	v->9	
ngslo	g->1	
ngslä	g->3	n->3	
ngslö	s->5	
ngsma	j->1	k->1	r->2	
ngsme	d->2	k->2	t->3	
ngsmi	n->1	
ngsmo	d->2	m->1	n->1	t->1	
ngsmä	s->2	
ngsmå	l->4	
ngsmö	j->3	n->1	
ngsni	v->5	
ngsno	r->1	
ngsny	c->1	
ngsom	r->10	
ngsor	g->2	
ngspa	k->1	n->1	r->2	
ngspe	r->3	
ngspl	a->17	i->6	
ngspo	l->21	
ngspr	i->1	o->45	
ngspu	n->11	
ngspå	f->1	
ngsre	g->3	k->5	p->2	s->8	
ngsri	k->15	
ngsru	n->1	
ngsrä	d->1	t->1	
ngsrå	d->1	
ngssa	m->2	
ngsse	d->1	k->3	
ngssi	f->1	t->1	
ngssk	a->2	e->3	i->5	r->1	y->3	
ngssp	r->1	
ngsst	a->2	r->15	ö->2	
ngssy	s->24	
ngssä	k->1	l->6	t->8	
ngst 	a->1	f->1	p->1	
ngst.	V->1	
ngsta	 ->2	g->7	
ngste	n->3	
ngstj	ä->5	
ngstm	ä->2	
ngstr	ö->1	
ngstä	t->1	
ngsum	m->1	
ngsut	r->4	s->1	ö->1	
ngsve	r->4	
ngsvi	l->3	s->30	
ngsvä	n->1	r->5	v->1	
ngsvå	g->1	
ngsys	t->2	
ngsär	e->1	
ngsät	t->1	
ngsår	e->1	
ngsåt	g->5	
ngsöv	e->1	
ngt a	v->1	
ngt b	a->2	o->1	
ngt d	e->3	ä->2	
ngt f	r->3	
ngt h	a->1	j->1	
ngt i	f->6	n->1	
ngt k	v->2	
ngt m	e->5	
ngt n	i->1	ä->1	
ngt s	i->3	o->4	
ngt u	n->1	t->1	
ngt v	i->1	
ngt ö	v->1	
ngt, 	p->1	
ngt.D	e->1	
ngt.M	e->1	
ngt.V	a->1	
ngtar	 ->1	
ngter	a->8	
ngtgå	e->11	
ngtid	s->4	
ngton	 ->2	.->1	?->1	s->1	
ngtvä	t->4	
nguer	 ->2	
ngvar	i->6	
ngäld	 ->1	
ngå e	t->1	
ngå i	 ->5	
ngå s	o->1	å->1	
ngå.A	t->1	
ngåen	d->53	
ngång	e->1	
ngår 	d->1	e->1	f->1	i->5	o->3	p->1	s->1	ä->1	
ngår.	D->1	V->1	
ngått	 ->3	.->1	s->2	
ngör 	b->1	
ngöri	n->2	
nhamn	 ->1	
nhand	l->1	
nhang	 ->20	,->6	.->8	e->13	
nhas 	b->1	
nhedr	a->2	
nhems	k->2	
nhet 	a->4	f->3	i->9	k->4	l->1	m->2	o->16	r->1	s->4	t->1	ä->2	
nhet"	 ->2	
nhet,	 ->12	
nhet.	A->1	D->5	E->2	F->1	H->1	I->4	J->3	M->2	R->1	S->1	T->1	V->2	
nhete	n->50	r->61	
nhetl	i->36	
nhets	a->1	c->3	l->2	o->1	u->3	
nhill	 ->1	
nho f	ö->1	
nho p	å->1	
nho s	o->1	
nho v	ä->1	
nho. 	D->1	
nhos 	i->1	
nhund	r->1	
nhäll	i->32	
nhämt	a->6	
nhäng	a->3	e->1	i->1	
nhåll	a->3	n->52	
nhård	a->1	
nhöjd	e->4	
ni 19	6->1	9->5	
ni 20	0->2	
ni al	l->4	
ni an	v->1	
ni ar	b->1	
ni at	t->18	
ni av	s->1	
ni be	d->1	k->2	r->1	s->1	t->2	
ni bl	i->1	
ni br	y->1	
ni bä	t->1	
ni de	t->2	
ni di	s->1	
ni dä	r->1	
ni då	 ->3	
ni ef	t->1	
ni en	 ->1	
ni er	 ->1	k->1	
ni fi	c->1	
ni fr	a->2	å->1	
ni få	 ->1	
ni fö	r->10	
ni ge	 ->1	n->1	
ni gö	r->3	
ni ha	d->1	f->1	r->17	
ni he	r->1	
ni hä	n->1	v->1	
ni hå	l->1	n->1	
ni i 	L->1	d->1	å->1	
ni in	g->2	l->2	s->1	t->7	
ni ju	s->3	
ni ka	n->3	
ni ko	m->6	n->2	
ni ku	n->1	
ni kä	n->5	
ni le	v->1	
ni lä	g->1	
ni lö	s->1	
ni me	n->2	
ni må	s->1	
ni nu	 ->2	
ni nä	m->6	
ni oc	h->4	k->1	
ni om	 ->2	
ni os	s->1	
ni pa	r->1	
ni pe	k->1	
ni på	s->1	
ni ra	t->2	
ni re	d->2	
ni rä	t->1	
ni sa	d->9	m->2	
ni se	 ->1	r->3	
ni sj	ä->2	
ni sk	a->2	i->1	r->1	u->2	
ni sl	u->1	
ni so	m->2	
ni st	ä->1	ö->1	
ni sä	g->4	k->1	
ni ta	g->1	l->1	r->3	
ni ti	l->1	
ni to	l->1	
ni un	d->1	
ni up	p->3	
ni ut	v->1	
ni va	r->4	
ni ve	t->8	
ni vi	l->9	
ni vä	l->1	n->1	
ni vå	g->1	
ni är	 ->6	
ni äv	e->1	
ni ön	s->1	
ni, b	e->1	
ni, d	e->1	
ni, f	r->3	ö->1	
ni, h	e->4	
ni, i	n->1	
ni, m	e->1	
ni, o	m->2	r->1	
ni, t	i->1	
ni.(P	a->1	
ni.Al	l->1	
ni.Dä	r->1	
niali	s->1	
nicer	a->2	
nied 	(->1	
nied.	K->1	
niefu	s->1	
nien 	9->1	a->1	i->1	m->1	o->4	s->3	t->1	ä->2	
nien,	 ->4	
nien.	I->1	P->1	V->1	
nien?	E->1	
niens	 ->2	
nier 	-->4	a->2	e->1	f->1	h->1	k->1	o->1	s->2	t->1	ä->1	
nier,	 ->2	
nier.	K->1	
niera	 ->5	d->2	r->1	s->2	t->2	
nieri	n->1	
niern	a->5	
niers	 ->2	
niesk	i->2	
niet 	a->1	
niet.	A->1	H->1	
nifes	t->1	
nifrå	n->2	
nig h	a->1	
nig i	 ->1	
nig o	m->1	
niga 	i->1	o->1	
niga,	 ->1	
niga.	 ->1	J->1	
nighe	t->12	
nigt 	v->1	
nik D	e->1	
nik s	a->1	k->1	o->3	
nik u	t->1	
nik- 	o->1	
nika 	f->1	
nikat	i->16	
niken	 ->3	s->1	
niker	 ->1	,->1	n->1	
nikt 	k->1	
nilat	e->2	
nimal	i->1	
nimbu	s->1	
nimer	a->1	
nimib	e->2	
nimif	i->1	
nimii	n->1	
nimik	a->1	o->1	r->2	
nimil	ä->1	ö->1	
nimin	i->1	o->2	
nimir	e->5	
nimis	-->1	
nimor	u->1	
nimum	 ->4	
nimus	-->1	
ninde	l->1	
nindu	s->1	
niner	 ->1	
ning 	(->4	-->6	1->2	3->1	6->1	D->1	E->1	I->2	T->1	V->1	a->221	b->9	d->10	e->13	f->79	g->4	h->11	i->74	k->8	l->2	m->50	n->8	o->120	p->40	r->2	s->81	t->41	u->8	v->12	ä->24	å->2	ö->2	
ning"	,->1	.->1	
ning)	 ->1	N->1	
ning,	 ->125	
ning.	 ->1	(->1	.->2	A->7	D->44	E->5	F->9	G->2	H->10	I->8	J->22	K->7	L->2	M->7	N->1	O->8	P->3	R->1	S->6	T->1	V->9	Ä->1	
ning:	 ->3	D->1	
ning;	 ->2	
ning?	D->1	J->1	T->1	Ä->1	
ninga	r->308	
ningd	y->1	
ninge	n->580	
ningf	l->1	
ningo	m->4	
ningp	o->2	
ningr	e->1	
nings	 ->2	-->7	a->14	b->5	c->2	d->2	e->3	f->68	g->5	h->2	i->10	k->32	l->60	m->17	n->5	o->7	p->52	r->13	s->41	t->12	u->3	v->41	å->6	ö->1	
ningt	v->4	
ninsp	e->1	
ninvå	n->1	
nio V	i->1	
nio b	e->2	
nio f	ö->1	
nio l	ä->1	
nio m	i->5	å->2	
nio p	u->1	
nio t	i->1	
nio; 	d->1	
nion 	d->1	e->1	f->2	h->1	i->2	k->1	m->2	o->1	s->2	u->1	ä->1	
nion,	 ->5	
nion.	D->3	F->2	S->1	
niond	e->1	
nione	n->415	
nions	 ->1	-->1	f->1	m->2	n->1	s->1	u->1	
nipa.	E->1	
nipen	 ->1	
nippa	d->3	
niref	o->1	
nisat	i->42	o->1	
nisch	!->1	
niser	a->27	i->30	
nisk 	a->2	b->1	d->1	f->3	h->2	k->3	n->1	p->1	r->3	s->1	u->4	v->1	ö->2	
niska	 ->33	,->1	n->4	
nisko	f->2	h->3	l->3	r->82	s->1	
niskt	 ->8	
nism 	o->2	s->1	
nism,	 ->2	
nism.	D->1	J->1	
nisme	r->9	
nista	n->2	
niste	r->56	
nisti	s->7	
nistr	a->40	e->1	
nit d	e->1	
nit e	n->1	t->1	
nit f	r->2	
nit v	a->1	
nit, 	e->1	
nit.N	ä->1	
nitet	 ->5	,->4	.->2	:->1	e->2	
nitia	t->80	
nitie	r->2	
nitio	n->14	
nitis	k->1	
nitiv	 ->2	a->2	t->5	
nitor	i->1	
nits 	e->1	n->1	o->1	p->1	s->1	t->2	
nits,	 ->1	
nitt 	2->1	i->1	l->2	s->1	t->1	u->1	
nitt,	 ->1	
nitte	n->2	t->3	
nittl	i->1	
nitts	r->1	
nitud	 ->1	
nitum	.->1	
nitz 	i->1	
nitär	t->1	
nium 	b->1	s->1	
nium!	D->1	
nium.	A->1	S->1	
niver	s->4	
nivå 	-->1	a->3	d->1	f->5	g->2	h->1	i->4	m->4	n->1	o->7	p->2	s->9	u->3	v->1	ä->2	
nivå,	 ->13	
nivå.	A->1	B->1	D->7	F->1	G->1	H->2	J->4	M->1	N->1	P->1	V->1	
nivå;	 ->1	
nivå?	S->1	
nivåe	r->14	
nivåg	r->3	
nivån	 ->7	.->4	
nié u	t->1	
nj fö	r->2	
nj mo	t->1	
nj.De	 ->1	
nje (	B->1	
nje m	e->5	
nje o	c->1	
nje s	o->4	
nje.G	e->1	
nje.J	a->1	
njen 	b->1	h->1	i->1	
njen.	D->1	
njer 	9->1	b->1	d->1	e->1	f->7	g->1	i->5	k->2	n->3	o->5	s->5	u->1	v->1	ä->1	å->1	
njer"	.->1	
njer,	 ->6	
njer.	H->1	M->1	V->1	
njer:	 ->1	
njern	a->31	
njor 	o->1	
njunk	t->1	
njute	r->1	
njutn	i->1	
njuve	l->1	
njämk	a->1	
njäre	r->1	
njör 	-->2	
nk ba	r->1	
nk en	 ->1	
nk ho	n->1	
nk på	 ->1	
nk ra	k->1	
nk ti	l->1	
nk ut	a->1	
nk vä	g->1	
nk" f	ö->1	
nk- e	l->1	
nk.De	t->1	
nka a	r->2	t->1	v->1	
nka b	e->1	
nka d	e->2	
nka e	f->1	n->1	
nka h	j->1	o->1	
nka m	i->2	
nka n	å->1	
nka o	c->1	s->1	
nka p	å->16	
nka s	a->1	i->6	
nka v	a->1	
nka ö	v->2	
nka, 	s->1	
nka.E	n->1	
nka.Å	 ->1	
nkall	a->9	
nkand	e->288	
nkar 	f->1	k->2	o->4	s->3	
nkar,	 ->1	
nkar.	E->1	J->1	V->2	
nkara	?->1	
nkarn	a->2	
nkas 	t->1	v->1	
nkas,	 ->1	
nkata	s->1	
nkbar	a->2	h->1	t->1	
nke a	t->1	
nke l	e->1	
nke o	c->1	
nke p	å->40	
nke r	ö->1	
nke t	i->2	
nke ä	r->2	
nke, 	h->1	n->1	
nkeba	n->1	
nkefr	i->1	
nkegå	n->1	
nkel 	a->2	b->1	f->1	k->1	o->2	ä->2	
nkel.	E->1	V->1	Ä->1	
nkel:	 ->2	
nkelm	a->1	
nkeln	 ->1	,->1	
nkelr	i->1	
nkelt	 ->28	
nkelv	ä->2	
nken 	-->1	a->2	b->1	m->4	o->4	p->5	s->1	t->1	u->1	
nken,	 ->2	
nken.	M->1	
nken:	 ->1	
nkens	 ->1	
nkepo	l->1	
nker 	a->2	b->1	d->1	f->1	g->3	i->3	j->3	k->1	m->3	n->3	o->3	p->12	r->4	s->4	u->1	
nker,	 ->2	
nkern	 ->2	s->1	
nkers	 ->1	
nkerä	g->1	
nkesi	s->1	
nkfar	t->7	
nkfor	d->1	
nkför	v->1	
nkire	r->1	
nkit 	f->1	t->1	
nkla 	d->1	e->1	f->2	n->1	o->3	s->2	
nklad	e->1	
nklag	a->1	e->3	
nklar	 ->1	,->1	e->3	
nklas	 ->1	t->2	
nklat	s->1	
nklig	h->5	
nklin	g->1	
nklud	e->4	
nklus	i->17	
nkna 	t->1	
nknad	e->1	
nknar	 ->1	
nknat	 ->1	
nknin	g->15	
nknyt	n->1	
nko.T	y->1	
nkole	n->1	
nkoml	i->3	
nkomm	e->1	
nkomp	e->3	
nkoms	t->12	
nkons	e->1	
nkont	r->2	
nkonv	e->3	
nkopp	l->1	
nkra 	d->1	
nkrad	 ->1	e->2	
nkraf	t->22	
nkrar	 ->1	.->1	n->3	
nkren	g->2	
nkret	 ->18	:->1	a->37	i->2	
nkrik	e->39	
nkris	e->1	
nkräk	t->1	
nks o	c->2	
nks t	i->1	
nksam	h->2	
nksch	e->1	
nksek	r->1	
nkt (	8->2	
nkt -	 ->1	,->1	
nkt 1	 ->1	,->1	1->1	
nkt 2	 ->2	6->1	
nkt 4	 ->2	
nkt 5	,->1	
nkt 6	 ->1	
nkt 7	 ->1	
nkt D	 ->1	
nkt a	b->1	t->5	
nkt b	e->1	
nkt d	)->1	ä->3	
nkt e	)->1	t->1	
nkt f	e->1	r->1	y->1	ö->3	
nkt g	ä->3	ö->1	
nkt h	a->2	i->1	u->1	ä->1	
nkt i	 ->10	n->6	
nkt k	l->1	o->1	
nkt m	o->1	y->3	
nkt n	ä->2	
nkt o	c->4	m->2	
nkt p	å->29	
nkt r	i->1	
nkt s	i->1	k->1	o->19	
nkt t	r->1	v->1	
nkt u	t->1	
nkt v	a->1	i->2	
nkt ä	n->1	r->7	
nkt, 	"->1	d->1	e->1	f->1	m->2	n->1	o->2	s->4	t->1	
nkt. 	D->1	
nkt.A	v->1	
nkt.D	e->4	i->1	
nkt.I	 ->1	
nkt.M	a->1	e->1	i->1	
nkt.N	u->1	å->1	
nkt.P	r->1	
nkt.T	a->1	i->1	
nkt.V	a->1	i->2	å->1	
nkt: 	J->1	V->1	
nkt?E	u->1	
nkta 	a->2	e->1	f->3	
nkta,	 ->1	
nkta.	J->1	
nkte 	p->1	s->2	
nkten	 ->66	,->10	.->12	
nkter	 ->50	,->8	.->11	:->2	?->2	n->13	
nktio	n->41	
nktiv	a->1	
nkts 	a->1	e->2	i->1	
nktsp	r->1	
nktur	e->1	
nkurr	e->285	
nkänn	e->1	
nköp 	a->1	
nköps	b->1	
nkörs	p->1	
nlagt	 ->1	
nlamp	o->1	
nland	 ->1	,->4	.->2	
nlar 	f->1	
nlarn	a->1	
nleda	 ->21	,->1	n->5	s->4	
nledd	e->10	
nlede	r->8	
nledn	i->57	
nleds	 ->5	
nlett	 ->3	s->10	
nlig 	a->2	d->2	f->2	m->3	n->1	s->2	t->1	u->1	
nlig,	 ->1	
nlig.	J->1	
nliga	 ->30	,->2	.->1	r->2	s->1	
nlige	n->17	
nligg	a->1	
nligh	e->37	
nligt	 ->135	!->1	,->1	.->1	v->1	
nlita	t->1	
nlysn	i->1	
nlägg	 ->13	.->1	e->4	n->14	
nlämn	a->1	i->4	
nländ	e->1	s->5	
nlänk	a->1	
nlänt	.->1	
nlåst	a->1	
nlåta	 ->1	
nlöpa	 ->1	n->1	
nlöpe	r->3	
nlös 	k->1	
nmanö	v->1	
nmark	 ->17	,->3	.->4	s->2	
nmäla	 ->2	n->1	
nmäld	a->1	
nmäle	r->1	
nmäln	i->12	
nmäls	 ->2	
nmält	 ->1	
nmärk	a->1	n->10	t->1	
nmäss	i->2	
nmöte	t->2	
nn de	 ->1	
nn eu	r->1	
nn oc	h->1	
nn ti	l->1	
nn är	 ->1	
nn, d	e->1	
nn, e	t->1	
nn-gr	u->1	
nna -	 ->2	
nna E	u->1	
nna T	e->1	u->1	
nna a	k->1	m->2	n->15	r->5	s->1	t->6	v->4	
nna b	a->6	e->16	i->5	l->4	o->1	r->3	u->4	y->4	ä->1	ö->1	
nna c	a->1	e->1	
nna d	a->3	e->39	i->4	r->2	ö->1	
nna e	f->3	k->1	l->1	n->12	r->2	t->1	u->1	
nna f	a->4	i->2	o->3	r->71	u->3	å->6	ö->42	
nna g	a->4	e->25	r->7	å->5	ö->8	
nna h	a->4	e->1	i->1	j->2	o->2	y->1	ä->3	å->1	ö->1	
nna i	 ->1	d->1	f->1	g->1	k->1	n->21	
nna j	o->1	
nna k	a->26	l->1	o->27	r->2	u->1	v->6	ä->3	
nna l	a->2	e->4	i->2	u->1	y->1	ä->4	å->1	ö->8	
nna m	a->6	e->8	i->3	o->2	u->2	y->8	ä->1	å->3	ö->4	
nna n	e->1	y->3	å->2	
nna o	c->3	j->1	l->3	m->12	p->1	r->11	s->6	
nna p	a->4	e->1	l->3	o->6	r->26	u->9	å->4	
nna r	a->6	e->54	i->5	o->2	ä->5	ö->2	
nna s	a->3	e->8	i->17	j->5	k->7	l->3	m->2	n->1	o->4	p->6	t->28	u->2	v->2	y->2	ä->5	å->3	
nna t	a->6	e->7	i->9	o->1	r->2	v->1	y->13	ä->3	
nna u	l->1	n->5	p->11	r->1	t->18	
nna v	a->11	e->4	i->20	ä->5	å->4	
nna y	r->1	t->1	
nna ä	n->4	r->2	
nna å	k->1	s->1	t->13	
nna ö	d->2	k->1	p->1	v->4	
nna, 	B->1	i->1	v->1	ö->1	
nna. 	D->1	Å->1	
nna.-	 ->1	
nna.D	ä->1	
nna.J	a->3	
nna.O	m->1	
nna.U	t->1	
nna.V	i->2	
nna.Ä	r->1	
nna?S	v->1	
nnabi	s->1	
nnade	 ->6	
nnaga	v->3	
nnage	 ->1	r->1	t->1	
nnagi	v->3	
nnaki	s->2	
nnala	g->1	
nnamb	a->1	
nnan 	E->3	a->3	b->3	c->1	d->11	e->2	f->2	g->1	h->1	i->1	j->3	k->1	m->8	n->1	o->3	p->1	r->3	s->9	t->1	v->16	å->2	
nnan,	 ->4	
nnan.	L->1	
nnand	e->28	
nnans	t->2	
nnar 	d->2	i->3	k->1	l->1	n->1	o->1	r->1	v->1	
nnare	p->1	
nnars	 ->18	,->1	
nnas 	a->5	d->3	e->12	h->1	i->3	k->4	l->1	m->4	n->7	o->5	p->1	r->1	t->4	ä->1	
nnas!	E->1	
nnas,	 ->2	
nnas.	D->1	M->1	Å->1	
nnat 	-->1	E->1	I->1	a->2	b->5	d->4	e->1	f->14	g->5	h->2	i->7	j->1	k->8	l->4	m->2	o->3	p->4	r->3	s->11	t->5	u->6	v->4	ä->13	å->3	ö->1	
nnat,	 ->1	
nnat.	D->1	G->1	K->1	Ä->1	
nndra	g->1	
nne F	o->1	
nne a	n->1	t->2	v->1	
nne f	r->1	ö->3	
nne h	a->2	j->1	ö->1	
nne n	ä->1	
nne o	c->1	
nne p	å->2	
nne s	o->1	
nne t	i->1	
nne ä	r->2	
nne å	k->1	
nne! 	N->1	
nne, 	g->1	k->1	n->1	t->1	ä->1	
nne.D	e->1	
nne.J	a->1	
nneba	r->1	
nnebo	e->1	
nnebä	r->108	
nnebö	r->7	
nnedo	m->1	
nnefa	t->6	
nneha	r->2	v->1	
nnehå	l->78	
nnehö	l->4	
nnela	g->1	
nneli	g->1	
nneln	,->1	.->1	
nnelt	r->1	
nnen 	J->1	a->10	e->2	f->2	h->2	i->4	j->1	k->3	m->2	n->2	o->2	p->1	s->7	
nnen,	 ->2	
nnen.	B->1	D->1	J->2	O->1	
nnena	 ->1	
nnens	 ->11	
nner 	E->1	J->1	K->1	a->7	b->1	d->12	e->3	f->3	g->2	i->9	j->3	k->1	m->12	n->2	o->18	r->1	s->22	t->18	u->1	v->8	ä->2	ö->1	
nner,	 ->5	
nner.	 ->1	.->1	J->1	M->1	U->1	
nnerh	e->46	
nnerl	i->12	
nners	t->2	
nnes 	a->3	b->2	e->1	f->3	i->1	k->4	m->2	o->2	s->2	t->2	u->1	v->1	
nnes,	 ->1	
nnesm	a->1	ä->1	
nnesr	ö->1	
nnet 	m->1	
nnet.	D->1	F->1	
nnete	c->6	
nnevå	n->2	
nnhet	 ->1	
nnief	u->1	
nnien	 ->9	,->2	.->2	s->1	
nnier	 ->3	.->1	n->1	
nnies	k->2	
nniet	 ->1	.->2	
nnig 	h->1	o->1	
nniga	.->1	
nnigh	e->3	
nnigt	 ->1	
nning	 ->19	)->1	,->3	.->3	a->5	d->1	e->15	f->1	p->2	r->1	s->24	t->4	
nnisk	a->7	o->91	
nnit 	d->1	e->2	f->2	v->1	
nnit,	 ->1	
nnit.	N->1	
nnits	 ->7	,->1	
nnium	 ->1	!->1	.->1	
nnivå	 ->1	
nnlan	d->1	
nnlar	 ->1	n->1	
nnlig	a->2	
nnlys	n->1	
nnlän	d->1	
nnock	 ->12	,->6	.->3	s->3	
nnoli	k->9	
nnopr	o->2	
nnor 	a->1	e->1	f->1	i->10	o->14	s->9	t->1	
nnor,	 ->3	
nnor.	D->1	F->2	J->1	
nnor?	H->1	
nnorl	u->2	
nnorn	a->5	
nnors	 ->10	t->2	
nnova	t->6	
nns 2	4->1	
nns G	e->1	
nns S	O->1	
nns a	b->1	l->4	n->4	r->3	t->3	u->1	v->1	
nns b	e->3	i->1	l->1	
nns c	i->1	
nns d	a->1	e->51	o->1	ä->6	
nns e	k->1	m->1	n->32	t->18	x->1	
nns f	a->3	l->3	o->6	r->2	å->1	ö->10	
nns g	a->1	e->1	o->1	r->1	
nns h	i->1	o->1	u->1	ä->2	
nns i	 ->19	n->24	
nns j	u->2	
nns k	v->3	
nns l	u->1	
nns m	a->1	e->5	i->1	o->1	y->2	ä->1	å->11	ö->1	
nns n	a->1	i->1	u->2	ä->1	å->15	
nns o	c->7	l->1	m->2	s->1	t->1	
nns p	r->3	å->5	
nns r	e->5	i->4	ä->1	
nns s	a->2	e->1	k->3	m->1	o->1	t->2	ä->1	å->4	
nns t	i->8	r->1	v->6	
nns u	t->1	
nns v	e->1	i->4	
nns y	t->2	
nns ä	n->1	r->1	v->1	
nns å	t->1	
nns ö	k->1	v->1	
nns, 	b->1	d->1	m->1	
nns.D	e->2	ä->1	
nns.E	n->1	
nns.J	a->1	
nns.M	y->1	
nns.V	a->1	
nnsak	a->1	
nnsam	m->2	t->1	
nnska	p->1	
nnu a	l->1	
nnu e	n->9	t->3	
nnu f	l->1	
nnu h	å->2	ö->4	
nnu i	n->32	
nnu m	e->7	i->1	
nnu n	å->1	
nnu p	å->1	
nnu s	k->1	m->1	t->6	v->1	å->1	
nnu v	i->2	
nnu ä	l->1	
nnu.D	e->1	
nnu.K	o->2	
nnu.V	i->1	
nnu; 	i->1	
nnytt	i->2	
nnäer	;->1	
nnämn	d->2	
no Le	o->1	
no Pr	o->2	
no i 	e->1	
no ko	m->1	
no oc	h->1	
no om	 ->1	
no un	d->1	
no, T	a->1	
no, m	e->1	
no.Ja	g->1	
no.Or	d->1	
nock 	f->1	h->2	i->1	k->4	l->1	m->1	n->1	v->1	
nock,	 ->6	
nock.	 ->1	J->1	K->1	
nocks	 ->3	
nodla	r->2	
nodli	n->1	
nog a	t->3	
nog b	a->1	
nog d	e->1	i->1	
nog h	a->2	
nog i	 ->1	
nog k	a->1	
nog n	o->1	
nog o	c->1	
nog p	å->1	
nog ö	k->1	
nog, 	i->1	
nog.M	e->1	ö->1	
noga 	a->1	f->4	m->2	p->1	s->1	
noga,	 ->1	
noga.	J->1	V->1	
noggr	a->12	
nogra	f->2	
noise	 ->1	
nokul	t->3	
nolik	a->2	h->2	t->5	
noll,	 ->1	
nolln	i->1	
nollr	i->1	
nolog	i->3	
nom -	 ->1	
nom 2	8->1	
nom 5	b->1	
nom A	m->1	
nom D	i->1	
nom E	M->1	U->11	u->27	
nom F	ö->1	
nom G	e->1	
nom I	r->1	
nom L	i->1	
nom S	E->1	c->1	
nom V	ä->1	
nom W	i->1	
nom a	g->1	l->4	n->2	r->1	t->106	v->1	
nom b	a->1	e->2	i->2	u->1	ä->1	ö->1	
nom d	e->64	i->5	ä->1	
nom e	g->1	k->1	l->1	n->23	r->1	t->11	
nom f	e->1	i->1	l->1	r->1	u->1	y->1	ö->8	
nom g	e->9	
nom h	a->3	e->2	u->1	ä->1	
nom i	 ->2	n->8	
nom j	o->3	ä->1	
nom k	a->1	o->22	r->1	u->2	
nom l	a->1	i->1	y->1	ä->2	
nom m	e->3	i->3	y->6	å->2	
nom n	a->2	ä->1	å->2	
nom o	c->2	l->1	m->10	r->1	
nom p	o->2	r->3	u->1	å->2	
nom r	a->51	e->1	i->3	å->4	
nom s	a->3	e->2	i->1	j->1	k->2	o->2	p->1	t->6	ä->2	å->1	
nom t	a->1	i->9	r->1	v->2	
nom u	n->15	p->3	t->4	
nom v	a->1	e->1	i->10	ä->1	å->4	
nom y	t->1	
nom ä	n->1	r->1	
nom å	r->1	t->3	
nom ö	r->1	v->6	
nom, 	a->1	t->1	u->1	
nom. 	H->1	
nom.H	e->1	u->1	
nom.J	a->1	
nom.M	e->1	
nom.V	i->1	
nomar	b->2	
nombl	i->5	
nombr	o->2	
nomdr	i->6	
nomen	 ->1	,->2	.->1	e->2	
nomer	 ->1	
nomeu	r->1	
nomfö	r->161	
nomgi	c->1	
nomgr	i->4	
nomgå	 ->1	.->1	n->3	r->4	t->2	
nomi 	-->1	a->1	m->5	o->12	ä->1	
nomi,	 ->2	
nomi.	D->2	F->1	
nomi?	 ->1	
nomie	r->8	
nomin	 ->20	,->2	.->5	e->3	s->3	
nomis	k->215	t->4	
nomlä	s->2	
nområ	d->1	
nomsk	i->1	
nomsl	a->3	
nomsn	i->11	
nomsy	r->3	
nomtä	n->1	
non e	f->1	
non f	ö->2	
non o	c->1	
non, 	i->1	
non.E	n->1	
non?K	a->1	
noner	.->1	
nonym	 ->2	.->1	a->1	i->1	
nopol	 ->8	,->1	.->1	f->3	i->3	s->1	
nopro	g->2	
nor a	t->1	
nor e	l->1	
nor f	a->1	
nor i	 ->7	n->3	
nor o	c->14	
nor s	k->1	o->7	t->1	
nor t	i->1	
nor, 	g->1	s->2	
nor.D	e->2	
nor.F	ö->3	
nor.J	a->2	
nor.V	å->1	
nor?H	u->1	
norda	m->4	
norde	u->1	
nordi	r->2	s->1	
nordk	u->1	
nordl	i->4	
nordn	a->4	i->5	
nordt	y->1	
nordv	ä->1	
norer	a->4	
norit	e->22	
norlu	n->2	
norm 	d->1	f->2	k->2	o->1	ö->1	
norma	 ->17	.->1	l->11	t->2	
norme	r->32	
normt	 ->7	
norna	 ->3	.->1	s->2	
norr?	V->1	
norra	 ->4	
nors 	d->5	l->1	p->1	r->1	s->1	ö->1	
norst	ä->2	
nos h	a->1	
nos i	n->1	
nos o	r->1	
nos t	a->1	
nos! 	J->1	
nos, 	a->1	h->1	
notan	;->1	
noter	a->27	n->1	
notis	 ->1	
notti	 ->1	
novat	i->6	
novem	b->11	
nover	a->1	i->2	
now-h	o->1	
npass	a->10	n->4	
nporn	o->2	
nprin	c->2	
nprob	l->1	
nprän	t->1	
npunk	t->31	
npå d	e->1	
nr 1 	f->1	
nr 12	 ->1	4->1	
nr 17	6->2	
nr 28	 ->1	
nr 29	 ->1	
nr 30	 ->1	
nr 31	 ->1	
nr 32	.->1	
nr 33	 ->1	2->1	
nr 35	 ->1	
nr 36	 ->1	
nr 37	 ->1	
nr 38	 ->1	
nr 39	 ->1	
nr 40	 ->1	
nr 41	 ->1	
nr 42	 ->1	
nr 43	.->1	
nr 44	 ->1	
nr 45	 ->1	
nr 46	 ->1	
nr 5 	f->1	
nr 6 	f->1	
nr 7.	F->1	
nr 8 	f->1	
nr 9 	f->1	
nra k	o->1	
nra o	m->10	
nrad 	A->1	
nrar 	o->1	
nras 	a->1	
nre a	n->2	
nre e	u->2	
nre g	r->1	
nre m	a->69	
nre v	a->8	ä->1	
nrege	l->1	
nreni	n->1	
nresa	 ->3	,->1	n->1	
nresu	r->1	
nrike	s->13	
nrikt	a->20	n->24	
nry F	o->1	
nryms	 ->1	
nrätt	a->54	n->2	
nråde	n->1	
nröja	 ->4	s->1	
nröjt	s->1	
nrött	.->1	
ns - 	a->1	
ns 24	 ->1	
ns 28	:->1	
ns BN	I->2	P->1	
ns EU	-->1	
ns Eu	r->2	
ns Ge	n->1	
ns He	l->1	
ns Is	r->1	
ns SO	L->1	
ns VD	 ->1	
ns XX	V->1	
ns ab	s->2	
ns ad	m->1	
ns ag	e->2	
ns ak	t->1	
ns al	l->10	t->1	
ns am	b->1	
ns an	a->1	d->7	f->1	g->1	l->1	n->1	s->11	t->1	v->1	
ns ar	b->15	g->1	k->1	
ns at	t->11	
ns au	k->1	
ns av	 ->8	g->3	s->1	
ns ba	c->1	r->1	
ns be	f->3	g->7	h->6	r->1	s->6	t->23	v->1	
ns bi	d->1	l->1	
ns bl	.->1	o->2	
ns br	i->1	
ns bu	d->7	
ns by	r->1	
ns bä	s->1	
ns bå	d->2	
ns ce	n->1	
ns ci	r->1	
ns da	g->12	
ns de	 ->3	b->6	l->3	m->3	n->3	t->48	
ns di	r->5	
ns do	c->1	k->3	m->2	
ns dä	r->7	
ns dö	d->1	
ns ef	f->3	t->3	
ns eg	e->5	n->1	
ns ek	o->18	
ns el	l->1	
ns em	b->1	e->1	
ns en	 ->32	d->2	h->3	s->1	
ns et	t->18	
ns eu	r->1	
ns ex	e->1	i->1	p->1	t->1	
ns fa	k->2	l->1	m->2	n->1	r->3	
ns fe	l->1	m->1	
ns fi	n->3	s->1	
ns fl	e->4	o->1	
ns fo	n->1	r->9	t->1	
ns fr	a->8	i->2	ä->2	å->9	
ns fu	n->3	
ns fy	r->1	
ns få	 ->1	
ns fö	l->2	r->76	
ns ga	r->1	s->1	
ns ge	m->8	n->4	r->1	
ns go	d->3	
ns gr	a->2	u->5	ä->2	ö->1	
ns gä	r->1	
ns gå	n->1	
ns ha	m->3	n->3	v->1	
ns he	l->1	
ns hi	n->1	s->2	t->2	
ns ho	s->1	t->1	
ns hu	r->1	v->1	
ns hä	l->2	n->2	r->4	
ns hå	l->1	
ns i 	A->1	E->3	F->1	I->1	a->1	b->3	d->3	e->2	f->3	r->2	s->4	v->3	ä->2	
ns id	é->1	
ns ik	r->1	
ns im	m->1	
ns in	f->1	g->18	i->2	k->1	l->1	n->4	r->5	s->15	t->21	v->3	
ns jo	r->2	
ns ju	 ->1	r->3	v->1	
ns ka	n->2	
ns ko	l->3	m->4	n->23	r->1	
ns kr	a->2	i->2	
ns ku	l->3	m->1	n->1	
ns kv	a->6	
ns kä	n->1	r->1	
ns la	g->9	n->4	
ns le	d->1	g->1	
ns li	g->1	k->1	v->2	
ns lj	u->1	
ns lo	p->2	
ns lu	c->1	
ns lä	g->2	m->1	n->5	s->1	
ns lö	f->1	
ns ma	n->3	r->2	t->1	
ns me	d->53	l->10	s->1	t->3	
ns mi	l->2	n->3	s->1	
ns mo	n->1	t->4	
ns my	c->4	
ns mä	n->1	
ns må	l->6	n->11	
ns mö	j->4	r->1	
ns na	m->4	t->2	
ns ne	g->1	
ns ni	 ->1	v->2	
ns nu	 ->2	v->6	
ns ny	f->1	
ns nä	r->2	
ns nå	g->16	
ns nö	d->1	
ns ob	e->3	
ns oc	h->30	k->6	
ns od	j->1	
ns oi	n->2	
ns ol	i->2	
ns om	 ->21	)->1	.->4	b->1	f->2	r->5	
ns or	d->10	g->2	o->3	
ns os	ä->1	
ns ot	i->2	v->1	
ns pa	r->10	s->1	
ns pe	n->1	r->1	
ns pl	a->2	
ns po	l->10	p->1	s->1	ä->1	
ns pr	a->1	e->3	i->5	o->4	
ns på	 ->9	p->1	
ns ra	n->1	p->15	
ns re	a->1	d->4	f->2	g->23	k->1	p->1	s->9	
ns ri	k->4	s->4	
ns ro	c->1	l->7	
ns ru	t->1	
ns rä	k->6	t->12	
ns rå	d->1	
ns rö	r->1	
ns sa	k->2	m->14	
ns sc	i->1	
ns se	g->1	k->2	n->1	x->1	
ns si	d->17	n->1	t->2	
ns sj	ä->1	
ns sk	a->3	i->1	o->2	u->3	y->1	ä->3	ö->1	
ns sl	a->2	u->5	
ns sm	å->1	
ns sn	a->3	
ns so	c->3	m->14	
ns sp	e->3	å->1	
ns st	a->4	e->1	o->3	r->15	u->1	y->1	ä->3	å->4	ö->6	
ns sv	a->3	
ns sy	n->3	
ns sä	k->2	n->1	r->3	t->3	
ns så	 ->1	d->1	l->2	
ns ta	k->2	l->1	n->1	
ns te	k->1	n->2	r->4	x->2	
ns ti	d->2	l->13	
ns tj	ä->7	
ns to	t->1	
ns tr	a->1	e->1	o->4	
ns tu	r->1	
ns tv	i->2	å->4	
ns un	i->1	
ns up	p->8	
ns ur	s->5	
ns ut	a->1	b->1	f->3	g->1	m->4	r->3	s->1	t->16	v->16	
ns va	d->1	r->3	t->1	
ns ve	r->9	t->1	
ns vi	 ->1	c->1	d->3	k->5	l->5	n->1	s->2	t->5	
ns vo	l->1	
ns vä	g->6	k->1	l->2	n->1	r->3	
ns yt	a->1	t->8	
ns äg	a->3	g->1	
ns än	d->4	
ns är	 ->7	
ns äv	e->1	
ns ål	d->2	
ns år	h->1	l->2	
ns ås	i->3	
ns åt	e->1	g->3	m->1	
ns öd	e->3	
ns ök	a->2	
ns ör	e->1	
ns öv	e->9	
ns!Vi	 ->1	
ns, b	l->1	ö->1	
ns, d	e->5	å->1	
ns, e	l->1	
ns, f	r->4	
ns, j	a->1	
ns, m	e->2	i->2	ä->1	
ns, n	ä->2	å->1	
ns, o	c->8	m->3	
ns, p	a->1	
ns, s	o->4	
ns, t	y->1	
ns, v	i->1	ä->1	
ns, ä	r->2	
ns- o	c->6	
ns.De	t->10	
ns.Dä	r->2	
ns.En	 ->1	
ns.Eu	r->1	
ns.Fö	r->1	
ns.I 	s->1	
ns.Ja	g->3	
ns.Lå	t->1	
ns.Ma	n->1	
ns.Me	n->1	
ns.My	n->1	
ns.Oa	v->1	
ns.So	m->1	
ns.Va	r->1	
ns/de	n->1	
ns: h	ö->1	
ns; v	i->1	
ns?.H	e->1	
ns?Et	t->1	
ns?Ja	,->1	
nsa a	n->2	
nsa d	e->2	
nsa m	i->1	
nsa p	a->1	
nsa s	i->1	t->2	
nsa t	i->1	v->1	
nsa u	p->2	t->1	
nsa, 	f->1	
nsad 	a->1	d->2	e->2	g->1	o->2	s->1	t->4	
nsad,	 ->1	
nsad.	D->1	J->1	V->1	
nsade	 ->9	.->1	
nsaff	ä->2	
nsaka	r->1	
nsam 	a->4	b->1	c->1	d->4	e->3	f->2	g->1	h->1	i->2	l->2	m->6	p->1	r->6	s->10	t->1	u->1	v->2	å->2	
nsam,	 ->1	
nsaml	i->8	
nsamm	a->134	e->1	
nsamr	ä->1	
nsamt	 ->26	,->1	.->1	
nsana	l->1	
nsand	e->3	
nsar 	d->1	e->1	m->1	o->1	t->1	u->1	
nsarb	e->8	
nsas 	m->1	t->4	
nsat 	a->1	b->1	f->1	i->1	m->1	s->1	t->1	
nsat.	D->1	F->1	H->1	
nsati	o->3	
nsats	 ->6	,->4	.->3	e->33	s->3	
nsatt	 ->2	.->2	
nsavg	ö->1	
nsavt	a->1	
nsbeg	r->3	
nsber	ä->1	
nsbes	t->6	
nsbev	i->2	
nsbol	a->1	
nsbri	s->1	
nsbut	i->1	
nsch 	f->1	o->1	s->1	
nsch.	E->1	
nsch?	F->1	
nsche	n->2	r->2	
nsdag	 ->1	.->1	:->1	e->1	s->1	
nsdeb	a->2	
nsdep	a->1	
nsdir	e->1	
nsdok	u->1	
nsdom	s->1	
nsdug	l->2	
nsdöm	t->1	
nse a	t->8	
nse d	e->2	
nse h	u->1	
nse m	e->4	
nse o	m->1	
nse v	a->3	i->1	
nse, 	i->1	
nse.E	n->1	
nse; 	j->1	
nseen	d->11	
nsekv	e->61	
nseme	l->3	
nsen 	(->2	-->2	2->1	a->14	b->4	d->4	e->1	f->6	g->2	h->3	i->19	k->3	l->1	m->9	n->1	o->9	p->3	r->1	s->20	t->8	u->4	v->3	ä->3	ö->1	
nsen,	 ->13	
nsen.	 ->2	A->2	D->11	F->1	H->3	I->1	J->2	L->1	M->1	N->1	O->3	R->2	S->1	T->1	V->7	
nsen?	F->1	
nsenN	ä->1	
nsenl	i->1	
nsens	 ->17	,->1	
nser 	4->1	a->116	b->1	d->18	e->4	f->15	h->2	i->9	j->33	k->6	l->1	n->2	o->16	p->1	r->2	s->9	u->4	v->20	ä->2	ö->1	
nser,	 ->6	
nser.	 ->1	(->1	9->1	A->1	H->1	I->1	J->1	O->1	V->2	
nser?	E->1	M->1	V->1	
nsera	 ->4	d->5	n->1	r->2	s->1	t->2	
nseri	n->1	
nsern	a->36	
nserv	a->7	
nses 	d->1	m->1	u->1	v->2	
nsett	 ->2	
nseur	o->1	
nsfor	u->1	
nsfri	a->1	h->2	
nsfrä	m->1	
nsfrå	g->5	
nsfun	k->1	
nsför	d->2	f->1	h->1	k->2	m->2	s->14	
nsgru	n->1	
nshau	s->1	
nshin	d->10	
nshäm	m->2	
nsibi	l->1	
nsidi	g->4	
nsiel	l->28	
nsier	a->16	i->34	
nsifi	e->3	
nsikt	.->1	e->4	
nsin 	h->3	k->1	m->1	o->1	p->1	s->1	t->2	ä->1	
nsin.	B->1	
nsind	u->1	
nsini	t->1	
nsinn	e->2	
nsinr	i->1	
nsins	a->1	
nsion	 ->6	,->1	.->5	e->13	s->1	ä->1	
nsisk	 ->1	t->1	
nsist	e->6	
nsite	t->1	
nsiti	o->1	v->1	
nsitl	a->2	ä->1	
nsitr	u->1	
nsitt	r->1	
nsiv 	k->1	s->1	t->1	
nsiva	 ->2	r->1	
nsivt	 ->6	
nsiär	e->1	
nsjov	i->17	
nsk T	V->1	
nsk b	a->1	
nsk d	a->1	
nsk k	v->1	
nsk l	a->1	ä->1	
nsk n	a->1	
nsk p	a->1	r->1	
nsk r	ä->1	
nsk s	t->1	
nska 	a->13	b->8	d->16	e->7	f->19	g->2	h->6	i->2	k->16	l->4	m->16	n->1	o->17	p->6	r->14	s->21	t->5	u->2	v->3	
nska,	 ->3	
nska.	D->1	E->2	P->1	V->2	
nskad	 ->5	e->8	
nskaf	f->1	
nskam	p->1	
nskan	 ->12	.->1	a->1	d->2	
nskap	 ->35	"->3	,->8	.->9	:->1	e->139	l->36	s->86	
nskar	 ->29	,->1	.->2	
nskas	 ->5	,->1	
nskat	 ->8	,->1	.->2	s->3	t->1	
nske 	I->1	a->2	b->3	d->4	f->4	g->1	h->2	i->10	k->6	l->5	m->2	n->3	o->5	r->2	s->2	t->3	v->5	ä->6	
nske,	 ->1	
nskem	å->3	
nskil	d->25	t->3	
nskli	g->43	
nskni	n->41	
nskom	m->16	n->3	
nskon	f->9	k->1	t->8	
nskos	t->2	
nskra	f->36	
nskri	t->3	v->2	
nskrä	m->1	n->11	
nskt 	b->1	f->1	k->1	s->1	u->1	v->1	
nskt.	(->1	
nskta	l->1	
nskul	t->6	
nskur	s->6	
nskvä	r->10	
nsla 	-->1	a->7	f->1	g->1	m->3	
nsla"	.->1	
nsla,	 ->1	
nslag	 ->13	e->9	n->7	s->1	
nsled	a->11	
nslen	,->1	.->1	
nsler	 ->1	
nsles	k->1	n->4	
nslie	r->1	
nslig	 ->12	a->7	t->2	
nslog	s->1	
nslol	a->1	
nslom	ä->1	
nslor	 ->4	.->1	
nslut	a->5	e->5	i->2	n->17	
nsläg	r->1	
nslå 	m->1	
nslåd	a->1	
nslår	 ->1	
nslås	 ->2	
nsmed	b->1	e->1	l->3	
nsmin	i->2	
nsmom	e->1	
nsmyn	d->8	
nsmäl	t->1	
nsmän	n->5	
nsmäs	s->1	
nsmål	 ->1	
nsmöt	e->1	
nsnac	k->2	
nsnin	g->19	
nsniv	å->2	
nsoli	d->3	
nsomr	å->3	
nsord	f->1	n->1	
nspak	e->1	
nspar	k->1	
nspek	t->12	
nspel	n->1	
nspir	e->3	
nspla	n->2	
nspol	i->79	
nspor	t->108	
nspri	d->1	n->4	s->1	
nspro	c->5	j->1	
nsprå	k->7	
nsrad	 ->1	
nsram	 ->1	
nsreg	e->3	l->9	
nsrel	a->1	
nsrol	l->1	
nsrät	t->43	
nssam	h->5	m->1	t->1	
nssch	e->1	
nssek	t->1	
nssit	u->1	
nsska	d->1	n->1	
nssky	d->2	
nsstr	a->1	ö->1	
nsstä	m->20	
nsstö	r->1	
nssvå	r->1	
nssys	t->6	
nst -	 ->1	
nst 1	0->1	2->1	
nst 3	 ->2	
nst 4	0->1	
nst a	r->1	
nst b	e->1	
nst d	ä->2	
nst f	r->1	
nst i	 ->2	n->1	
nst l	i->1	
nst m	i->1	å->1	
nst n	ö->1	
nst o	c->3	m->1	
nst p	e->1	å->1	
nst r	ö->1	
nst s	a->1	e->1	k->2	t->1	
nst u	n->1	t->1	
nst v	a->2	
nst å	t->1	
nst, 	d->1	e->1	h->1	
nst.J	a->2	
nsta 	g->2	m->1	s->1	v->1	
nstab	u->1	
nstag	a->2	
nstak	a->5	
nstal	l->1	t->1	
nstan	s->37	
nstat	 ->1	e->40	l->5	
nstee	n->5	
nstef	e->1	ö->5	
nstek	n->2	
nstel	e->1	
nstem	a->5	ä->34	
nsten	 ->2	,->2	e->1	
nstep	r->1	
nster	 ->42	"->1	,->8	.->13	n->9	r->3	s->1	
nstes	e->2	
nstfu	l->1	
nstgö	r->3	
nstig	a->1	t->2	
nstil	l->3	
nstin	k->2	r->1	
nstit	u->158	
nstjä	n->1	
nstma	r->1	
nston	e->27	
nstor	a->2	
nstra	 ->1	t->3	
nstre	a->8	r->3	s->2	t->1	
nstru	e->5	k->32	m->52	
nsträ	n->46	
nstrå	l->1	
nstsv	a->1	
nstäl	l->58	
nstäm	d->1	m->22	
nstän	d->5	
nståe	n->1	
nsult	a->2	b->1	e->2	
nsume	n->61	
nsumt	i->2	
nsund	e->3	
nsupp	f->1	
nsutb	y->3	
nsuts	ä->2	
nsvar	 ->69	,->23	.->27	?->1	a->10	e->57	i->54	s->70	
nsver	k->1	
nsvil	j->1	l->9	
nsvän	l->1	
nsvär	d->10	t->2	
nsyn 	g->1	i->1	o->4	t->65	v->1	ä->2	
nsyn,	 ->1	
nsyn.	A->1	S->2	
nsyn;	 ->1	
nsyne	n->4	
nsyns	t->2	
nsäga	r->1	
nsäke	r->3	
nsämn	e->1	
nsäre	n->2	
nsätt	 ->3	,->1	n->5	
nsåg 	a->7	d->2	e->1	o->1	s->1	
nsåte	r->1	
nsåtg	ä->1	
nsöka	 ->1	n->1	r->6	
nsökn	i->1	
nsökt	 ->1	
nsöve	r->12	
nsövn	i->1	
nt (t	.->1	
nt - 	e->1	f->1	i->1	o->1	s->1	t->1	v->1	
nt 19	9->2	
nt As	s->1	
nt Cl	i->1	
nt Eu	r->2	
nt al	l->5	
nt an	a->1	s->1	v->3	
nt ar	r->1	
nt at	t->16	
nt av	 ->54	
nt ba	k->1	r->1	
nt be	s->2	
nt bi	g->1	
nt bo	r->1	
nt br	i->1	
nt bu	d->1	
nt bö	r->2	
nt ce	n->1	
nt de	 ->1	b->2	n->2	t->1	
nt di	s->1	
nt ek	o->1	
nt el	l->3	
nt en	 ->2	b->1	
nt et	t->1	
nt ex	a->1	e->2	
nt fa	k->1	l->4	
nt fi	n->1	
nt fr	a->1	å->4	
nt fu	l->1	
nt fy	s->1	
nt fö	r->44	
nt ga	r->1	
nt ge	 ->2	n->2	
nt gr	u->1	
nt gä	l->2	
nt ha	 ->2	r->7	
nt he	l->1	
nt ho	p->1	
nt hu	r->1	s->1	
nt hå	l->1	
nt i 	P->1	d->5	e->1	f->4	h->1	p->1	s->2	v->2	
nt id	e->1	
nt if	r->1	
nt ig	e->1	
nt in	b->1	f->1	i->1	n->2	o->2	r->1	t->5	
nt ka	n->4	o->1	
nt ko	m->3	n->2	r->3	
nt kr	a->1	i->1	
nt ku	n->1	
nt kv	i->1	
nt kä	n->1	
nt le	d->1	
nt li	t->1	
nt lj	u->1	
nt lö	p->1	
nt ma	t->1	
nt me	d->6	n->1	r->1	
nt mi	g->1	
nt mo	t->2	
nt må	s->3	
nt mö	j->1	
nt nu	,->1	
nt ny	t->1	
nt nä	r->1	
nt nå	d->1	g->1	
nt oc	h->25	k->2	
nt om	 ->8	k->1	r->2	
nt pl	a->1	
nt pr	a->1	e->1	i->1	o->1	
nt pu	n->1	
nt på	 ->5	
nt re	g->1	p->1	
nt sa	k->1	m->1	
nt se	 ->1	d->1	r->1	t->2	x->1	
nt si	g->2	
nt sj	ä->2	
nt sk	a->2	u->2	
nt sl	a->1	
nt sn	a->1	
nt so	c->1	m->36	
nt st	a->1	r->1	ä->1	ö->2	
nt sv	å->1	
nt sy	n->1	s->1	
nt sä	t->12	
nt så	 ->2	
nt ta	n->1	r->1	
nt te	k->1	o->1	x->1	
nt ti	l->15	t->1	
nt tv	å->1	
nt un	d->6	
nt up	p->2	
nt ur	 ->1	
nt ut	 ->1	a->2	s->2	
nt va	r->2	
nt ve	t->1	
nt vä	n->1	
nt vå	l->1	
nt äm	n->1	
nt än	n->1	
nt är	 ->5	
nt åt	e->1	
nt ön	s->1	
nt öv	e->3	
nt!"J	a->1	
nt, L	a->1	
nt, S	o->1	
nt, a	t->1	v->1	
nt, b	e->1	
nt, d	e->3	v->1	ä->1	
nt, e	l->1	t->1	
nt, f	r->1	å->1	ö->1	
nt, g	e->1	
nt, h	a->1	e->1	
nt, i	 ->2	n->4	
nt, k	o->1	
nt, l	i->1	
nt, m	e->3	
nt, o	c->5	
nt, r	a->1	ä->1	
nt, s	ä->1	å->1	
nt, u	t->2	
nt, v	i->1	
nt-Ex	u->1	
nt. V	i->1	
nt.De	n->1	s->2	t->10	
nt.En	 ->1	
nt.Eu	r->1	
nt.Fr	a->1	
nt.Fö	r->3	
nt.He	r->3	
nt.I 	m->1	n->1	s->1	v->1	
nt.Ja	,->1	g->5	
nt.Lå	t->1	
nt.Ma	x->1	
nt.Me	d->1	n->1	
nt.Nä	r->1	
nt.OK	,->1	
nt.Pl	ä->1	
nt.Sa	m->1	n->1	
nt.Så	 ->2	
nt.Vi	 ->3	
nt: U	n->1	
nt: v	i->1	
nta -	 ->1	
nta 1	0->1	
nta M	a->1	
nta N	a->1	
nta S	h->1	t->1	
nta a	n->1	r->1	v->2	
nta b	e->2	i->4	
nta d	e->5	
nta e	l->2	n->6	t->4	
nta f	o->21	r->2	ö->2	
nta h	å->1	
nta i	 ->4	
nta k	o->2	r->1	v->1	
nta l	a->1	
nta m	a->1	e->1	o->1	y->2	ö->1	
nta n	a->10	å->1	
nta o	l->1	s->1	
nta p	r->1	å->4	
nta r	e->1	å->1	
nta s	a->1	i->1	t->18	
nta t	i->3	y->1	
nta u	t->1	
nta ä	n->2	
nta å	t->1	
nta, 	r->1	
nta. 	V->1	
nta.D	e->1	
ntabl	a->1	
ntabr	i->3	
ntade	s->1	
ntag 	a->2	f->2	g->1	i->3	o->1	t->1	v->1	ä->1	
ntag,	 ->4	
ntag.	I->1	O->1	
ntag?	F->1	
ntaga	n->14	r->3	
ntage	n->3	t->3	
ntagi	t->22	
ntagl	i->1	
ntagn	a->4	
ntags	b->1	f->3	m->1	r->3	t->2	
ntain	e->1	
ntakt	 ->4	.->1	e->12	
ntal 	a->4	b->2	f->6	i->1	k->4	l->2	m->5	n->1	p->2	r->4	s->6	å->1	ö->3	
ntal,	 ->1	
ntala	 ->4	
ntale	t->19	
ntali	t->1	
ntals	 ->11	
ntami	n->2	
ntan 	p->4	
ntan.	J->1	
ntan?	Ä->1	
ntana	 ->1	
ntand	e->2	
ntans	v->6	
ntant	 ->2	e->11	
ntar 	a->2	b->3	d->2	e->2	f->3	i->1	j->3	k->2	m->11	n->1	o->4	p->6	s->10	v->4	ä->1	
ntar,	 ->1	
ntar.	D->1	
ntare	r->21	
ntari	k->9	s->18	t->3	u->1	
ntas 	a->2	f->2	g->2	k->1	m->1	n->1	p->1	r->1	s->2	
ntas,	 ->2	
ntas.	O->1	
ntasi	f->1	n->1	
ntast	i->9	
ntat 	i->2	l->1	m->2	o->1	p->1	s->1	
ntat.	T->1	
ntate	t->1	
ntati	o->13	v->5	
ntav 	ö->1	
nte -	 ->3	
nte 1	9->1	
nte B	e->1	
nte E	U->2	u->1	
nte a	c->9	k->1	l->31	n->15	r->1	s->1	t->59	u->4	v->17	
nte b	a->91	e->27	i->1	l->13	o->3	r->2	ö->4	
nte c	h->1	
nte d	e->48	i->2	r->2	ä->2	ö->2	
nte e	f->1	l->2	n->40	r->1	t->12	x->3	
nte f	a->10	i->17	o->9	r->8	u->6	ä->1	å->17	ö->55	
nte g	a->4	e->16	j->3	l->10	o->9	ä->4	å->13	ö->15	
nte h	a->98	e->49	i->2	u->3	ä->5	å->3	ö->6	
nte i	 ->25	f->2	g->1	l->1	n->17	s->1	
nte j	u->1	
nte k	a->55	l->2	o->29	r->1	u->13	ä->1	ö->1	
nte l	a->1	e->6	i->3	u->1	y->6	ä->38	å->8	ö->2	
nte m	e->26	i->18	o->3	y->5	å->4	ö->6	
nte n	e->1	i->2	o->2	u->2	ä->5	å->26	ö->11	
nte o	b->1	c->3	f->1	l->1	m->22	p->2	r->2	
nte p	a->2	l->2	o->1	r->4	å->37	
nte r	a->3	e->11	i->1	u->1	ä->12	å->5	ö->2	
nte s	a->6	e->8	j->3	k->45	l->2	n->3	o->4	p->2	t->7	v->3	y->1	ä->10	å->10	
nte t	a->23	i->32	j->1	r->4	u->3	v->2	y->1	ä->6	
nte u	n->7	p->23	r->1	t->19	
nte v	a->29	e->3	i->9	o->2	ä->5	å->2	
nte ä	g->1	n->9	r->74	v->1	
nte å	l->1	s->1	t->4	
nte ö	k->2	n->2	p->1	v->7	
nte!D	e->1	
nte!M	e->1	
nte, 	a->3	e->1	h->2	i->1	m->1	o->3	v->2	ä->2	
nte.A	n->1	
nte.B	e->1	
nte.D	e->2	ä->1	
nte.H	e->2	
nte.J	a->2	
nte.S	å->1	
nte.V	i->2	
nte.Å	 ->1	r->1	
nte: 	v->1	
nte?F	ö->1	
nte?H	ä->1	
ntegr	a->16	e->23	i->3	
ntekn	i->3	
ntell	e->3	i->5	t->1	
ntels	e->5	
ntemo	t->27	
nten 	I->1	S->1	a->1	e->1	f->4	h->1	i->9	k->2	n->2	o->5	u->1	v->1	ä->1	
nten"	.->1	
nten)	 ->1	
nten,	 ->6	
nten.	D->2	E->1	H->1	V->1	Å->1	
nten?	J->1	
ntens	 ->4	i->12	
ntent	i->1	
nter 	a->1	f->5	h->2	i->5	k->1	m->1	o->5	s->2	t->1	
nter,	 ->2	
nter-	k->1	
nter.	D->2	E->1	I->1	J->1	V->2	
ntera	 ->74	,->1	.->1	d->8	n->2	r->19	s->15	t->8	
nteri	m->8	n->40	
ntern	 ->5	a->118	e->11	t->4	
nterp	a->1	
nterv	e->7	j->3	
ntes.	F->1	
ntet 	-->4	1->2	M->1	a->26	b->13	c->1	d->10	e->4	f->26	g->11	h->25	i->30	j->3	k->16	l->5	m->10	n->5	o->44	p->3	r->5	s->33	t->7	u->4	v->10	ä->9	å->1	
ntet,	 ->37	
ntet-	 ->1	
ntet.	B->1	D->13	F->1	H->1	J->4	K->1	L->1	M->2	P->1	S->1	V->3	
ntet:	 ->1	
ntet?	D->1	
ntets	 ->103	
ntext	e->1	
ntfrå	g->6	
nti -	 ->1	
nti f	ö->5	
nti h	a->2	
nti i	 ->3	g->1	
nti k	o->1	
nti o	c->2	m->1	
nti p	å->1	
nti s	å->1	
nti v	a->1	
nti! 	J->2	U->1	
nti, 	d->1	m->1	ä->1	
nti-g	e->1	
nti-i	r->1	
nti-r	a->1	
nti.H	ä->1	
nti.J	a->1	
nti.V	i->1	
ntial	 ->1	,->1	.->1	
ntibe	d->1	
ntide	m->1	
ntiel	l->8	
ntier	 ->10	a->1	i->4	n->5	
ntieu	r->1	
ntifa	s->3	
ntifi	e->14	q->1	
ntifo	l->1	n->2	
ntika	 ->1	
ntiko	l->1	
ntikr	y->2	
ntil 	n->1	
ntile	r->1	
ntili	s->1	
ntime	t->1	
ntimt	 ->1	
ntimö	g->1	
ntin 	a->1	f->1	m->1	
ntine	n->5	
nting	 ->57	,->3	.->2	e->10	
ntins	 ->1	
ntinu	e->2	
ntion	 ->4	,->1	e->34	i->1	s->1	
ntiqu	e->1	
ntise	k->2	m->3	
ntisk	 ->2	a->4	
ntisy	s->1	
ntita	t->4	
ntite	t->8	
ntitr	u->1	
ntkat	e->1	
ntkus	t->1	
ntlig	 ->33	,->1	.->1	a->76	e->57	g->17	h->29	t->35	
ntnin	g->8	
ntog 	b->1	d->1	e->3	k->3	l->4	o->1	p->1	r->2	
ntogs	 ->8	,->2	
ntole	r->4	
ntom 	i->1	
ntons	 ->1	
ntor 	e->1	f->2	h->1	o->1	
ntor,	 ->2	
ntore	n->1	t->1	
ntorg	a->1	
ntpol	i->2	
ntpra	t->1	
ntra 	f->1	h->1	i->1	k->2	o->1	p->1	s->2	t->1	u->1	v->1	
ntra,	 ->1	
ntrad	 ->1	
ntrak	t->4	
ntral	 ->7	-->6	.->2	a->20	b->8	e->2	f->1	i->24	t->6	
ntran	 ->1	d->2	
ntrap	r->1	
ntrar	 ->8	
ntras	 ->3	t->2	
ntrat	 ->1	i->16	
ntrea	l->2	
ntrel	a->1	
ntrep	r->5	
ntrer	a->15	
ntres	s->120	
ntret	 ->1	
ntrod	u->6	
ntrol	,->1	.->1	l->178	
ntrov	e->4	
ntrum	 ->5	!->1	,->2	e->1	
ntryc	k->15	
nträd	e->36	
nträf	f->26	
nträt	t->1	
ntrån	g->1	
nts a	n->1	v->5	
nts b	u->1	
nts e	n->1	
nts f	ö->1	
nts h	a->1	
nts i	 ->1	n->2	
nts m	e->2	å->1	
nts o	r->1	
nts p	å->1	
nts t	i->1	
nts v	a->1	
nts ä	r->1	
nts, 	a->1	ä->1	
nts.D	e->1	
nts.J	a->1	
ntsat	s->1	
ntsbe	s->1	
ntsfo	r->1	
ntsif	f->1	
ntska	n->1	
ntsko	l->1	
ntsky	d->5	
ntsle	d->28	
ntsut	s->2	
nttil	l->1	
ntuel	l->21	
ntunn	e->1	
nture	r->1	
ntusi	a->3	
ntvar	o->1	
ntver	k->2	
ntvän	l->1	
ntydd	e->2	
ntydi	g->4	
ntyg 	o->1	
ntyga	 ->3	
ntyra	 ->3	r->5	s->1	
ntäkt	s->5	
ntära	 ->2	
ntóni	o->1	
ntöre	n->1	r->1	
ntörs	o->1	
nu - 	a->1	
nu 34	 ->1	
nu Er	i->1	
nu al	l->1	
nu an	s->1	
nu at	t->5	
nu av	 ->1	
nu be	f->1	h->2	t->1	
nu bl	i->3	o->1	
nu de	f->1	s->1	t->2	
nu di	s->2	
nu dö	p->1	
nu ef	t->1	
nu eg	e->1	
nu en	 ->12	
nu et	t->8	
nu eu	r->1	
nu fa	k->1	t->1	
nu fi	n->3	
nu fl	e->1	
nu fr	a->1	å->1	
nu få	r->1	t->2	
nu fö	r->10	
nu ge	m->1	n->1	r->2	t->1	
nu gä	l->3	
nu gå	 ->3	
nu gö	r->3	
nu ha	r->13	
nu hå	l->1	r->2	
nu hö	g->4	r->1	
nu i 	p->1	s->1	v->1	
nu ig	e->1	
nu in	n->3	t->35	
nu ka	n->5	
nu ko	m->5	n->1	
nu li	g->1	
nu ly	s->1	
nu lä	g->1	s->1	t->1	
nu me	d->1	r->7	
nu mi	n->1	
nu mä	r->1	
nu må	s->8	
nu nu	m->1	
nu nä	r->8	
nu nå	t->1	
nu oc	h->3	k->1	
nu of	f->1	t->1	
nu om	s->1	
nu pl	a->1	
nu pr	i->1	ö->1	
nu på	 ->1	.->1	g->2	
nu ru	l->1	
nu rå	d->2	
nu rö	s->1	
nu se	r->1	s->1	
nu si	f->1	
nu sk	a->4	e->1	u->1	ö->1	
nu sl	å->1	
nu sm	i->1	
nu so	m->1	
nu sp	e->1	
nu st	a->1	r->1	ä->1	å->3	ö->5	
nu sv	å->1	
nu sä	g->1	t->1	
nu så	 ->2	
nu ta	g->2	l->1	r->2	
nu ti	l->3	
nu ty	d->2	v->1	
nu un	d->1	
nu up	p->3	
nu va	d->1	
nu ve	m->1	r->1	
nu vi	d->2	k->2	l->1	s->1	
nu äl	d->1	
nu än	 ->1	t->5	
nu är	 ->9	,->1	
nu åt	e->1	
nu, e	f->1	
nu, i	 ->1	
nu, m	e->2	
nu, u	n->1	
nu, ö	v->1	
nu..T	a->1	
nu.De	t->1	
nu.Ja	g->1	
nu.Ko	m->1	n->1	
nu.Lå	t->1	
nu.Vi	 ->2	
nu: g	ö->1	
nu; i	 ->1	
nu?Ja	g->1	
nuari	 ->12	,->3	.->1	
nuc s	e->1	
nuerl	i->2	
nuft 	g->1	
nuft.	V->1	
nufte	t->1	
nufti	g->11	
nulli	t->1	
nuläg	e->1	
num f	r->1	
num h	a->1	
num i	 ->1	
num ä	n->1	
num.D	e->1	
numer	a->5	
numme	r->2	
nunno	r->1	
nuppr	o->4	
nus 2	0->1	
nus f	y->1	
nus t	j->1	
nusdi	m->1	
nusgr	a->2	
nussl	a->1	
nut f	ö->2	
nut n	ä->1	
nut.(	P->1	
nut.)	F->1	
nut.J	a->1	
nuten	 ->3	
nuter	 ->3	,->1	.->6	
nutet	 ->1	
nutna	 ->2	
nutpu	n->1	
nuts-	b->1	
nutta	 ->2	
nutve	c->1	
nuvar	a->45	
nvald	.->1	
nvand	r->18	
nvape	n->12	
nvara	n->4	
nvaro	 ->2	,->1	n->1	
nveck	l->2	
nvent	 ->1	a->1	i->23	
nverg	e->5	
nverk	a->7	
nvers	,->1	
nvest	e->15	
nvete	t->1	
nvikt	 ->3	e->2	
nvink	e->11	l->1	
nvisa	 ->9	d->6	r->7	s->4	t->1	
nvish	e->3	
nvisn	i->10	
nvist	 ->1	
nvit 	f->1	
nvolv	e->9	
nväg 	e->6	k->1	o->1	
nväg,	 ->1	
nväg.	A->1	M->1	
nväga	r->9	
nvägs	n->2	o->1	
nvänd	 ->1	a->64	b->9	e->31	n->62	s->20	
nvänt	 ->5	a->2	s->5	
nvärd	a->1	
nvåna	r->9	
ny bi	l->1	
ny eu	r->1	
ny fa	s->1	
ny fo	r->1	
ny fö	r->2	
ny gr	a->1	
ny hä	r->1	
ny in	f->1	s->1	
ny ke	m->1	
ny ko	m->3	
ny ku	l->3	
ny kv	a->1	
ny la	g->1	
ny le	d->1	
ny li	v->1	
ny my	n->1	
ny oc	h->1	
ny ol	j->1	
ny pe	r->2	
ny rö	s->2	
ny se	k->1	
ny si	t->1	
ny sp	e->1	
ny st	o->1	
ny sy	n->1	s->1	
ny ty	p->1	
ny up	p->1	
ny ve	t->1	
ny vi	g->1	t->1	
nya "	l->1	
nya 8	1->1	
nya E	U->1	u->2	
nya a	r->9	t->1	v->2	
nya b	e->6	i->6	u->1	y->1	
nya d	e->2	i->2	o->1	
nya e	u->1	x->1	
nya f	e->1	r->3	ö->6	
nya g	e->2	r->1	
nya i	m->1	n->3	
nya j	o->1	
nya k	l->1	o->16	
nya l	a->1	e->1	i->1	ä->4	
nya m	a->1	e->8	i->1	o->1	y->2	å->1	ö->3	
nya n	o->1	ä->1	
nya o	b->1	c->2	m->2	r->1	
nya p	a->1	e->3	r->9	
nya r	a->1	e->10	i->2	u->1	ä->2	
nya s	i->1	p->1	y->4	ä->1	
nya t	e->4	i->1	j->2	y->1	
nya u	p->1	t->2	
nya v	e->2	i->1	å->1	
nya ä	n->2	
nya å	r->1	t->5	
nya, 	u->1	
nya; 	k->1	
nyand	e->1	
nyans	e->1	t->2	
nyar 	l->1	
nyas 	o->1	
nyast	e->1	
nybar	 ->4	,->1	a->34	
nybil	s->2	
nycke	l->8	
nydan	a->1	
nye o	r->1	
nyels	e->6	
nyeta	b->1	
nyfas	c->1	
nyför	v->1	
nyhet	 ->1	.->2	e->9	s->1	
nykte	r->2	
nyktr	a->1	
nylib	e->1	
nylig	e->29	
nym m	e->1	
nym s	o->1	
nym.D	e->1	
nyma 	B->1	
nymit	e->1	
nynaz	i->6	
nyo s	k->1	
nyon 	1->1	s->1	
nyon,	 ->1	
nypla	n->1	
nyska	p->1	
nyss 	a->1	b->1	e->1	g->1	n->1	o->3	s->2	
nyss,	 ->2	
nyss.	S->1	
nyta 	a->1	b->1	d->1	m->1	s->1	
nyter	 ->2	
nytni	n->1	
nyts 	t->1	
nytt 	a->1	b->2	e->1	f->3	g->1	i->3	k->2	l->1	m->2	o->2	p->5	s->11	t->1	u->1	v->1	å->2	ö->1	
nytt,	 ->3	
nytt.	D->2	J->1	
nytta	 ->14	,->1	.->4	n->1	
nytti	g->13	
nyttj	a->41	
nytto	-->1	a->1	
nyval	d->1	
nyårs	a->1	
nz Fi	s->3	
nz Fl	o->2	
nz be	t->1	
nz et	t->1	
nz fr	å->1	
nz fö	r->1	
nz oc	h->5	k->1	
nz om	 ->1	
nz to	g->1	
nz)(T	a->1	
nz).H	e->1	
nz, L	a->3	
nzFru	 ->1	
nzbet	ä->1	
nzes-	C->1	
nzále	z->1	
nÄrad	e->1	
näcka	 ->1	s->1	
näer;	 ->1	
nägna	 ->1	
nälla	 ->1	
nälle	t->1	
nämli	g->43	
nämna	 ->24	,->1	n->1	r->2	s->2	
nämnd	a->8	e->18	
nämne	r->5	
nämni	n->3	
nämns	 ->8	.->1	
nämnt	 ->9	,->2	.->2	s->6	
nämnv	ä->1	
nämt 	a->1	
när -	 ->2	
när A	n->1	
när B	a->8	o->1	
när C	E->1	
när E	u->1	
när K	i->5	
när M	a->1	o->13	
när N	i->1	
när P	a->17	r->1	
när R	e->2	
när S	c->1	o->1	
när V	i->4	
när W	a->1	
när a	l->7	n->1	t->1	
när b	e->2	l->1	
när c	o->1	
när d	e->197	i->1	o->1	
när e	n->7	x->1	
när f	ä->1	ö->6	
när g	e->1	i->1	
när h	a->13	
när i	 ->1	
när j	a->14	
när k	a->1	o->6	
när l	o->1	
när m	a->19	e->2	i->1	ä->1	
när n	a->1	i->5	y->1	å->3	
när o	c->1	
när p	e->1	
när r	e->3	
när s	o->3	
när t	i->1	
när v	e->2	i->40	ä->1	
när ä	r->1	v->1	
när ö	v->2	
när! 	1->1	B->1	C->1	D->2	E->3	F->1	I->2	J->6	L->2	N->2	O->1	T->1	U->1	V->4	Ä->1	
när!.	H->1	
när!E	r->1	
när!J	a->1	
när, 	a->8	b->3	d->1	f->5	h->5	j->3	k->13	l->1	m->8	n->2	o->2	p->1	r->1	s->4	t->1	u->1	v->6	ä->10	
när. 	N->1	
när.D	e->2	
när.G	e->1	
när.J	a->6	
när.V	i->1	
nära 	5->1	a->1	b->1	d->1	f->9	h->1	k->1	m->2	o->1	p->1	r->1	s->7	
nära,	 ->1	
nären	 ->37	,->4	.->2	s->3	
närer	 ->9	!->1	n->10	
närfr	å->1	
närhe	t->5	
närin	g->12	
närma	 ->2	n->1	r->20	s->13	
närme	l->1	
närmn	i->5	
närpe	r->1	
närs 	h->1	
närsy	n->1	
närva	r->46	
näsdu	k->1	
nästa	 ->29	.->1	n->17	
nät k	a->1	
nät o	c->1	s->1	
nät s	k->1	o->1	
nät. 	D->1	
näten	 ->2	
nätet	 ->2	
nätst	r->1	
nätte	r->1	
nätve	r->11	
nävar	e->1	
nå an	s->1	
nå da	g->1	
nå de	 ->3	n->2	s->2	t->5	
nå ek	o->2	
nå en	 ->17	h->2	i->1	
nå et	t->6	
nå fa	s->1	
nå fr	a->5	
nå ge	m->1	
nå hö	g->1	
nå me	d->2	
nå må	l->1	
nå nå	g->1	
nå på	 ->2	
nå re	s->1	
nå si	n->1	
nå vå	r->5	
nå yt	t->1	
nå än	d->1	
nå åt	e->1	
nå ön	s->1	
nå, n	ä->1	
nå. D	e->1	
nå.Fr	u->1	
nå.Ja	g->1	
nå.Sl	u->1	
nåbar	 ->2	
nåd a	t->1	
nåda 	d->1	
nådda	 ->3	
nådde	 ->2	s->1	
någon	 ->110	,->2	.->1	s->14	t->38	
någor	l->1	
något	 ->183	,->2	.->6	?->1	
några	 ->147	
nåla 	b->1	f->1	
nåla,	 ->1	
nålar	e->2	
når d	e->4	i->1	
når e	n->4	t->1	
når m	o->1	y->1	å->1	
når s	a->1	
når v	i->1	
nårig	a->1	
nårin	g->1	
nås b	ä->1	
nås e	n->1	
nås g	e->1	
nås i	 ->1	n->1	
nås.F	ö->1	
nås.L	a->1	
nått 	e->3	g->1	k->1	m->1	n->2	s->2	u->2	v->1	
nått,	 ->1	
nått.	P->1	
nåtts	 ->3	.->2	
nçois	 ->1	
nève 	1->1	
nève,	 ->1	
nèvek	o->1	
nödbe	d->1	
nöden	s->1	
nödig	 ->2	.->1	a->3	t->6	
nödin	s->1	
nödsi	t->1	
nödvä	n->124	
nöja 	m->1	o->5	s->2	
nöjak	t->2	
nöjd 	m->1	p->1	
nöjda	 ->6	,->3	
nöje 	B->1	E->1	f->1	o->1	
nöjer	 ->1	
nöjet	 ->2	
nöjt 	o->1	
nör t	a->1	
nör, 	B->1	
nörsk	a->2	
nöste	r->19	
nöt.D	e->1	
nötkö	t->3	
nötsk	a->1	
nötte	r->1	
növad	e->1	
növit	t->1	
növra	r->1	
o (KO	M->2	
o - d	e->1	
o - e	n->1	
o - t	i->1	
o 199	8->1	
o Cad	i->5	
o Eur	o->1	
o Leo	n->1	
o Pro	d->2	
o Roj	o->1	
o Sán	c->1	
o Tom	é->2	
o Tra	n->1	
o Val	l->3	
o Vit	o->1	
o acc	e->1	
o ang	a->1	
o att	 ->8	
o bea	k->1	
o bes	l->2	
o bla	n->1	
o bär	 ->1	
o det	.->1	
o dis	k->1	
o då,	 ->1	
o ett	 ->1	
o far	 ->1	
o fat	t->1	
o fra	m->1	
o frå	n->1	
o ful	l->1	
o för	 ->15	b->1	e->2	s->1	
o god	t->1	
o gra	d->2	
o gån	g->3	
o har	 ->4	
o hår	d->1	
o i a	l->1	
o i d	e->1	
o i e	k->1	t->1	
o i f	r->3	
o i h	a->1	
o i l	a->1	
o i m	a->1	
o i n	å->1	
o int	e->1	
o kan	 ->2	
o kom	m->1	
o kva	r->1	
o käm	p->1	
o led	a->1	
o län	d->1	
o med	 ->1	
o mel	l->1	
o mil	j->6	
o min	u->1	
o mål	a->1	
o mån	a->2	
o mås	t->1	
o när	 ->2	
o någ	o->3	
o och	 ->16	
o ock	s->2	
o om 	l->1	s->1	u->1	
o per	 ->2	
o pun	k->1	
o på 	d->1	g->1	k->2	
o påp	e->1	
o res	p->1	
o sad	e->1	
o saf	e->1	
o sin	e->1	
o ski	s->1	
o sku	l->1	
o som	 ->14	,->1	
o så 	m->1	r->1	
o til	l->5	
o tim	m->1	
o tre	,->1	
o und	e->2	
o uta	n->1	
o utt	a->1	
o var	 ->1	a->1	
o vik	t->1	
o vil	j->1	
o väl	k->1	
o änd	r->1	
o är 	b->1	d->1	e->2	g->1	o->2	
o äve	n->2	
o år 	f->1	i->1	n->1	s->1	
o år,	 ->1	
o åre	n->2	
o års	 ->1	
o åte	r->1	
o öpp	e->1	
o öve	r->1	
o!All	t->1	
o, As	i->1	
o, He	l->1	
o, Ta	n->1	
o, Wy	e->1	
o, an	s->1	
o, at	t->1	
o, de	n->1	t->3	
o, dä	r->1	
o, el	l->1	
o, et	t->2	
o, fö	r->2	
o, he	l->1	
o, hu	v->1	
o, i 	d->1	e->1	
o, ko	m->1	
o, me	d->1	n->1	
o, mo	t->1	
o, oc	h->5	
o, or	d->1	
o, sa	m->1	
o, se	r->1	
o, so	m->6	
o, st	i->1	
o, sy	r->1	
o, ti	l->2	
o, vi	l->2	
o, än	d->1	
o- oc	h->1	
o-Pla	t->4	
o-aff	ä->1	
o-ana	l->1	
o-pro	t->1	
o-råd	e->1	
o. De	n->1	
o.- (	P->1	
o.Att	 ->1	
o.Avs	l->1	
o.Bet	ä->1	
o.Des	s->1	
o.Det	 ->2	t->2	
o.Där	a->1	
o.Eur	o->1	
o.Fle	r->1	
o.För	 ->1	s->2	
o.Her	r->2	
o.Hur	 ->1	
o.Jag	 ->5	
o.Kna	p->1	
o.Kom	m->1	
o.Låt	 ->1	
o.Men	 ->1	
o.När	 ->2	
o.Och	 ->1	
o.Om 	d->1	j->1	
o.Ord	e->1	
o.Sed	a->1	
o.Tro	t->1	
o.Ty 	e->1	
o.Vi 	b->1	m->3	ä->1	
o.m. 	a->2	d->1	i->1	ä->2	
o.m.,	 ->1	
o/Oil	-->1	
o: vi	 ->1	
o; de	t->1	
o? De	n->1	
o?Hur	 ->1	
oNäst	a->1	
oU, n	ä->1	
oU-ra	m->1	
oa fö	r->1	
oa os	s->1	
oa si	g->1	
oacce	p->31	
oad ö	v->3	
oade 	a->1	s->1	
oaklu	k->1	
oakta	t->1	
oakti	o->1	v->12	
oalit	i->14	
oanal	y->1	
oande	 ->7	.->2	
oanst	a->1	
oansv	a->5	
oanvä	n->1	
oar e	l->1	
oar k	o->1	
oar o	s->1	
oar s	i->2	
oard,	 ->1	
oares	,->1	
oater	 ->1	
oavbr	u->2	
oavse	t->8	
oavsi	k->2	
ob Sö	d->2	
obak,	 ->1	
obaks	o->1	
obal 	n->1	
obala	 ->4	n->6	
obali	s->5	
obalt	 ->1	,->1	
obase	n->1	
obb e	f->1	
obb o	c->1	
obb, 	s->1	v->1	
obby,	 ->1	
obbya	r->1	
obbyb	i->1	
obbyg	r->2	
obbyi	s->2	
obbym	a->1	
obbyn	 ->3	
obbyv	e->1	
obebo	e->1	
obefo	g->1	
obegr	i->3	ä->2	
obeha	g->2	
ober 	1->6	f->1	m->1	
obero	e->50	
obert	 ->1	
oberä	t->1	
obest	r->1	ä->1	
obesv	a->3	
obetä	n->1	
obili	s->7	
obin,	 ->1	
objek	t->1	
oblem	 ->71	,->13	.->22	:->1	;->2	?->1	a->5	e->65	o->3	
obles	 ->1	
oblig	a->14	
oboda	 ->2	s->1	
obser	v->2	
oc-di	r->1	
oc-tr	a->1	
oca C	o->1	
ocedu	r->1	
ocent	 ->75	,->2	.->10	a->2	s->5	
ocess	 ->22	"->1	,->2	.->13	?->1	e->66	r->3	u->1	
och "	U->1	s->1	t->1	
och (	A->1	
och -	 ->3	o->3	
och 0	 ->1	
och 1	-->1	0->2	3->1	4->1	6->1	7->2	9->13	
och 2	 ->1	,->1	.->1	0->3	1->3	2->1	5->1	7->1	9->1	
och 3	.->1	0->2	3->1	4->1	5->1	:->1	
och 4	.->1	1->2	5->4	7->1	8->2	
och 5	 ->1	.->1	3->1	
och 6	0->1	8->1	
och 7	 ->4	,->2	
och 8	 ->1	,->1	2->6	6->2	9->1	
och 9	 ->2	2->1	4->1	
och A	l->2	m->1	n->1	
och B	P->1	a->1	e->1	r->2	u->1	
och C	.->1	E->1	a->1	y->1	
och D	a->2	e->2	
och E	L->2	U->4	d->1	l->2	m->1	r->1	t->1	u->23	
och F	N->1	P->1	i->2	r->11	
och G	a->2	e->1	o->1	r->3	
och H	e->1	i->1	u->1	
och I	I->2	n->4	r->2	s->5	t->1	
och J	a->1	ö->1	
och K	a->1	i->6	o->1	u->1	
och L	a->3	e->5	
och M	A->1	a->3	e->1	
och N	o->1	y->1	
och O	L->1	n->1	
och P	P->1	S->2	a->9	o->2	r->1	
och R	a->3	
och S	a->10	c->1	j->1	o->1	p->1	t->2	w->1	y->8	
och T	a->4	s->1	u->1	y->2	
och U	z->1	
och V	i->1	ä->1	
och W	y->1	
och X	 ->1	
och a	c->1	d->2	g->2	k->4	l->18	m->4	n->58	r->15	s->4	t->150	v->32	
och b	a->13	e->52	i->10	l->8	o->5	r->15	u->3	y->2	ä->4	å->1	ö->6	
och c	a->2	e->6	h->2	
och d	a->3	e->449	i->11	j->4	o->9	r->3	u->1	y->1	ä->83	å->23	ö->1	
och e	f->33	g->1	j->1	k->22	l->1	n->90	r->16	t->33	u->9	x->4	
och f	a->14	e->3	i->12	l->10	o->7	r->83	u->9	y->2	ä->1	å->12	ö->167	
och g	a->7	e->43	i->3	j->1	l->3	o->2	r->10	ä->1	å->4	ö->17	
och h	a->44	e->54	i->1	j->4	o->11	u->15	y->2	ä->8	å->16	ö->6	
och i	 ->72	b->3	c->2	d->5	f->1	k->1	l->1	m->2	n->141	r->1	s->2	
och j	a->139	o->5	u->7	ä->1	
och k	a->21	i->1	l->4	n->1	o->128	r->18	u->7	v->10	ä->6	ö->1	
och l	a->17	e->16	i->11	j->1	o->9	u->1	y->3	ä->14	å->19	ö->2	
och m	a->21	e->142	i->39	o->24	u->1	y->8	ä->12	å->22	ö->9	
och n	a->11	e->8	i->8	o->5	u->9	y->13	ä->14	å->5	ö->6	
och o	a->4	b->2	c->8	d->1	e->2	f->6	j->1	k->4	l->8	m->39	n->1	p->2	r->8	s->5	t->1	u->3	
och p	a->25	e->9	l->3	o->17	r->32	å->29	
och r	a->7	e->66	i->9	o->4	u->1	ä->61	å->39	ö->1	
och s	a->43	e->29	i->10	j->6	k->29	l->21	m->2	n->4	o->131	p->9	t->61	u->5	v->12	y->16	ä->33	å->27	ö->2	
och t	.->1	a->20	e->6	h->1	i->59	j->4	o->6	r->18	u->17	v->3	y->14	ä->3	
och u	n->25	p->24	t->57	
och v	a->49	e->22	i->120	ä->26	å->11	ö->1	
och y	n->1	r->1	t->5	
och Ö	V->1	s->6	
och ä	g->2	n->12	r->10	v->30	
och å	 ->4	k->1	s->3	t->29	
och ö	k->3	m->1	n->1	p->13	r->1	s->4	v->20	
och)D	e->1	
och, 	d->1	f->3	h->1	i->1	n->1	r->1	s->4	t->1	u->1	
och.J	a->1	
och/e	l->1	
ochI 	o->1	
ochII	.->1	
ochis	t->1	
ochs 	i->1	
ocial	 ->30	-->1	a->78	d->15	f->26	i->34	p->4	t->18	
ocier	i->1	
ociet	y->1	
ocilo	v->1	
ocioe	k->3	
ock a	l->1	t->10	v->1	
ock d	e->3	
ock e	f->1	j->1	n->1	
ock f	r->3	å->1	ö->2	
ock g	a->1	r->1	
ock h	a->2	u->1	
ock i	 ->1	n->7	
ock k	a->2	l->1	o->3	
ock l	ä->2	
ock m	y->2	å->1	
ock n	u->1	y->1	å->1	
ock o	c->3	
ock p	a->1	
ock s	k->2	t->2	v->1	ä->2	
ock t	i->1	v->1	ä->1	
ock u	t->1	
ock v	i->5	ä->1	
ock ä	n->1	
ock å	t->2	
ock" 	-->1	
ock, 	R->1	i->2	m->1	s->3	t->1	
ock. 	M->1	
ock.J	a->1	
ock.K	i->1	
ocka 	f->2	t->1	
ockad	 ->1	.->1	i->1	
ockan	 ->1	.->1	
ockar	 ->1	
ockbi	l->1	
ocker	a->3	i->1	
ocket	.->1	
ockho	l->3	
ocks 	d->1	p->1	r->1	
ocksk	ö->1	
också	 ->570	,->10	.->5	
ockup	a->2	e->3	
oco, 	e->1	
od ad	m->1	
od an	l->1	
od at	t->3	
od av	 ->3	.->1	
od bi	l->1	
od bö	r->1	
od de	t->3	
od dä	r->1	
od ef	t->2	
od en	b->1	
od fa	m->1	
od fi	c->1	n->1	
od fr	å->1	
od få	r->1	
od fö	r->14	
od ha	r->1	
od i 	f->1	j->1	k->1	m->1	s->1	
od id	é->2	
od in	s->1	t->1	
od ja	g->1	
od jo	r->1	
od ko	m->2	
od le	d->1	
od me	d->3	
od mi	n->1	
od my	c->1	
od ny	l->1	
od om	 ->2	
od pr	o->1	
od på	 ->3	
od re	s->1	
od rö	s->1	
od sk	r->1	
od so	m->8	
od ta	r->1	
od ti	d->5	
od tr	o->1	
od tä	c->1	
od up	p->1	
od vi	 ->1	l->1	
od är	 ->4	
od åt	e->1	
od, e	n->1	
od, f	a->1	
od, m	e->1	
od, n	ä->1	
od, v	i->1	
od.De	 ->1	
od.Fa	k->1	
od.Vi	 ->1	
od?- 	(->1	
oda a	n->1	r->1	v->2	
oda c	h->1	
oda e	x->1	
oda f	ö->8	
oda g	r->1	
oda h	u->1	ä->1	
oda i	d->1	
oda k	v->1	
oda l	i->1	o->1	
oda n	y->1	
oda o	c->3	
oda p	l->2	
oda r	e->4	
oda s	a->1	
oda t	i->3	
oda v	i->3	
oda.V	a->1	
odac 	b->2	o->1	
odac"	,->1	
odac-	s->1	
odafo	n->1	
odas 	u->2	
odas.	B->1	D->2	
odda.	 ->1	
odde 	a->1	d->3	p->4	
odds 	e->1	
odelb	a->1	
odell	 ->3	"->2	.->1	e->6	
oden 	1->6	2->13	J->1	b->1	e->1	f->3	h->3	i->2	k->1	o->3	s->1	v->1	ä->1	
oden,	 ->3	
oden.	 ->1	A->1	D->1	H->1	K->1	M->1	S->1	
odens	 ->2	
oder 	d->1	h->1	i->1	o->4	p->1	s->2	v->2	ä->1	
oder,	 ->4	
oder.	A->1	D->3	I->1	K->1	
odera	t->1	
oderm	a->1	
odern	 ->5	,->1	a->8	i->24	t->1	
oders	k->3	m->1	
odert	i->1	
odet 	a->4	i->1	s->1	
odfil	m->1	
odi a	t->2	v->1	
odi b	e->1	
odi h	a->2	
odi i	n->1	
odi l	o->1	ä->1	
odi o	c->5	
odi s	o->1	
odi t	a->2	
odi, 	v->1	
odi.S	o->1	
odi.V	i->1	
odi; 	m->1	
odifi	e->5	
odiga	 ->3	
odigt	 ->1	
odins	k->1	
odis 	l->1	p->2	s->1	u->1	v->2	
odisk	a->14	u->1	
odjur	 ->1	,->1	
odkän	d->25	n->46	t->18	
odlar	e->2	n->1	
odlig	e->12	
odlin	g->2	
odo.D	e->1	
odo.H	e->1	
odo.O	m->1	
odont	 ->1	
odose	d->1	
ods a	n->1	
ods b	å->1	
ods i	n->1	
ods l	i->1	
ods o	c->1	
ods p	å->18	
ods s	k->2	o->2	
ods t	a->1	
ods v	e->1	
ods ö	k->1	
ods, 	t->1	
ods. 	D->1	
ods.B	e->1	
ods.D	e->1	
ods.U	n->1	
ods; 	b->1	
odsNä	s->1	
odset	 ->1	s->1	
odta 	a->1	d->2	f->1	g->1	n->1	u->1	ä->3	
odta.	D->1	
odtag	b->15	i->2	
odtar	 ->3	
odtas	 ->4	.->3	
odtog	 ->1	s->1	
odtyc	k->6	
oduce	n->22	r->9	
odugl	i->1	
odukt	 ->5	,->1	e->14	i->31	s->2	
odwil	l->1	
oebbe	l->1	
oedte	r->14	
oeffe	k->2	
oeffi	c->1	
oefte	r->1	
oegen	t->5	
oek s	o->1	
oekon	o->9	
oelig	?->1	
oelva	 ->1	
oende	 ->93	"->1	,->3	.->10	f->2	k->1	r->1	s->1	t->12	v->6	
oenig	h->4	
oense	 ->4	
oerhö	r->12	
oersä	t->1	
oet a	t->1	
oetis	k->1	
oette	r->5	
oetti	c->1	
of - 	a->1	
of av	 ->1	
of el	l->1	
of ex	t->1	
of fö	r->5	
of ha	d->1	r->1	
of i 	f->1	
of in	n->1	t->1	
of ku	n->1	
of li	k->1	
of oc	h->1	k->1	
of so	m->4	
of th	e->1	
of ut	a->1	
of äg	t->1	
of, h	a->1	
of, m	e->1	
of, o	c->1	
of, s	o->1	
of.De	t->1	
of.Dä	r->1	
of.En	d->1	
of.Ja	g->1	
ofala	 ->1	
ofant	l->2	
ofdra	b->1	
ofede	r->1	
ofelb	a->1	
ofem 	å->2	
ofen 	d->1	g->1	i->1	l->1	m->4	o->1	u->2	v->1	ä->1	
ofen,	 ->5	
ofen.	D->1	F->1	
ofer 	a->1	e->1	h->2	i->5	m->2	p->1	s->3	u->1	ä->1	
ofer"	 ->1	
ofer,	 ->5	
ofer.	D->2	N->1	V->2	
ofern	a->4	
ofess	i->1	o->6	
offen	s->3	t->77	
offer	 ->9	,->3	t->1	
offic	i->5	
offra	d->1	r->1	
offre	n->14	
ofhjä	l->1	
ofi o	c->1	
ofi s	o->1	
ofi, 	m->1	
ofil 	u->1	
ofil.	D->1	L->1	
ofils	k->1	
ofin 	i->1	
ofin-	r->2	
ofina	n->1	
ofisk	a->1	
ofobi	n->1	
ofred	.->1	
ofrån	k->3	
ofsit	u->1	
ofstr	a->1	
ofstö	d->2	
oft l	a->1	
ofta 	a->3	b->4	d->1	e->1	f->3	g->2	h->5	i->2	k->1	l->1	m->1	n->2	o->4	s->8	t->2	u->3	v->1	ä->5	
ofta.	O->1	
oftar	e->3	
oftas	t->1	
ofull	s->2	
oföra	k->1	
oförd	e->2	
oföre	n->5	t->1	
oförf	ö->1	
oförk	l->1	
oförl	å->2	
oförm	å->5	
oförs	i->1	k->1	t->1	
ofört	j->1	r->1	
oförä	n->2	
og 19	9->1	
og ak	t->1	
og at	t->4	
og av	 ->1	
og ba	r->1	
og be	f->1	g->2	
og de	 ->1	n->2	t->1	
og di	s->1	
og en	 ->3	
og er	,->1	
og et	t->3	
og ev	e->1	
og fa	s->1	
og fr	a->1	
og fö	r->3	
og ha	d->1	r->1	
og he	l->1	
og hä	n->1	
og i 	B->1	b->1	d->4	h->1	k->1	
og in	t->1	
og ka	n->1	
og ko	m->3	
og la	g->4	
og lä	r->1	
og ma	n->1	
og me	d->7	l->2	
og må	n->2	
og ni	 ->1	
og no	t->1	
og oc	k->2	
og om	 ->1	b->1	
og pa	r->1	
og på	s->1	
og re	d->1	s->2	
og rå	d->1	
og si	n->1	
og so	m->4	
og st	o->1	ä->1	
og ti	l->3	
og up	p->9	
og vi	s->1	
og är	 ->1	
og åt	g->1	
og ök	a->1	
og, i	 ->1	
og, o	c->1	
og, v	i->1	
og.Da	l->1	
og.De	n->1	
og.Fr	å->1	
og.Fö	r->1	
og.Ha	n->1	
og.Ja	g->2	
og.Me	n->1	
og.Mö	j->1	
og.Nä	r->1	
og.Sa	m->1	
oga a	t->4	v->1	
oga f	å->1	ö->4	
oga m	e->2	
oga p	å->1	
oga s	å->1	
oga ö	v->1	
oga, 	m->1	
oga.J	a->1	
oga.V	i->1	
ogad.	M->1	
ogade	.->1	s->1	
ogam 	g->1	
ogam,	 ->1	
ogand	e->11	
ogans	 ->1	
ogant	 ->1	
ogar 	d->1	e->1	m->1	ö->5	
ogar,	 ->1	
ogar.	T->1	
ogarn	a->7	
ogat 	f->1	r->1	t->1	
ogati	v->1	
ogau 	f->3	o->1	s->3	
ogau,	 ->5	
ogau.	E->1	
ogauM	e->1	
ogaub	e->1	
ogaus	 ->3	
ogber	o->1	
oge f	ö->1	
oge, 	m->1	
ogen 	h->1	m->5	n->1	p->2	å->1	
ogen,	 ->2	
ogen.	D->2	K->1	
ogena	 ->1	,->1	
ogenh	e->27	
ogeno	m->2	
ogent	 ->1	.->1	
oger 	a->1	o->1	
oget 	h->1	s->1	
oggra	n->12	
ogi -	 ->2	
ogi o	c->2	
ogi..	 ->1	
ogi.V	å->1	
ogik 	o->1	
ogik,	 ->2	
ogik.	F->1	H->1	V->1	
ogike	n->2	
ogin,	 ->1	
ogisk	 ->5	a->18	t->11	
ogjor	d->1	
ogkul	t->1	
ogm e	l->1	
ogmat	i->1	
ograf	i->14	
ogram	 ->75	,->17	.->20	?->2	a->1	f->1	m->108	p->11	r->1	u->1	v->1	
ogres	s->1	
ogrik	e->1	
ogrun	d->3	
ogs -	,->1	
ogs a	l->1	v->4	
ogs b	o->1	
ogs d	e->1	
ogs e	n->1	
ogs i	 ->3	
ogs k	l->2	
ogs m	e->3	
ogs n	ä->1	
ogs o	c->2	
ogs p	å->1	
ogs s	o->1	
ogs t	i->1	
ogs u	n->1	p->2	
ogs, 	a->1	f->1	
ogsar	b->1	
ogsav	v->1	
ogsbr	u->6	
ogser	a->1	
ogsfa	s->1	
ogsko	m->1	
ogsom	r->1	
ogspo	l->1	
ogsse	k->4	
ogsut	r->1	
ogsvå	r->1	
ogsäg	a->2	
oguei	r->1	
ogynn	s->1	
ogård	a->1	
ogör 	f->1	
ogöra	 ->4	
ogöre	l->3	
ogörs	 ->1	
ohand	e->3	
ohere	n->1	
ohjam	o->1	
ohjäl	p->1	
ohol,	 ->1	
ohämm	a->1	
ohövl	i->1	
oigen	k->1	
oij-v	a->1	
oinsk	r->2	
ointr	e->4	
oire 	h->1	
oire,	 ->1	
oire-	A->1	
oirmo	u->1	
ois M	i->1	
oise 	G->1	
oisk 	k->1	
oissy	s->1	
oisti	s->2	
ojala	 ->2	
ojali	s->4	t->1	
ojekt	 ->29	,->6	.->2	?->2	a->2	e->23	
ojkan	 ->1	
ojkot	t->1	
ojos 	a->1	
ojust	 ->3	,->1	.->2	
ojäml	i->5	
ojämn	.->1	a->1	
ok av	 ->1	
ok de	t->1	
ok fö	r->2	
ok gj	o->1	
ok he	l->1	
ok i 	h->1	
ok me	d->1	
ok oc	h->2	
ok om	 ->7	
ok sa	d->1	
ok sk	u->1	
ok so	m->2	
ok ti	l->1	
ok är	 ->2	
ok, d	e->1	
ok, f	ö->1	
ok, k	o->1	
ok, m	e->1	
ok, s	å->1	
ok.De	t->1	
ok.Hu	r->1	
ok.Ja	g->1	
ok.Ta	c->1	
ok.Vi	 ->1	
oka h	å->1	
oka s	o->1	
okal 	a->1	b->1	n->2	s->3	
okala	 ->31	
okali	s->3	
okalp	a->1	
okalt	 ->2	
okast	 ->1	
okat 	m->2	
okat.	H->1	
okate	r->2	
oken 	a->3	e->1	f->6	i->3	m->3	o->7	s->6	u->1	ä->1	
oken,	 ->1	
oken.	D->2	H->1	M->1	
oken:	 ->1	
okens	 ->1	
okeri	n->1	
okig 	s->1	
okigt	 ->1	
oklad	 ->1	
oklam	e->1	
oklan	d->2	
oklar	 ->2	.->1	a->2	h->5	t->2	
oko C	a->5	
okoll	 ->6	.->3	e->17	
okonf	l->1	
okont	r->2	
okor 	a->1	
okrat	 ->2	e->22	i->114	
okred	i->2	
okrig	e->1	
okrit	i->1	
okrän	k->1	
okslu	t->1	
oksta	v->1	
okt d	e->2	
okt s	ä->2	
okt v	å->1	
oktob	e->8	
okult	u->3	
okume	n->46	
okunn	i->2	
okuns	k->1	
okus 	f->1	
okus.	D->1	
okuse	r->3	
okänd	 ->1	
okäns	l->1	
ol at	t->1	
ol av	v->1	
ol be	h->1	
ol dä	r->1	
ol fö	r->2	
ol i 	A->1	E->1	
ol in	t->1	
ol me	d->1	
ol må	s->1	
ol oc	h->9	
ol so	m->4	
ol ti	l->1	
ol vi	d->1	
ol, d	e->1	
ol, e	t->1	
ol, i	 ->1	
ol, o	c->1	m->1	
ol, p	o->1	
ol, t	o->1	
ol- o	c->1	
ol-fö	r->1	
ol.De	n->1	
ol.Et	t->1	
ol.Eu	r->1	
ol.He	r->1	
ol.Kä	r->1	
ol.Me	n->1	
ol; f	ö->1	
ola d	e->2	
ola f	ö->1	
ola s	i->1	
ola v	i->1	
ola ä	r->1	
ola, 	s->1	
oladd	a->1	
olag 	o->1	s->2	
olag,	 ->1	
olage	n->6	t->2	
olagl	i->4	
olan 	1->1	s->2	u->1	v->1	
olan,	 ->1	
olan.	S->1	U->1	
olan?	H->1	
olana	 ->2	,->2	
olanh	ö->4	
olar 	a->1	d->1	i->1	m->2	s->2	v->2	ä->3	
olar,	 ->1	
olar.	D->1	V->1	
olarn	a->8	
olars	 ->2	
olavt	a->1	
olbes	 ->2	
oldat	e->2	
oldio	x->5	
ole p	o->1	
olemi	k->1	
olen 	a->3	b->1	e->2	f->1	h->3	i->7	m->1	n->1	o->3	p->1	s->2	t->1	u->2	
olen,	 ->5	
olen.	D->2	I->1	S->1	U->1	V->2	
olens	 ->8	
olera	 ->5	.->1	n->11	
olere	r->7	
oleri	n->1	
oleum	 ->1	
olf H	i->2	
olfen	 ->2	.->2	
olfrå	g->1	
olfst	r->3	
olför	e->2	
oliba	k->1	
olicy	,->1	a->1	d->1	f->1	
olida	r->30	
olide	r->3	
olig 	f->2	ö->2	
olig,	 ->1	
oliga	 ->2	
olige	n->6	
oligt	 ->5	
olik 	m->1	
olik.	D->1	
olik:	 ->1	
olika	 ->114	,->1	.->1	
olike	r->2	
olikh	e->7	
olikt	 ->4	,->1	
olint	r->1	
olis,	 ->1	
olis.	V->1	
olis;	 ->1	
olisa	k->1	
olise	n->5	r->3	
olisi	ä->1	
olisk	 ->2	,->1	.->1	a->2	
olism	 ->1	y->2	
oliss	a->1	t->1	
olisv	ä->1	
olita	n->1	
oliti	c->1	k->309	s->223	
oliv 	k->1	t->1	
oliv.	I->1	
olja 	f->1	i->2	s->1	
olja,	 ->2	
olja.	T->1	
oljan	 ->2	,->1	
oljeb	e->1	o->4	ä->8	
oljef	ö->1	
oljei	n->3	
oljek	o->2	
oljes	k->1	
oljet	a->8	r->2	
oljeu	t->2	
olk a	t->1	
olk b	l->1	o->1	
olk h	a->1	
olk i	 ->2	
olk o	c->2	
olk r	e->1	
olk s	k->1	o->2	
olk t	v->1	
olk u	p->1	
olk, 	d->1	
olk.A	t->1	
olk.D	e->1	
olk.M	e->1	
olk.O	c->1	
olk.V	i->4	
olka 	d->1	f->1	m->1	u->1	
olkad	e->1	
olkar	 ->3	n->2	
olkas	 ->4	,->1	.->1	
olkat	s->1	
olken	 ->2	s->4	
olkes	t->1	
olket	 ->5	,->1	.->1	:->1	i->2	s->4	
olkfr	o->1	
olkgr	u->2	
olkhä	l->9	
olkli	g->1	
olkni	n->57	
olkom	r->6	
olkon	v->1	
olkpa	r->10	
olkre	g->1	p->3	
olkrä	t->1	
olks 	f->1	s->2	
olkst	y->1	
olksw	a->1	
olksä	g->1	
olkva	l->2	
oll -	 ->1	
oll E	u->1	
oll a	n->1	t->3	v->17	
oll d	e->2	
oll f	o->1	r->1	ö->6	
oll g	e->1	ö->1	
oll i	 ->16	n->3	
oll k	a->1	o->1	
oll m	å->1	
oll n	y->1	ä->2	
oll o	c->6	m->1	
oll p	å->1	
oll s	o->11	t->1	
oll u	t->1	
oll v	a->1	i->2	o->1	
oll ä	r->3	
oll ö	v->5	
oll!J	a->1	
oll, 	a->1	d->1	f->2	h->1	i->1	m->1	n->1	o->3	p->1	s->3	u->1	v->2	ä->2	
oll- 	o->1	
oll.D	e->5	
oll.E	n->1	
oll.F	i->1	r->1	
oll.H	ä->1	
oll.I	 ->1	n->1	
oll.J	a->3	
oll.K	o->2	
oll.M	å->1	
oll.P	r->1	å->1	
oll.S	m->1	o->1	
oll.T	a->1	ä->1	
oll.U	t->1	
oll.V	i->3	å->1	
oll: 	e->1	
ollan	t->1	
ollar	 ->3	,->3	;->1	n->2	
olleg	a->62	e->127	i->4	o->3	
ollek	t->10	
ollen	 ->20	,->1	.->5	Ä->1	
oller	 ->14	.->6	;->1	a->34	n->5	
ollet	 ->12	.->4	
ollfu	n->1	
ollis	i->3	
ollma	k->1	
ollmy	n->1	
ollmä	r->1	
ollmö	j->2	
ollni	n->1	s->1	
ollom	r->1	
ollor	g->1	
ollri	s->1	
ollsb	e->1	
ollsy	s->3	
ollut	i->1	s->14	
ollve	r->1	
ollyw	o->1	
olm d	e->1	
olm, 	h->1	
olm.H	e->1	
oln o	c->1	
olog,	 ->1	
ologi	 ->3	n->1	s->26	
oloni	a->1	
olor 	o->1	s->1	
olor,	 ->1	
oloss	a->1	
olpe 	p->1	
ols a	r->1	
ols m	e->1	
ols u	p->1	
olsav	g->1	
olsbu	r->1	
olsfa	l->1	
olsfö	r->1	
olsit	u->1	
olska	 ->3	n->1	
olske	n->1	
olspr	o->1	
olssy	s->1	
olstv	i->1	
olsut	s->1	
olsvä	s->1	
olt ö	v->6	
olta 	o->1	ö->2	
olthe	t->2	
olunt	a->4	
olut 	a->1	b->5	d->1	e->1	f->3	i->8	l->1	m->2	n->10	r->1	s->2	t->2	ä->1	
oluta	 ->3	
oluti	o->100	
olv å	r->1	
olver	a->9	
olvet	 ->1	
olyck	a->19	l->4	o->16	s->9	
olym 	a->1	o->1	
olyme	n->1	r->1	
olymp	i->1	
olzma	n->2	
olämp	a->1	l->3	n->1	
olöst	a->2	
om "E	q->1	u->1	
om "K	v->1	
om "n	å->1	
om "o	r->1	
om "v	a->1	
om "ö	p->1	
om - 	a->3	k->1	m->1	o->1	p->1	t->1	v->2	
om 1 	0->1	
om 15	0->1	
om 16	 ->1	
om 19	8->1	9->1	
om 20	 ->2	
om 28	 ->1	
om 3-	l->2	
om 31	4->1	
om 35	 ->2	0->1	
om 40	 ->2	0->1	
om 45	 ->1	
om 5b	-->1	
om 6,	0->1	
om Ag	u->1	
om Ah	e->1	
om Al	a->1	p->1	
om Am	o->1	s->2	
om Ap	a->1	
om At	l->1	
om BS	E->1	
om Ba	r->1	
om Be	l->1	r->5	
om Bl	a->1	
om Bo	w->1	
om Br	i->1	y->1	
om CE	N->1	
om Ce	y->1	
om Co	c->1	x->1	
om Da	 ->1	l->1	n->2	
om De	 ->1	
om Di	m->1	
om Du	t->1	
om EG	-->3	
om EM	U->1	
om EU	 ->11	,->1	-->2	.->3	:->2	
om Eh	u->1	
om El	l->1	
om Er	i->1	
om Et	i->1	
om Eu	r->72	
om FB	I->1	
om FP	Ö->1	
om Fl	o->1	
om Fr	a->2	
om Fö	r->4	
om GU	S->1	
om Ga	l->1	
om Ge	n->2	
om Go	l->1	o->1	
om Gr	e->2	
om Ha	i->3	t->2	
om He	d->1	
om Hi	t->1	
om IN	T->1	
om In	d->1	
om Ir	l->1	
om Is	r->1	
om It	a->2	
om Jo	n->2	
om Jö	r->2	
om Ka	u->1	
om Ko	s->4	u->1	
om La	n->6	
om Li	b->1	
om Ll	o->1	
om Ma	l->1	r->1	
om Mc	C->1	N->1	
om Ne	d->1	
om Of	f->1	
om PP	E->1	
om Pa	k->1	l->1	y->1	
om Po	r->1	w->3	
om Pr	o->1	
om Ra	c->1	
om Ri	c->1	
om Ro	t->1	
om SE	K->1	
om Sc	h->2	
om Se	i->2	
om Sj	ä->1	
om Sk	o->1	
om Sp	e->1	
om Ta	m->1	
om Th	e->3	
om Ti	b->2	
om To	r->1	t->1	
om Tu	r->4	
om Vä	r->1	
om Wa	l->2	
om Wi	e->1	
om a 	p->1	
om ab	s->2	
om ad	v->2	
om ag	e->3	r->1	
om al	d->1	l->52	
om am	b->1	e->1	
om an	d->9	f->2	g->3	k->1	l->2	n->2	o->1	s->25	t->13	v->8	
om ap	p->1	
om ar	b->17	g->1	r->1	t->2	
om as	y->3	
om at	t->334	
om av	 ->14	f->2	g->6	k->2	l->2	s->10	t->1	v->2	
om b)	 ->1	
om ba	k->2	l->1	n->1	r->3	
om be	a->2	d->8	f->8	g->7	h->29	k->10	m->1	o->1	r->14	s->26	t->15	v->6	
om bi	d->7	l->2	n->1	o->1	t->1	
om bl	.->2	a->2	e->2	i->2	y->1	
om bo	r->12	s->2	t->1	
om br	i->3	o->4	u->1	y->2	å->3	
om bu	d->3	
om by	g->1	r->1	
om bä	r->5	t->2	
om bå	d->5	
om bö	c->1	r->14	t->1	
om c)	 ->1	
om ca	n->1	
om ce	n->1	
om ch	a->1	o->1	
om co	r->1	
om da	g->6	
om de	 ->152	,->1	b->2	c->1	f->2	l->6	m->6	n->142	r->1	s->33	t->271	
om di	a->1	f->1	o->1	r->7	s->7	
om dj	ä->1	
om do	g->1	m->4	
om dr	a->12	i->3	y->1	
om du	b->1	
om dy	k->1	
om dä	r->8	
om då	 ->4	l->1	
om dö	d->1	e->1	m->1	
om ef	f->3	t->5	
om eg	e->4	n->1	
om ej	 ->1	
om ek	o->5	
om el	e->1	l->1	
om em	e->1	
om en	 ->164	d->6	e->5	h->1	l->3	s->3	
om er	 ->3	a->4	k->1	s->1	t->4	ö->1	
om et	t->98	
om eu	r->8	
om ex	 ->1	a->2	c->2	e->9	p->1	
om fa	d->1	k->3	l->7	r->1	s->11	t->8	
om fe	m->2	
om fi	c->1	n->38	s->4	
om fj	o->1	
om fl	a->1	e->5	y->5	
om fo	d->1	l->2	n->1	r->16	s->1	
om fr	a->27	e->6	i->8	u->2	ä->1	å->16	
om fu	l->1	n->3	s->1	
om fy	l->1	r->1	
om fä	l->1	r->1	
om få	r->6	t->3	
om fö	l->7	r->201	
om ga	m->1	r->5	v->1	
om ge	 ->2	m->18	n->14	r->9	s->4	t->1	
om gi	c->1	l->1	v->1	
om gj	o->10	
om gl	o->1	
om go	d->8	
om gr	a->2	i->2	u->10	ä->2	
om gä	l->22	
om gå	r->9	t->2	
om gö	m->1	r->33	
om ha	 ->1	d->3	m->3	n->42	r->143	s->1	v->2	
om he	d->1	l->51	r->3	
om hi	n->2	t->12	
om hj	ä->6	
om ho	b->1	n->10	t->3	
om hu	m->2	r->32	
om hy	s->1	
om hä	l->2	n->16	r->13	v->4	
om hå	l->7	r->1	
om hö	g->4	r->3	
om i 	B->1	E->1	H->1	N->1	T->2	U->1	a->2	b->1	d->26	e->2	f->12	g->1	h->6	l->1	m->2	n->1	o->2	p->5	r->3	s->15	t->1	v->6	å->1	
om ic	k->4	
om id	é->1	
om if	a->1	r->1	
om ig	e->1	
om ih	å->1	
om in	 ->1	b->1	d->6	f->12	g->11	i->1	k->1	l->9	n->28	o->4	r->5	s->4	t->99	v->3	
om is	r->1	
om ja	g->133	
om jo	r->6	
om ju	 ->5	s->8	
om jä	m->2	r->1	
om ka	n->54	p->4	r->5	
om ke	m->1	
om kl	a->2	
om ko	d->1	l->4	m->138	n->28	r->10	s->5	
om kr	a->3	i->6	ä->17	
om ku	l->7	n->1	r->1	
om kv	i->1	
om kä	n->6	r->6	
om kö	p->1	r->1	
om la	d->4	g->12	n->2	
om le	d->30	g->1	t->1	v->6	
om li	b->2	g->16	k->4	t->2	v->16	
om lj	u->1	
om lo	k->1	
om ly	c->2	d->1	f->1	k->1	s->1	
om lä	c->1	g->7	k->1	m->10	n->4	t->1	
om lå	g->2	n->1	
om lö	s->2	
om ma	i->1	j->2	k->1	n->87	r->3	x->1	
om me	d->40	l->2	n->2	r->3	s->1	
om mi	l->8	n->17	s->4	t->1	
om mo	d->3	t->11	
om mu	s->1	
om my	c->7	n->8	
om mä	n->13	r->1	
om må	h->1	l->2	n->4	s->25	
om mö	j->51	
om na	r->1	t->9	z->3	
om ne	d->2	g->1	k->1	
om ni	 ->55	,->5	.->1	o->1	
om no	r->1	
om nu	 ->24	m->1	
om ny	 ->1	a->2	l->2	s->1	t->1	
om nä	m->5	r->6	s->1	
om nå	g->26	
om nö	d->1	t->1	
om oa	c->1	
om ob	e->2	
om oc	h->18	k->18	
om of	f->3	t->4	
om og	e->1	
om ol	i->3	j->2	y->1	
om om	 ->23	b->1	e->1	f->4	l->1	r->9	s->1	ö->1	
om on	ö->1	
om or	d->11	i->1	o->2	s->3	
om os	s->4	
om ot	i->1	
om pa	r->23	
om pe	k->2	n->2	r->3	
om pl	a->4	
om po	l->5	s->1	ä->1	
om pr	a->2	e->3	i->7	o->10	
om pu	b->1	m->1	
om på	 ->25	g->1	m->1	p->1	t->2	v->8	
om ra	d->1	m->51	p->1	s->2	t->1	
om re	d->34	f->8	g->23	l->7	p->1	s->12	t->1	v->2	
om ri	k->4	m->2	s->8	
om ro	l->1	
om ru	l->2	s->1	
om ry	g->1	s->1	
om rä	c->1	k->1	t->13	
om rå	d->35	
om rö	r->13	s->3	v->1	
om s.	k->1	
om sa	d->2	g->4	k->5	m->33	n->1	t->2	
om sc	h->1	
om se	d->5	g->2	k->2	n->1	r->5	x->1	
om si	n->6	t->5	
om sj	u->2	ä->1	ö->1	
om sk	a->69	e->12	i->3	o->5	r->7	u->25	y->5	ö->1	
om sl	o->1	u->5	
om sm	å->3	
om sn	a->2	e->1	
om so	c->2	l->1	m->3	
om sp	e->8	o->1	r->2	
om st	a->14	e->1	i->1	o->2	r->10	y->3	ä->14	å->22	ö->14	
om su	b->4	
om sv	a->3	
om sy	f->8	n->2	s->8	
om sä	g->2	k->14	r->3	t->1	
om så	 ->16	d->8	l->1	t->1	
om sö	k->1	r->2	
om t.	e->2	o->1	
om ta	g->2	l->6	r->6	s->5	x->1	
om ti	b->1	d->11	l->60	o->1	
om tj	ä->3	
om to	g->5	l->5	
om tr	a->16	e->3	o->2	ä->5	
om tu	r->1	
om tv	e->1	å->4	
om ty	c->2	d->5	n->1	s->1	v->2	
om tä	c->2	n->1	p->1	
om un	d->17	i->22	
om up	p->35	
om ur	 ->1	s->7	
om ut	.->1	a->5	b->5	d->1	e->1	f->7	g->11	j->1	l->2	m->2	n->1	r->1	s->12	t->13	v->11	ö->1	
om va	d->16	g->1	l->3	n->4	r->35	
om ve	d->1	l->1	m->2	r->17	t->4	
om vi	 ->253	,->3	?->1	a->1	d->10	k->1	l->38	n->1	s->24	t->5	
om vo	n->3	r->2	
om vr	ä->1	
om vu	x->1	
om vä	c->2	g->3	l->4	n->2	r->1	s->1	
om vå	r->17	
om yr	k->1	
om yt	t->3	
om Ös	t->4	
om äg	e->2	n->1	t->1	
om än	 ->4	d->15	n->4	t->3	
om är	 ->176	
om ät	e->1	
om äv	e->14	
om åk	t->1	
om ål	a->1	i->1	
om år	e->3	s->1	
om ås	t->1	y->4	
om åt	e->17	g->4	m->1	
om öa	r->1	
om ök	a->3	
om öm	s->1	
om ön	s->1	
om öp	p->7	
om ör	o->1	
om ös	t->2	
om öv	e->16	r->1	
om!Tr	o->1	
om".D	e->1	
om) o	m->1	
om); 	a->1	
om, a	n->1	t->3	v->1	
om, d	e->7	
om, e	f->2	n->2	
om, f	r->1	
om, g	r->1	
om, h	a->1	e->2	
om, i	 ->4	
om, j	a->1	u->1	
om, k	v->1	
om, l	e->1	
om, m	e->2	
om, n	i->1	ä->1	
om, o	c->4	m->1	
om, p	å->1	
om, s	a->1	o->2	ä->1	
om, t	r->1	
om, u	p->1	t->3	
om, v	a->1	i->3	
om, ä	r->1	v->5	
om- o	c->1	
om. D	å->1	
om. H	u->1	
om.Av	s->1	
om.De	 ->1	n->2	s->1	t->5	
om.Dä	r->1	
om.EK	S->1	
om.Ex	p->1	
om.He	r->1	
om.Hu	r->1	
om.In	f->1	
om.Ja	g->7	
om.Me	d->1	n->3	
om.Nä	r->1	
om.Oc	h->1	
om.St	a->1	
om.Så	 ->1	
om.Vi	 ->3	
om/ri	k->1	
omI. 	f->1	
omade	 ->1	
omagn	a->1	
omane	r->1	
omano	 ->2	
omar 	a->2	f->3	i->2	o->1	ö->1	
omar,	 ->3	
omar.	B->1	H->1	
omarb	e->2	
omare	 ->2	,->1	.->2	
omark	o->1	
omarn	a->8	
omate	r->1	
omati	,->1	k->1	s->16	
omb h	a->1	
omb.A	n->1	
ombad	s->1	
ombar	d->1	
ombat	t->2	
ombed	s->1	
omben	 ->1	
omber	 ->1	,->1	
ombes	ö->2	
ombet	t->2	
ombex	p->1	
ombin	a->1	
ombli	c->5	
ombni	n->1	
ombor	d->1	
ombro	t->2	
ombud	 ->2	s->10	
omdef	i->1	
omdir	i->1	
omdri	v->6	
omdöm	e->2	
omede	l->18	
omedg	ö->2	
omedv	e->1	
omen 	a->1	b->1	i->2	o->3	s->1	t->1	ö->1	
omen,	 ->3	
omen.	D->1	
omene	r->3	t->2	
oment	 ->3	.->2	
omer 	N->1	v->1	
omer,	 ->3	
omera	d->4	
omern	a->1	
omes,	 ->1	
omet 	s->1	
omete	r->1	
omeur	o->4	
omfat	t->83	
omfly	t->1	
omfor	m->3	s->1	
omfån	g->2	
omför	 ->8	a->120	b->7	d->5	h->1	s->12	t->9	
omger	 ->1	
omgic	k->1	
omgiv	a->1	n->1	
omgri	p->4	
omgå 	e->1	
omgå.	F->1	
omgåe	n->1	
omgån	g->5	
omgår	 ->3	.->1	
omgåt	t->2	
omhul	d->1	
omi -	 ->1	
omi a	t->1	
omi m	e->5	
omi o	c->12	
omi ä	r->1	
omi, 	l->1	m->1	
omi.D	e->2	
omi.F	ö->1	
omi? 	O->1	
omier	 ->1	,->1	.->1	n->5	
omin 	-->1	d->1	i->2	k->2	o->10	s->4	
omin,	 ->2	
omin.	C->1	D->1	L->1	M->1	V->1	
omina	n->1	
omine	r->10	
omins	 ->3	
omisk	 ->45	a->142	t->28	
omiss	 ->6	,->5	.->2	a->2	e->1	f->2	l->1	r->2	t->1	
omist	l->1	y->4	
omkri	n->15	
omlas	t->1	
omlig	 ->1	a->6	e->1	g->1	t->9	
omlok	a->2	
omläs	n->2	
omma 	a->9	d->5	e->4	f->13	h->2	i->23	l->3	m->11	n->3	o->1	p->4	r->2	s->3	t->12	v->1	å->1	ö->5	
omma,	 ->1	
omma.	J->2	O->1	
omman	d->55	
ommar	 ->1	e->1	l->1	
ommas	 ->1	
ommel	s->15	
ommen	.->1	;->1	d->45	t->37	
ommer	 ->714	,->4	.->4	s->8	
ommet	 ->2	.->3	
ommis	s->1150	
ommit	 ->37	,->3	.->2	s->2	t->59	
ommon	 ->1	
ommor	 ->1	,->1	
ommun	.->1	a->3	e->10	i->19	
ommöb	l->1	
omna 	e->2	f->1	h->1	i->2	m->1	o->1	r->3	s->1	t->1	
omna,	 ->1	
omna.	T->1	
omnan	d->1	
omnar	 ->27	.->1	
omnas	 ->1	
omofo	b->1	
omoge	n->2	
omora	l->1	
omord	e->7	
omorg	a->2	
omose	x->1	
ompas	s->1	
ompen	s->10	
ompet	e->11	
ompla	n->1	
omple	m->10	t->14	x->4	
ompli	c->12	m->4	
ompon	e->4	
ompro	m->22	
omprö	v->8	
omrin	g->1	
omrum	 ->1	,->1	
områd	e->316	
omrös	t->42	
oms f	ö->1	
oms s	ä->1	
oms- 	o->2	
oms-,	 ->1	
omsa 	d->2	u->1	
omsar	 ->1	
omsbr	o->1	
omsfr	å->3	
omsfu	l->1	
omsgr	ä->1	
omshe	m->1	
omski	n->1	
omsla	g->3	
omslu	t->3	
omsni	t->11	
omsor	g->9	
omspl	i->1	
omspä	n->1	
omsrä	t->1	
omst 	f->1	i->1	o->1	p->3	u->1	
omste	n->2	r->6	
omstf	ö->1	
omsth	ä->1	
omstk	ä->1	
omsto	l->86	
omstr	a->1	i->4	u->10	
omstä	l->1	n->34	
omstå	e->2	
omsve	p->1	
omsvä	t->1	
omsyr	a->3	
omsät	t->8	
omtal	a->1	
omtän	k->1	
omull	,->1	
omvan	d->5	
omväg	 ->1	e->1	
omväl	v->4	
omvän	d->4	t->1	
omväx	l->1	
omán,	 ->1	
omäss	i->1	
omål 	o->1	t->1	
omåle	t->1	
omé o	c->1	
omé p	e->1	
oméav	t->1	
oméko	n->1	
omés 	R->1	
omöjl	i->16	
on (A	5->5	
on (f	ö->2	
on - 	e->1	m->1	o->2	s->1	
on 12	/->3	4->2	
on 19	6->1	
on 34	.->1	
on 52	0->1	
on 57	,->1	
on Ac	t->1	
on Bo	e->1	
on Ei	e->1	
on Ha	r->1	
on I 	o->1	
on Pr	o->2	
on VI	I->2	
on Va	l->3	
on Wo	g->17	
on al	l->2	
on an	d->1	l->2	n->6	s->2	t->2	
on ap	p->1	
on ar	a->1	
on at	t->6	
on av	 ->24	f->2	s->1	
on be	d->1	g->1	k->1	s->2	t->3	
on bi	t->1	
on bl	i->1	
on bo	r->1	
on bä	r->2	
on bö	r->1	
on ch	a->1	
on de	l->2	n->1	
on dä	r->8	
on då	l->1	
on ef	f->3	t->3	
on el	l->2	
on en	 ->2	b->1	d->1	s->1	
on et	t->1	
on eu	r->1	
on fa	r->1	
on fo	r->1	
on fr	å->5	
on fu	n->1	
on få	r->1	
on fö	l->1	r->32	
on ge	n->3	
on gr	u->1	
on gå	n->7	r->1	
on gö	r->1	
on ha	 ->1	d->2	r->10	
on ho	s->1	
on hä	r->2	v->1	
on hö	r->1	
on i 	E->3	F->1	K->2	L->2	S->1	a->1	b->2	d->7	e->1	m->1	p->2	r->2	s->3	v->1	
on id	é->1	
on in	f->2	n->4	o->6	r->1	s->1	t->3	
on ja	g->1	
on ju	r->1	s->2	
on ka	n->12	t->1	
on kl	.->12	
on ko	l->2	m->9	n->4	
on la	g->2	w->1	
on li	g->1	k->1	
on ly	s->1	
on lö	n->1	
on m.	m->1	
on me	d->15	l->3	n->1	
on mi	l->1	n->1	
on mo	d->1	t->3	
on my	c->1	
on må	n->1	s->1	
on mö	j->2	
on ne	g->1	
on ni	 ->1	
on ny	t->4	
on nä	r->2	
on oc	h->40	k->1	
on of	f->1	
on ol	i->1	j->1	y->1	
on om	 ->16	,->1	.->1	f->1	p->1	
on or	d->1	g->1	
on ov	a->1	
on pe	r->2	
on pl	a->2	
on pr	o->1	
on på	 ->14	m->1	p->1	
on re	d->2	s->1	
on ri	s->2	
on ro	l->1	
on rä	t->3	
on sa	k->1	m->3	
on se	t->1	
on sk	a->2	i->2	r->2	u->6	ö->1	
on so	m->71	r->1	
on sp	e->1	
on st	a->5	ä->1	ö->1	
on sy	s->1	
on sä	k->1	t->1	
on så	 ->2	d->2	l->1	s->2	
on ta	l->3	r->1	
on ti	l->22	
on tj	ä->1	
on tr	o->1	
on ty	v->1	
on tä	v->1	
on un	d->2	
on up	p->5	
on ur	 ->1	
on ut	g->1	t->2	
on va	r->1	
on ve	c->1	r->1	t->2	
on vi	 ->4	f->1	l->1	
on vå	r->1	
on än	 ->1	
on är	 ->11	
on år	 ->2	
on åt	e->2	g->1	
on öv	e->1	
on" p	å->1	
on) (	K->2	
on, 5	0->1	
on, D	u->1	
on, L	o->1	
on, O	l->1	
on, P	a->1	
on, S	h->1	
on, a	t->1	v->1	
on, b	a->1	e->1	l->1	
on, d	e->2	v->1	ä->2	
on, e	f->2	l->1	n->3	t->1	
on, f	i->1	ö->2	
on, h	a->1	o->1	
on, i	 ->1	g->1	n->2	
on, k	o->1	ä->2	
on, m	e->4	
on, n	u->1	ä->1	
on, o	c->10	m->2	
on, p	å->1	
on, s	a->1	o->6	å->2	
on, t	r->1	
on, u	t->1	
on, v	i->4	
on, ä	r->2	v->1	
on- o	c->1	
on-Ha	r->1	
on. D	e->1	
on. I	 ->1	
on. O	c->1	
on. R	å->1	
on.14	 ->1	
on.Av	s->1	
on.Br	i->1	
on.DE	B->1	
on.De	 ->2	n->7	t->9	
on.Dä	r->2	
on.Då	 ->1	
on.En	 ->1	l->1	
on.Ev	e->1	
on.Fl	e->1	
on.Fr	å->1	
on.Fö	l->1	r->2	
on.Gä	l->1	
on.Ha	n->1	
on.He	r->6	
on.I 	a->1	d->4	f->1	s->1	
on.Ja	c->1	g->13	
on.Ko	m->2	
on.Lå	t->1	
on.Me	n->1	
on.Mi	n->2	
on.Mö	j->1	
on.Ni	 ->1	e->1	
on.Om	 ->3	
on.Sa	m->1	
on.Se	d->1	
on.So	c->1	m->1	
on.Så	 ->1	
on.Ti	l->1	
on.Tr	o->1	
on.Un	d->1	
on.Va	d->4	l->1	
on.Vi	 ->10	l->1	
on.Å 	e->1	
on/år	)->1	,->1	
on: D	e->1	
on: a	t->1	
on: i	 ->1	
on; v	i->1	
on? D	e->1	
on? I	n->1	
on?De	n->1	
on?Ja	,->1	
on?Ka	n->2	
on?Ko	m->1	
on?Vi	 ->1	
on?Äv	e->1	
onNäs	t->1	
ona a	t->8	
ona d	e->5	
ona e	k->1	n->1	
ona h	u->1	
ona i	g->1	
ona n	å->1	
ona o	c->1	
ona s	o->1	
ona t	r->1	v->3	
ona v	a->1	i->1	
onade	 ->4	.->2	s->1	
onakr	y->1	
onal 	C->1	d->1	f->1	i->2	m->1	o->2	p->1	r->1	s->2	u->2	v->2	
onal,	 ->2	
onal-	s->2	
onal.	D->1	P->1	S->1	V->1	
onala	 ->44	
onale	k->4	n->1	
onalf	ö->3	
onali	s->21	t->7	
onall	i->1	
onalp	o->39	r->1	
onalr	e->3	ä->1	
onals	o->1	t->5	y->1	
onalt	 ->1	
onalu	t->1	
onand	e->1	
onans	l->1	
onapr	o->2	
onar 	C->1	a->3	k->1	p->1	v->1	
onar,	 ->1	
onas 	S->2	o->1	
onat 	d->1	o->1	
onat,	 ->2	
onat.	J->1	
onati	o->1	
onazi	s->2	
onbeh	a->1	
onbli	c->15	
oncen	t->31	
oncep	t->7	
oncer	n->2	
oncis	 ->1	t->1	
onckh	e->14	
ond c	i->1	
ond f	ö->4	
ond k	o->1	
ond s	o->2	
onda 	d->1	i->1	m->1	
ondag	e->2	
onde 	d->1	o->1	å->1	ö->2	
onde.	M->1	
onden	 ->26	,->9	.->5	N->1	s->4	
onder	 ->14	,->1	.->3	n->51	
ondgå	r->2	
ondit	i->1	
ondme	d->3	
ondo.	F->1	
ondon	 ->1	,->2	.->1	
ondsk	a->1	
ondsp	r->3	
ondup	p->1	
one a	n->1	t->1	
one b	l->1	
one d	e->1	
one e	k->1	
one f	o->1	
one g	ä->1	
one h	a->1	
one i	 ->2	n->3	
one j	a->1	
one k	a->1	o->1	
one l	o->1	
one n	ä->2	å->1	ö->1	
one o	m->1	
one r	y->1	
one s	å->1	
one t	o->1	
one v	a->1	i->1	
one-M	a->1	
one-s	t->1	
onell	 ->49	,->3	.->2	a->195	t->28	
onema	n->3	
onen 	(->5	-->6	C->1	E->1	I->1	P->1	a->102	b->36	d->9	e->15	f->77	g->21	h->60	i->80	k->63	l->9	m->31	n->11	o->109	p->25	r->18	s->87	t->23	u->21	v->22	ä->42	å->3	ö->4	
onen!	N->1	
onen"	.->1	
onen)	N->1	
onen,	 ->103	
onen.	 ->3	(->1	)->6	.->7	1->1	A->2	B->1	D->31	E->5	F->5	G->1	H->11	I->4	J->12	K->2	L->2	M->6	N->5	O->3	P->5	R->2	S->3	T->1	U->2	V->14	Ä->2	
onen:	 ->1	
onen;	 ->3	
onen?	H->1	K->1	V->1	Ä->1	
onenJ	a->2	
onens	 ->374	,->1	
onent	 ->1	e->3	i->1	
oner 	(->1	-->4	K->1	[->1	a->12	b->9	d->10	e->25	f->16	g->5	h->9	i->29	j->1	k->7	l->2	m->33	n->1	o->35	p->7	r->1	s->49	t->16	u->3	v->3	ä->3	å->1	
oner,	 ->42	
oner.	 ->1	(->1	A->1	B->1	D->11	F->1	G->1	H->2	I->6	J->8	K->2	L->1	M->1	N->1	S->1	T->1	V->4	Ä->1	
oner;	 ->1	
oner?	-->1	H->1	J->1	V->1	
onerN	ä->1	
onera	 ->4	d->6	n->1	r->2	s->2	
oneri	n->11	
onerl	i->2	
onern	a->181	
oners	 ->5	
onet.	D->1	
oneta	r->1	
onetä	r->6	
onfed	e->1	
onfer	e->170	
onfes	s->1	
onfid	e->2	
onfis	k->2	
onfli	k->16	
onfro	n->1	
ongen	 ->1	
ongiv	a->2	
ongre	s->1	
ongsb	e->1	
onhun	d->1	
oni o	c->2	
oni s	ä->1	
oni.(	P->1	
onial	i->1	
onik-	 ->1	
onind	e->1	
oning	 ->4	.->1	
onise	r->15	
onisk	 ->8	a->4	t->1	
onism	 ->1	,->1	.->1	
onist	i->2	
onito	r->1	
onjun	k->1	
onjuv	e->1	
onjär	e->1	
onkre	t->58	
onkur	r->285	
onlam	p->1	
onlig	 ->4	a->11	e->16	h->2	t->1	
onmär	k->2	
onmäs	s->1	
onmöt	e->2	
onnam	b->1	
onnäe	r->1	
onodl	a->2	i->1	
onoku	l->3	
onom 	-->1	2->1	d->1	e->1	f->2	h->1	m->2	n->1	o->3	p->1	s->3	t->4	ö->1	
onom,	 ->2	
onom.	 ->1	H->1	J->1	M->1	
onome	n->3	r->1	
onomi	 ->20	,->2	.->3	?->1	e->8	n->30	s->219	
onopo	l->17	
onrad	 ->1	
ons b	e->1	
ons f	r->1	
ons i	n->1	
ons p	a->1	
ons r	e->1	
ons s	c->1	v->1	
ons t	i->1	r->1	
ons v	e->1	ä->1	
ons- 	o->4	
onsaf	f->2	
onsan	a->1	
onsar	b->8	
onsav	t->1	
onsbo	l->1	
onsbr	i->1	
onsda	g->5	
onsdi	r->1	
onsdo	k->1	
onsdö	m->1	
onsek	v->61	
onser	v->7	
onsfo	r->1	
onsfr	i->2	
onsfu	n->1	
onsfö	r->19	
onsha	u->1	
onshi	n->8	
onsin	 ->10	.->1	d->1	s->1	
onska	m->1	n->1	
onsko	m->1	n->2	s->2	
onskr	a->1	
onsku	r->6	
onsle	d->11	
onslä	g->1	
onsme	d->4	
onsmo	m->1	
onsmä	s->1	
onsmö	t->1	
onsni	v->2	
onsol	i->3	
onsor	d->1	
onspa	r->1	
onspl	a->2	
onspo	l->3	
onspr	i->1	o->5	
onsra	d->1	
onsre	g->3	
onsro	l->1	
onsrä	t->12	
onssa	m->7	
onssc	h->1	
onsse	k->1	
onssk	a->1	
onsst	r->2	
onssy	s->5	
onst 	o->1	
onst,	 ->1	
onsta	b->1	n->4	t->40	
onste	k->2	r->1	
onsti	g->3	l->3	t->23	
onstj	ä->1	
onstr	a->3	e->3	u->36	
onsul	t->5	
onsum	e->61	t->2	
onsun	d->3	
onsup	p->1	
onsut	b->3	
onsvi	l->1	
onsäg	a->1	
onsäm	n->1	
onsåt	e->1	
ont a	t->1	
ont o	m->1	
ont.S	å->1	
ontai	n->1	
ontak	t->17	
ontal	a->2	s->1	
ontam	i->2	
ontan	?->1	a->1	t->3	
ontat	i->1	
ontel	l->1	
onten	 ->1	"->1	,->1	
onter	a->3	i->9	
ontex	t->1	
onti 	-->1	h->2	i->3	k->1	o->1	p->1	v->1	
onti!	 ->3	
onti,	 ->2	
onti.	J->1	V->1	
ontin	e->5	g->39	u->2	
ontor	 ->4	,->1	e->2	
ontra	k->4	p->1	s->2	
ontre	a->2	
ontro	l->180	v->4	
onven	t->24	
onver	g->5	
onvik	t->4	
onym 	m->1	s->1	
onym.	D->1	
onyma	 ->1	
onymi	t->1	
onzál	e->1	
onär 	-->2	A->1	B->9	K->5	M->13	N->1	P->17	R->2	S->2	V->4	W->1	a->1	f->2	h->1	i->1	m->1	o->1	s->1	
onär!	 ->29	.->1	E->1	J->1	
onär,	 ->74	
onär.	 ->1	D->2	G->1	J->6	V->1	
onäre	n->46	r->19	
onärs	 ->1	
onåri	n->1	
onödi	g->11	
oo fr	a->1	
ood o	m->1	
oodfi	l->1	
oods 	a->1	
oodwi	l->1	
ooij-	v->1	
ool, 	e->1	
oområ	d->1	
ooper	a->1	
oos a	t->1	
op al	l->1	
op be	t->1	
op de	t->1	
op fö	r->1	
op oc	h->1	
op om	 ->1	
op pe	r->1	
op si	n->1	
op sk	a->1	
op ti	l->1	
op ut	a->1	
op än	n->1	
op, A	r->3	
op, e	n->1	
op, o	c->1	
op, p	å->1	
op-sh	o->1	
op.De	t->1	
op.In	r->1	
op.Ja	g->1	
op.So	m->1	
opa -	 ->2	
opa a	l->2	t->5	v->1	
opa b	e->1	
opa d	ä->1	
opa e	f->1	n->3	
opa f	i->1	o->1	å->1	ö->3	
opa h	a->11	
opa i	 ->6	n->3	
opa k	a->5	o->3	u->1	v->1	
opa m	e->8	å->4	ö->1	
opa n	ä->1	
opa o	c->18	s->1	
opa p	å->3	
opa r	e->2	
opa s	k->4	n->1	o->19	p->1	å->1	
opa t	a->1	r->1	y->2	
opa u	n->2	r->1	t->1	
opa v	a->1	e->1	i->4	ä->1	
opa ä	r->11	
opa!A	v->1	
opa!F	r->1	
opa".	J->1	
opa, 	K->1	S->1	b->1	d->5	e->3	f->1	h->1	i->1	n->1	o->11	s->4	t->1	v->3	ä->2	
opa..	 ->1	(->1	
opa.1	8->1	
opa.D	e->15	
opa.E	n->1	t->1	
opa.F	r->2	ö->1	
opa.H	e->6	
opa.I	 ->2	
opa.J	a->8	
opa.M	a->1	e->1	å->1	
opa.N	ä->1	
opa.O	c->1	
opa.P	r->1	
opa.R	e->1	
opa.T	r->1	y->1	
opa.U	n->1	
opa.V	a->1	i->9	
opa.Ä	v->1	
opa; 	e->1	
opa?H	e->1	
opa?V	a->1	i->1	
opaNä	s->1	
opade	m->2	
opaga	n->3	
opage	r->1	
opagr	u->1	
opako	n->1	
opami	n->1	
opani	v->1	
opapa	r->166	
opar 	e->1	i->1	p->1	
opart	i->2	
oparå	d->1	
opas 	b->2	c->1	d->2	e->2	f->8	g->1	h->2	k->2	l->1	m->8	n->2	o->1	p->1	r->1	s->9	t->2	u->1	v->2	
opatj	ä->1	
opava	l->3	
opeis	e->2	k->710	
opera	h->1	t->11	
opere	r->1	
opet 	p->2	
opia 	t->1	
opien	 ->1	,->2	
opier	a->1	
opilo	t->1	
opini	o->4	
oplas	t->1	
opol 	a->2	i->2	m->2	o->6	s->2	t->1	
opol,	 ->3	
opol.	E->1	H->1	
opol;	 ->1	
opola	v->1	
opolf	r->1	ö->2	
opoli	n->1	s->2	
opolk	o->1	
opols	 ->3	i->1	
oport	i->9	
opoul	o->5	
opp -	 ->1	
opp a	n->1	v->1	
opp f	r->1	ö->7	
opp h	a->2	
opp i	 ->1	
opp p	å->1	
opp s	o->1	
opp, 	o->1	
opp..	(->1	
oppa 	a->1	i->2	t->1	ö->1	
oppad	e->2	
oppar	 ->1	
oppas	 ->95	,->4	
oppe 	i->1	
oppen	 ->7	.->1	
oppet	 ->8	,->2	
oppla	 ->1	d->1	s->2	
oppli	n->2	
opplö	s->1	
oppmö	t->12	
oppni	n->12	
oppon	e->3	
oppor	t->2	
oppos	i->2	
oprak	t->1	
oprog	r->2	
oproj	e->1	
oprop	o->2	
oprot	o->2	
optim	a->3	i->4	
optio	n->1	
opula	r->1	
opuli	s->4	
opulä	r->2	
opyri	g->1	
opå b	a->1	
opé o	c->1	
opéer	 ->4	,->2	n->3	
or - 	d->1	l->1	n->1	
or Fr	a->1	
or Mo	n->2	
or Te	s->1	
or Ts	a->2	
or al	l->1	
or an	d->1	g->1	s->1	
or ar	b->1	
or at	t->85	
or av	 ->9	s->1	
or be	h->1	s->4	t->9	
or bi	l->2	
or bl	o->1	
or bo	r->1	
or br	i->2	
or bö	r->3	
or ch	o->1	
or de	 ->5	l->10	r->1	s->1	t->4	
or dj	u->1	
or dä	r->7	
or dö	d->1	l->1	
or ef	t->2	
or eg	e->1	
or el	l->4	
or en	 ->1	e->1	h->1	
or er	k->1	
or eu	r->1	
or fa	k->2	r->1	s->1	
or fi	c->1	
or fo	r->2	
or fr	a->1	i->1	å->5	
or fö	r->27	
or ga	g->1	
or ge	m->1	n->1	t->1	
or gr	å->1	
or gä	l->1	
or gö	r->1	
or ha	 ->1	d->1	n->1	r->9	
or hi	n->1	
or hj	ä->3	
or hä	n->2	
or hö	g->1	
or i 	B->1	D->1	E->2	F->1	I->1	K->1	P->1	S->1	a->1	d->4	e->3	f->1	g->1	j->1	m->1	r->1	s->5	t->1	u->1	v->1	
or in	d->1	f->1	l->1	n->2	o->5	s->1	t->17	v->1	
or ja	g->23	
or jo	r->2	
or ju	 ->1	
or ka	n->3	t->2	
or ko	m->1	s->1	
or le	v->1	
or li	v->2	
or lö	p->1	
or ma	j->4	n->1	r->1	s->1	
or me	d->8	l->1	n->1	r->2	
or mi	g->1	
or my	c->1	
or mä	n->2	
or må	n->2	s->2	
or ni	 ->4	
or no	g->1	
or nä	r->1	
or oc	h->65	k->5	
or om	 ->15	s->1	
or or	o->2	
or pe	r->1	
or po	l->2	
or pr	ö->1	
or på	 ->20	
or re	f->2	g->1	s->2	
or ro	l->1	
or sa	d->1	m->1	
or se	d->2	n->1	
or sj	ä->1	
or sk	a->3	y->1	
or so	m->94	
or st	ä->1	ö->1	
or sy	m->1	
or så	 ->1	l->1	s->1	
or ti	l->24	
or tj	ä->1	
or tr	ä->1	
or un	d->1	
or up	p->8	
or ur	 ->1	
or ut	a->2	f->1	g->1	m->2	s->6	t->1	v->1	
or va	d->1	k->1	r->3	
or ve	t->2	
or vi	 ->6	d->1	k->3	l->2	
or vä	c->1	g->1	
or än	 ->1	d->2	
or är	 ->10	l->1	
or äv	e->1	
or öv	e->2	
or) o	c->1	
or, a	t->1	
or, b	l->2	
or, e	l->1	n->2	
or, f	r->2	ö->1	
or, g	a->1	ö->1	
or, h	e->1	
or, i	 ->1	n->5	
or, k	a->2	o->1	
or, m	e->10	ä->3	
or, n	y->1	ä->1	
or, o	c->9	m->1	r->1	
or, p	e->1	
or, r	e->1	ä->1	
or, s	a->3	i->1	j->1	o->10	t->1	ä->2	å->2	
or, t	i->2	
or, u	t->5	
or, v	i->2	
or, ä	r->1	v->3	
or. D	e->1	
or..(	E->1	
or.Al	l->1	
or.Br	e->1	
or.De	 ->2	n->7	t->14	
or.Dä	r->1	
or.Et	t->1	
or.Fe	m->1	
or.Fr	u->2	å->1	
or.Fö	r->6	
or.Ge	n->1	
or.He	r->2	
or.Hu	v->1	
or.Ja	c->1	g->11	
or.Ka	n->1	
or.Ko	m->2	
or.Li	k->1	
or.Ma	n->1	
or.Me	d->1	n->1	
or.My	l->1	
or.Na	t->1	
or.Ny	a->1	
or.Nä	r->1	
or.Oc	h->2	
or.Re	f->1	
or.Sa	m->2	
or.Ti	l->1	
or.Ty	v->1	
or.Ve	m->1	
or.Vi	 ->5	s->1	
or.Vå	r->1	
or.Äv	e->1	
or.ÖV	P->1	
or: d	e->1	
or: f	ö->1	
or: o	m->1	
or: t	i->1	
or; j	a->1	
or?, 	r->1	
or?Ha	r->1	
or?Hu	r->1	
or?Är	 ->1	
ora 1	6->1	
ora a	k->1	l->1	m->1	n->2	r->3	v->1	
ora b	e->5	y->1	
ora d	e->3	r->2	
ora e	k->2	n->1	u->2	
ora f	r->3	ö->44	
ora g	e->1	r->6	
ora h	e->1	i->1	
ora i	 ->1	n->7	
ora k	a->1	e->1	o->1	
ora m	i->1	ä->2	ö->1	
ora n	ä->1	
ora o	c->5	l->3	m->1	r->2	
ora p	e->2	o->1	r->10	
ora r	e->1	i->2	
ora s	a->1	i->1	k->4	o->2	p->1	t->1	u->3	v->4	y->1	
ora t	e->1	i->1	o->1	r->2	
ora u	t->3	
ora v	a->1	i->1	ä->1	å->1	
ora å	r->1	t->2	
ora, 	o->1	v->1	
ora.E	n->1	
ora.M	e->1	
ora.V	a->1	
ora?A	n->1	
orad 	e->1	u->1	
orade	 ->2	.->1	
oral 	s->1	
oral,	 ->1	
orale	n->1	
orali	s->5	
orand	e->1	
orar 	a->1	d->1	e->1	v->1	
orat 	-->1	a->1	e->1	f->1	m->2	v->1	
orat,	 ->3	
orat.	D->1	H->1	
orate	n->1	t->12	
orati	n->4	
orato	r->3	
orats	 ->1	
orber	a->1	
orbet	t->1	
orbih	a->1	
orbri	t->14	
orbro	t->1	
orce 	b->1	
orcyk	l->4	
ord -	 ->1	
ord I	n->2	
ord a	n->1	t->2	v->1	
ord b	l->1	
ord e	f->1	
ord f	ö->6	
ord i	 ->4	n->2	
ord j	a->1	
ord k	o->1	r->1	u->1	
ord m	e->1	
ord n	ä->1	
ord o	c->8	m->3	
ord s	o->6	
ord t	a->1	e->1	i->2	
ord v	a->1	i->2	
ord, 	m->1	o->2	s->1	
ord-f	ö->1	
ord.B	e->1	
ord.E	u->1	
ord.U	n->1	
ord.V	i->2	
ord: 	"->2	
orda 	e->1	p->1	r->1	u->1	v->1	
orda,	 ->1	
ordad	.->1	
ordal	a->4	y->2	
ordam	e->4	
ordan	d->1	i->1	s->1	
ordar	 ->2	
ordbr	u->56	ä->1	
ordbä	v->10	
orde 	a->2	b->5	d->9	e->5	f->6	g->2	h->9	i->11	j->1	k->8	m->5	n->2	o->1	p->1	r->6	s->5	t->4	u->5	v->13	
orde,	 ->1	
orde.	D->1	N->1	
ordea	u->1	
orden	 ->3	.->1	s->2	t->25	
order	l->5	n->1	
ordes	 ->5	
ordet	 ->20	.->2	
ordeu	r->1	
ordfö	r->216	
ordin	ä->1	
ordir	l->2	
ordis	k->4	
ordit	a->1	
ordku	s->1	
ordla	d->1	
ordli	g->4	s->1	
ordmå	n->1	
ordna	 ->7	d->9	n->2	r->5	s->2	t->3	
ordni	n->155	
ordon	 ->32	,->8	.->9	?->1	N->1	e->7	s->7	
ordra	 ->3	n->7	r->2	s->5	t->1	
ordre	 ->1	
ordri	f->2	k->2	n->1	
ordsk	a->1	
ordsu	t->1	
ordti	d->1	
ordty	s->1	
ordvr	ä->1	
ordvä	n->1	s->1	
ore b	r->1	ä->1	
ore d	e->5	
ore e	n->3	t->2	x->1	
ore f	a->2	ö->1	
ore h	e->1	
ore i	 ->1	n->1	t->1	
ore l	ä->1	
ore m	e->2	
ore o	l->1	m->1	r->1	
ore p	a->1	
ore t	i->1	
ore v	a->1	
ore ö	n->1	
orea 	b->1	o->2	
oreal	i->2	
orebo	a->1	
oredl	i->1	
oregl	e->1	
orela	t->1	
oren 	e->2	f->7	i->1	k->2	o->3	p->1	t->1	
oren,	 ->1	
oren.	D->1	E->1	J->1	V->1	
orena	 ->1	n->5	r->12	s->1	
oreni	n->9	
orenz	 ->12	)->2	,->3	F->1	b->1	
orer 	-->1	a->3	d->1	f->1	g->1	i->3	o->3	s->14	u->1	ä->2	
orer,	 ->2	
orer.	D->1	J->1	T->1	V->1	
orera	 ->3	s->1	
orern	a->10	
orest	i->1	
oret 	f->1	
oreti	s->2	
orför	e->2	
org a	v->1	
org o	c->1	m->6	
org s	a->1	
org t	i->1	
organ	 ->15	"->1	,->6	.->1	e->9	i->61	
orgar	 ->1	d->1	e->71	n->88	s->7	
orge 	o->1	
orge,	 ->1	
orger	l->3	
orgli	g->3	
orgmä	s->2	
orgon	 ->27	,->2	.->6	d->2	
orgsf	u->1	
orhav	e->1	
orhet	s->1	
ori 8	 ->2	
ori o	c->2	
ori s	k->1	
ori v	a->1	
oria 	-->1	f->1	i->1	o->2	s->1	
oria,	 ->2	
oria.	D->1	Ä->1	
oriel	l->5	
orien	 ->5	s->2	t->6	
orier	 ->4	,->1	.->3	n->2	
oriet	"->1	,->2	
origi	n->2	
orik 	n->1	
orik,	 ->1	
orik.	F->1	
orike	r->1	
orikt	i->3	
oriml	i->5	
orind	u->2	
oring	 ->1	
orino	 ->3	,->1	.->2	s->1	
oris 	P->1	
orise	r->2	
orisk	 ->8	,->1	.->1	a->17	e->1	t->7	
orism	.->2	
oriso	n->3	
orist	a->1	e->6	h->1	
orita	s->1	
orite	r->32	t->72	
oritl	e->1	
orium	 ->2	,->3	.->5	
ork v	i->1	
orka,	 ->1	
orkan	 ->1	e->2	
orkap	i->1	
orkni	n->1	
orld 	W->1	
orlig	e->2	
orlun	d->3	
orlär	l->1	
orm a	t->2	v->24	
orm b	e->1	
orm d	a->1	ö->1	
orm e	l->1	
orm f	ö->3	
orm i	 ->3	
orm j	u->1	
orm k	a->1	o->3	
orm l	ö->1	
orm o	c->3	
orm p	å->1	
orm s	k->2	o->4	p->1	
orm v	i->2	ä->1	
orm ä	r->1	
orm ö	v->1	
orm, 	e->2	f->1	m->1	o->2	s->1	u->1	ä->1	
orm.D	e->1	
orm.E	G->1	
orm.M	e->1	
orm.N	u->1	
orm.S	a->1	
orm.V	i->1	
orm.Ä	r->1	
orm: 	e->1	
orma 	M->1	b->3	d->3	e->1	f->2	k->3	m->3	p->1	s->5	u->1	ö->1	
orma.	O->1	
ormad	e->1	
ormal	a->2	i->4	t->5	
orman	d->4	s->1	
ormar	 ->7	b->3	n->13	
ormas	 ->3	
ormat	 ->2	i->74	s->1	
ormel	l->16	
ormen	 ->13	,->2	.->3	s->5	
ormer	 ->55	,->3	.->12	a->26	i->17	n->18	
ormfä	l->1	
ormfö	r->2	
ormis	t->1	
ormni	n->26	
ormon	b->1	
ormpa	k->1	
ormpr	o->14	
ormst	ä->1	
ormt 	a->2	e->1	h->1	m->1	u->1	v->1	
ormul	e->18	
ormåt	g->1	
orn -	 ->2	
orn b	ö->1	
orn e	l->1	n->1	
orn f	i->1	o->1	ö->1	
orn i	 ->2	
orn k	a->1	
orn o	c->5	
orn s	a->1	t->1	ä->1	
orn u	n->1	
orn ä	r->2	
orn).	D->1	
orn, 	a->1	e->1	f->1	i->3	m->1	o->2	s->2	v->1	
orn.D	e->4	
orn.F	ö->3	
orn.H	e->1	
orn.K	o->1	
orn.M	i->1	
orn?A	n->1	
orna 	3->1	d->5	f->8	h->1	i->12	k->2	l->1	m->6	n->1	o->10	p->4	s->7	t->3	u->1	v->3	ä->4	
orna,	 ->10	
orna.	D->5	I->1	K->1	M->1	N->1	S->1	V->2	
orna?	E->1	
ornas	 ->7	
ornet	.->1	
ornog	r->2	
orns 	a->1	p->1	s->2	
oro -	 ->1	
oro E	u->1	
oro b	l->1	
oro d	i->1	
oro f	u->1	ö->4	
oro i	 ->3	
oro l	e->1	
oro n	ä->2	
oro o	c->3	m->1	
oro p	å->1	
oro s	o->12	
oro ä	r->2	v->1	
oro ö	v->1	
oro, 	d->1	f->1	s->1	ä->1	
oro.A	t->1	
oro.B	e->1	
oro.F	l->1	ö->1	
oro.J	a->2	
oro.O	m->1	
oro.T	r->1	
oro.V	i->1	
oroa 	f->1	o->1	s->1	
oroad	 ->3	e->2	
oroan	d->9	
oroar	 ->4	
oroli	g->6	
oron 	-->1	f->2	ä->1	ö->1	
orosm	o->4	
orovä	c->2	
orpet	 ->2	
orpol	i->1	
orpus	 ->5	
orr?V	i->1	
orra 	T->1	d->2	o->1	
orrai	n->2	
orrec	t->1	
orrek	t->27	
orren	 ->1	
orres	p->1	
orrey	 ->3	
orrid	o->2	
orrum	p->2	
orrup	t->7	
ors a	r->1	
ors b	e->1	r->1	y->1	
ors d	e->5	ö->1	
ors e	n->1	
ors f	r->3	ö->2	
ors g	o->1	
ors h	a->4	ä->3	
ors i	 ->4	n->3	
ors k	o->2	
ors l	e->1	i->1	
ors o	c->4	
ors p	l->1	
ors r	ä->2	
ors s	i->1	o->2	ä->2	å->1	
ors t	i->2	o->1	
ors u	t->1	
ors y	r->1	
ors ö	k->1	
ors, 	a->1	m->1	o->2	p->1	s->1	ä->1	
ors.D	e->5	
ors.J	a->1	
ors.M	e->1	
ors.T	y->1	
ors.U	t->1	
ors.V	i->2	
orsak	 ->1	.->2	a->18	e->15	
orsan	a->1	
orsbe	s->1	
orsda	g->8	
orse 	f->1	o->1	s->1	
orse,	 ->1	
orse.	D->1	V->1	
orsel	!->1	
orsin	r->1	
orska	l->2	r->5	s->1	
orskn	i->35	
orskr	o->1	
orsla	g->2	
orsli	n->1	
orst 	c->1	
orstä	d->2	
orsöv	e->1	
ort -	 ->1	
ort E	G->1	
ort a	l->1	n->12	t->4	v->25	
ort b	e->1	i->1	l->1	ä->1	ö->2	
ort d	e->13	ä->1	
ort e	g->1	n->4	r->1	t->8	x->1	
ort f	i->2	r->5	ö->14	
ort g	e->2	r->1	å->2	
ort h	a->4	i->1	ä->1	å->1	
ort i	 ->4	f->1	n->8	
ort k	a->1	l->1	n->1	o->1	r->2	u->1	
ort l	ä->2	
ort m	e->4	o->1	å->2	
ort n	e->1	ä->1	å->6	
ort o	c->24	l->1	m->10	
ort p	e->2	r->1	å->6	
ort r	e->3	i->1	
ort s	a->5	e->5	i->9	k->3	o->6	t->3	v->1	ä->3	å->2	
ort t	a->6	i->3	y->1	
ort u	n->2	p->1	t->3	
ort v	e->1	i->5	ä->1	
ort ä	r->2	
ort å	t->1	
ort ö	v->2	
ort) 	t->1	
ort, 	b->1	d->2	e->2	g->2	h->2	i->1	k->2	m->3	n->1	o->3	p->1	s->1	t->1	v->2	ä->2	
ort- 	o->1	
ort-s	t->2	
ort.D	e->6	i->1	å->1	
ort.E	n->1	
ort.I	 ->1	
ort.J	a->2	u->1	
ort.L	å->1	
ort.N	i->1	
ort.R	i->1	
ort.S	a->1	
ort.U	t->1	
ort.V	i->3	
ort: 	E->1	
ort?J	a->1	
ortNä	s->1	
orta 	f->3	o->1	t->1	
ortab	l->1	
ortad	e->1	
ortam	e->1	
ortas	t->1	
ortbe	s->2	
ortbi	l->1	
ortdi	r->1	
orten	 ->36	,->3	.->5	:->1	s->3	
orter	 ->20	,->5	.->7	a->22	i->1	n->9	
ortet	 ->15	.->1	s->3	
ortfa	l->6	r->89	t->2	
ortfe	d->1	
ortfr	å->1	
ortfö	r->1	
ortgr	u->1	
ortgå	.->2	e->3	
ortio	n->9	
ortko	s->2	
ortle	v->1	
ortma	r->1	
ortmo	n->1	
ortni	n->1	
ortnä	t->1	
ortom	 ->3	r->3	
orton	 ->8	d->1	
ortpr	i->1	o->1	
orts 	"->1	a->6	c->1	d->1	e->2	f->4	h->2	i->2	m->1	n->1	o->2	u->1	v->1	
orts,	 ->3	
orts.	J->2	
ortsa	t->12	
ortse	 ->4	r->1	t->1	
ortsi	f->1	k->4	
ortsk	r->1	
ortsä	k->7	t->82	
ortug	a->26	i->70	u->1	
ortun	i->2	
ortut	s->1	
ortvi	n->1	
ortyr	e->1	
orum 	f->1	h->1	i->1	o->1	
orum,	 ->1	
orume	t->1	
orv f	å->1	
orven	 ->3	.->2	
orwel	l->1	
oräkn	e->1	
orär 	o->1	
orärt	 ->1	
orätt	 ->1	v->9	
orêts	 ->1	
orös 	r->1	
orösa	 ->2	
oröst	 ->1	
os Da	m->1	
os EG	-->1	
os Eu	r->1	
os FP	Ö->1	
os Oz	,->1	
os RE	P->1	
os al	b->1	l->2	
os an	f->1	
os at	t->1	
os av	d->1	
os be	f->1	g->1	t->9	
os bl	a->1	
os de	 ->4	f->1	m->3	n->2	t->3	
os en	 ->1	d->1	e->1	
os ex	t->1	
os fa	r->1	
os fö	r->5	
os ha	r->1	
os in	b->1	s->1	t->1	
os kl	i->1	
os ko	m->6	
os le	d->1	
os me	d->3	
os mi	n->1	
os mä	n->1	
os må	n->1	
os nä	r->1	
os oc	h->8	
os or	d->3	
os os	s->3	
os pr	o->2	
os rå	d->1	
os se	r->1	
os si	n->2	
os st	ö->1	
os ta	l->1	
os ti	l->1	
os vu	x->1	
os vä	p->1	
os vå	r->1	
os yt	t->1	
os ås	i->1	
os! J	a->1	
os, a	t->1	
os, h	a->1	
os, k	a->1	
osamt	 ->2	
osann	o->1	
osats	e->1	
osatt	a->3	
osedd	a->1	
osenr	ö->1	
osexu	e->1	
osfär	e->1	
osion	e->1	
ositi	o->13	v->74	
osiv 	b->1	
osju 	i->1	
oskep	t->3	
oskop	,->3	
oskri	v->1	
oskva	,->1	
oskyd	d->1	
oslav	i->1	
osläk	t->1	
osmol	n->1	
osmom	e->3	
osnie	r->2	
osofi	 ->2	,->1	n->1	s->1	
osor,	 ->1	
osovo	 ->25	,->11	.->12	?->2	N->1	k->2	s->7	
ospic	e->1	
ospin	 ->1	
oss -	 ->1	
oss a	l->6	n->4	t->27	v->2	
oss b	e->1	
oss d	e->10	o->1	ä->6	å->2	
oss e	m->2	n->9	t->4	u->1	
oss f	r->4	ö->12	
oss g	e->3	ä->1	
oss h	a->3	o->1	u->1	ä->1	
oss i	 ->21	d->1	n->7	
oss k	a->1	o->2	
oss l	e->1	u->1	å->1	
oss m	e->8	o->1	y->2	å->1	
oss n	e->2	y->1	ä->2	å->1	
oss o	a->1	c->11	d->1	f->1	m->15	
oss p	a->1	o->1	å->11	
oss r	a->1	ä->1	
oss s	a->2	e->1	i->2	j->9	l->2	o->8	t->1	ä->1	å->3	
oss t	a->1	i->13	r->2	
oss u	n->4	p->1	t->3	
oss v	a->7	e->3	i->2	ä->1	
oss y	t->1	
oss ä	n->2	r->8	
oss å	t->10	
oss ö	v->3	
oss, 	T->1	a->1	f->2	g->1	h->1	m->3	o->2	s->1	v->2	ä->1	
oss.D	e->3	
oss.E	n->1	u->1	
oss.F	r->2	
oss.H	e->1	
oss.J	a->4	
oss.N	å->1	
oss.V	a->1	i->2	
oss.Ä	v->2	
oss: 	k->1	
oss?.	 ->1	
oss?V	i->1	
ossal	a->1	
ossar	 ->1	
osset	ê->2	
ossil	 ->1	a->2	
ossni	n->1	
osstê	t->1	
ost a	v->1	
ost f	ö->2	
ost o	c->1	
ost t	i->1	
ost u	t->1	
ost v	i->1	
ost-b	e->5	
ost.N	ä->1	
osta 	h->1	k->1	n->1	o->1	s->2	v->2	ä->1	
osta,	 ->2	
ostad	e->2	i->1	s->1	
ostar	 ->4	
ostas	i->1	
ostat	 ->2	e->1	
ostbi	l->1	
osten	 ->1	
oster	 ->3	.->2	n->1	
osteu	r->1	
osthå	l->1	
ostit	u->1	
ostna	d->108	
ostra	t->2	
ostro	n->3	
ostsa	m->2	
ostve	r->1	
ostäd	e->4	
osv. 	M->1	V->1	m->1	
osv.,	 ->1	
osv.?	A->1	
osv.S	v->1	
osynl	i->1	
osyst	e->4	
osäke	r->12	
osätt	a->2	n->3	
osårb	a->1	
ot - 	s->1	v->1	
ot -e	r->1	
ot 13	 ->1	
ot 5 	0->1	
ot Ai	d->1	
ot Da	n->1	
ot EG	-->1	
ot EU	 ->1	:->1	
ot Eu	r->7	
ot Fr	a->1	
ot Fö	r->2	
ot Gr	e->1	
ot Ha	d->1	i->2	
ot Is	r->1	
ot Jo	n->3	
ot Ka	r->1	
ot La	n->1	
ot Mo	n->1	
ot Ra	p->2	
ot So	u->1	
ot Ti	b->1	
ot To	d->1	
ot UN	M->1	
ot Wa	l->1	
ot Wu	l->1	
ot ab	s->1	
ot ai	d->1	
ot al	l->7	
ot an	n->5	s->3	t->1	v->1	
ot ar	b->2	
ot at	t->16	
ot av	 ->17	f->1	g->1	s->1	
ot ba	k->17	n->1	
ot be	d->2	s->1	t->3	
ot br	o->1	å->1	
ot bä	t->1	
ot bå	d->1	
ot de	 ->9	m->2	n->29	r->1	s->2	t->17	
ot di	r->2	s->2	
ot do	k->1	l->2	
ot ek	o->1	
ot el	l->1	
ot en	 ->13	
ot er	,->1	a->1	k->1	
ot et	t->7	
ot ex	c->1	e->1	t->2	
ot fe	l->1	
ot fo	r->2	
ot fr	a->1	e->1	u->1	ä->2	å->5	
ot fö	r->17	
ot ge	m->1	
ot gl	o->1	
ot ha	r->4	
ot he	l->1	
ot hi	n->1	
ot hu	m->1	r->1	
ot hä	l->1	r->1	
ot i 	d->2	f->1	k->1	s->2	u->1	
ot id	é->1	
ot in	 ->1	f->1	s->1	t->4	v->1	
ot ja	g->4	
ot ka	n->1	
ot kl	a->1	
ot ko	m->4	n->2	r->1	
ot kö	n->1	
ot la	n->1	
ot le	k->1	
ot li	k->1	
ot lo	j->1	
ot ly	s->1	
ot lä	g->1	m->2	
ot ma	r->3	s->1	
ot me	d->5	r->3	
ot mi	n->2	
ot mo	t->6	
ot my	c->4	
ot mä	n->1	r->1	
ot må	l->1	
ot na	r->1	t->1	z->1	
ot nä	r->1	s->1	t->1	
ot nå	g->1	
ot oc	h->1	
ot oe	g->1	
ot ok	l->1	
ot ol	i->1	j->1	y->1	
ot om	 ->8	.->1	
ot os	s->3	
ot pa	r->1	t->1	
ot pe	s->1	
ot po	l->2	t->1	
ot pr	e->1	i->3	o->1	
ot pu	n->1	
ot på	 ->4	
ot ra	d->1	s->1	
ot re	g->2	s->3	
ot rå	d->4	
ot sa	m->1	
ot se	r->1	
ot si	g->1	n->2	
ot sj	ö->1	
ot sk	a->2	e->1	i->1	u->2	
ot sl	a->3	u->2	
ot sn	a->1	
ot so	c->2	m->53	
ot sp	e->2	o->1	
ot st	a->1	i->1	r->2	y->1	ä->1	ö->2	
ot su	v->2	
ot sv	a->2	å->1	
ot sy	s->1	
ot sä	k->1	t->11	
ot så	d->3	
ot ta	b->1	l->1	n->1	
ot te	x->1	
ot ti	d->1	l->2	
ot tv	i->1	
ot un	i->2	
ot up	p->2	
ot ut	ö->1	
ot va	d->1	l->1	r->4	
ot ve	d->1	r->2	t->2	
ot vi	 ->2	d->2	l->1	s->6	
ot vä	l->1	
ot vå	r->4	
ot yt	t->1	
ot Ös	t->3	
ot än	d->1	
ot är	 ->2	
ot år	,->1	
ot åt	g->1	
ot ök	a->1	n->1	
ot öv	e->3	r->1	
ot! D	e->2	
ot! J	a->2	
ot! N	ä->1	
ot! S	o->1	
ot! V	a->1	
ot!De	t->1	
ot, Z	i->1	
ot, a	t->5	
ot, d	e->1	
ot, e	f->2	
ot, h	ä->2	
ot, o	c->1	
ot, s	i->1	o->1	
ot, t	r->1	
ot, u	p->1	
ot, v	i->1	
ot, ä	r->2	v->1	
ot. 7	 ->1	
ot.Al	l->1	
ot.De	t->2	
ot.Fr	u->2	
ot.Ja	g->2	
ot.Sl	u->1	
ot.Vi	 ->1	
ot.Än	d->1	
ot?Ne	j->1	
ota d	e->1	
ota f	ö->1	
ota h	o->1	
ota k	a->1	
otack	s->1	
otad.	M->2	
otade	 ->4	.->1	s->1	
otal 	b->1	m->1	o->1	t->1	
otal,	 ->1	
otal-	F->3	
otalF	i->1	
otala	 ->12	n->2	
otalb	e->1	l->1	
otale	t->1	
otalf	å->4	ö->1	
otali	t->2	
otals	 ->5	u->1	
otalt	 ->6	
otalv	o->1	
otan;	 ->1	
otand	e->1	
otar 	b->1	d->2	e->2	h->1	j->1	m->2	v->1	
otarb	e->1	
otas 	e->2	m->1	n->1	o->1	u->1	v->2	
otas.	V->1	
otat 	d->1	
otati	o->1	
otbil	d->1	
otbol	l->1	
ote Q	u->1	
oteke	n->2	
otekt	i->4	
otels	e->1	
oten 	A->2	B->1	L->1	R->1	a->3	f->3	h->3	i->2	k->1	m->2	o->1	s->2	t->3	
oten.	D->2	J->1	
otens	 ->2	
otent	i->6	
oter 	s->1	
oter.	 ->1	
otera	 ->6	d->3	r->9	s->1	t->8	
oteri	n->5	
otern	a->4	
otese	n->1	
otest	 ->2	,->1	a->2	e->4	
otet 	k->1	m->3	o->3	
oteti	s->1	
otful	l->1	
otfär	d->1	
otfäs	t->1	
otgån	g->1	
oth-B	e->7	
othar	 ->2	"->1	
other	"->1	
otika	 ->2	b->1	f->1	n->1	p->1	s->1	
otill	f->2	r->12	å->3	
otion	e->1	
otis 	d->1	
otisk	a->1	
otism	 ->2	.->3	
otiv 	i->1	t->1	
otiva	t->1	
otive	n->2	r->16	
otjän	s->1	
otnin	g->17	
oto k	a->1	
oto o	c->1	
oto-p	r->1	
oto.V	i->1	
otoko	l->26	
otopr	o->2	
otor 	o->1	
otor.	A->1	R->1	
otorc	y->4	
otori	n->2	
otos 	k->1	
otpar	t->4	
otpro	g->1	j->1	
otrol	i->2	
otryg	g->1	
ots a	l->13	t->21	
ots d	e->20	
ots e	n->1	
ots i	n->1	
ots k	a->1	
ots m	i->1	
ots p	r->1	
ots r	å->1	
ots s	o->1	v->1	
ots t	i->1	
ots v	i->1	
otsat	s->16	t->7	
otspå	r->2	
otstr	ä->1	
otsty	c->3	
otstå	n->10	r->2	
otsva	r->17	
otsys	t->1	
otsäg	a->1	e->7	
otsät	t->9	
ott a	n->2	r->1	t->1	v->1	
ott b	e->2	o->1	
ott d	e->1	i->1	
ott e	f->1	n->1	x->1	
ott f	r->1	ö->4	
ott h	e->1	u->1	
ott i	 ->3	n->1	
ott m	o->4	
ott n	y->3	
ott o	c->5	
ott p	å->3	
ott r	e->2	
ott s	a->1	k->1	o->6	t->1	y->2	
ott u	n->1	
ott ä	r->1	
ott, 	a->1	b->1	f->2	g->1	k->2	t->3	v->1	
ott.D	e->2	
ott.F	ö->1	
ott.I	 ->1	
ott.J	a->1	
ott.L	å->1	
ott.M	o->1	
ott.O	b->1	m->1	r->1	
ott.Ä	v->1	
otta 	o->1	t->1	
otta,	 ->1	
ottad	e->3	
ottag	a->11	i->3	n->2	
ottan	.->1	
ottar	 ->1	
ottas	 ->1	
ottat	s->2	
otten	 ->6	,->1	l->1	
otter	d->2	i->1	
ottet	 ->113	,->5	.->11	s->7	
ottgö	r->1	
otti 	g->1	
ottla	n->5	
ottmå	l->1	
ottna	r->3	
ottne	n->1	
ottor	n->1	
otts 	b->1	f->1	k->1	
ottsb	e->5	
ottsd	e->1	
ottsf	r->1	
ottsl	i->17	
ottsm	y->1	å->1	
ottso	f->2	
ottsp	a->1	
ottsr	u->1	
otull	a->1	
otum 	f->1	
oturi	s->1	
otuse	n->1	
otver	k->4	
otvet	y->2	
otvik	t->1	
otvil	l->1	
otviv	e->1	
otydl	i->4	
otänk	b->1	
otåli	g->1	
otåtg	ä->3	
ou fr	å->1	
ou oc	h->1	
ouchn	e->12	
ouk a	l->1	
oulad	a->1	
oulos	 ->5	
oumbä	r->4	
ounci	l->1	
oundg	ä->2	
oundv	i->4	
oup ,	 ->1	
oup d	e->1	
oura 	f->3	o->1	s->2	
oura,	 ->2	
ourg 	m->1	ö->1	
ourg.	J->1	L->1	V->1	
ouri.	B->1	
ourla	n->6	
ourna	l->2	
ourne	r->1	
ours 	d->1	
ousew	i->1	
ousko	u->1	
outhä	r->2	
outie	r->1	
outny	t->1	
oux-a	f->1	
ov at	t->1	
ov av	 ->12	,->1	.->1	s->1	
ov fö	r->4	
ov i 	K->1	
ov in	t->1	
ov ko	m->1	
ov ny	s->1	
ov oc	h->6	k->1	
ov på	 ->9	
ov so	m->1	
ov sy	f->1	
ov så	 ->1	
ov ti	l->8	
ov", 	d->1	
ov, a	t->1	
ov, n	å->1	
ov, ä	r->1	
ov. D	e->1	
ov.Av	s->1	
ov.De	t->1	
ov.He	r->1	
ov.Up	p->1	
ova a	t->2	
ovade	 ->3	.->1	
ovaki	e->1	
ovan,	 ->1	
ovan.	T->1	
ovana	 ->1	
ovani	f->1	
ovanl	i->1	
ovann	ä->2	
ovanp	å->1	
ovans	 ->1	t->1	
ovar 	-->1	a->1	
ovat 	-->1	E->1	a->2	t->1	
ovat.	Å->1	
ovati	o->4	v->2	
ovats	.->1	
ovemb	e->11	
oven 	e->1	i->1	o->1	p->1	ä->1	
oven.	S->1	
ovens	k->1	
over 	i->1	
over,	 ->1	
overa	r->1	
overh	e->1	
overi	n->3	
overs	e->2	i->2	
ovet 	-->1	a->32	f->1	i->1	ä->1	
ovet,	 ->2	
ovic 	i->1	
ovilj	a->2	
ovill	k->2	
ovins	 ->2	e->1	
ovis 	s->1	
ovis)	 ->1	
ovisa	s->1	t->2	
ovisb	e->9	
ovise	n->1	
ovisf	i->3	
ovisk	v->2	
ovisn	i->1	
oviso	r->2	
oviss	h->1	
ovjet	t->1	
ovkar	t->1	
ovkon	s->1	
ovo (	K->2	
ovo T	r->1	
ovo a	t->1	
ovo b	ä->1	
ovo f	r->1	ö->2	
ovo h	a->1	
ovo i	n->1	
ovo k	a->1	ä->1	
ovo m	e->1	
ovo o	c->7	
ovo t	i->1	
ovo u	t->1	
ovo v	a->1	
ovo ä	r->3	
ovo, 	e->2	h->1	i->1	m->2	o->3	s->1	v->1	
ovo.-	 ->1	
ovo.A	v->1	
ovo.D	e->2	
ovo.E	u->1	
ovo.F	ö->1	
ovo.H	e->1	
ovo.K	o->1	
ovo.L	å->1	
ovo.M	e->1	
ovo.O	c->1	
ovo.V	i->1	
ovo? 	D->1	
ovo?H	u->1	
ovoNä	s->1	
ovoko	n->1	
ovokr	i->1	
ovord	a->2	
ovos 	a->1	d->1	e->1	l->1	m->1	s->1	y->1	
ovsid	a->1	
ovsko	n->2	
ovsma	n->2	
ovsmä	n->3	
ovste	s->1	
ovvär	d->2	
ovytt	r->1	
oväck	a->3	
oväde	r->1	
ovädr	e->1	
ovälk	o->1	
ovänl	i->1	
ovärd	i->15	
oväse	n->1	
ovådl	i->1	
ovård	 ->1	,->1	
ow ti	l->1	
ow-ho	w->1	
owe.E	u->1	
owe.V	i->1	
ower 	k->1	
ower,	 ->2	
owis 	h->1	n->1	
owitt	s->1	
own a	v->1	
own ä	r->1	
own, 	m->1	
ox oc	h->1	
ox sa	d->1	
ox!Ja	g->1	
ox, j	a->1	
ox, s	o->1	
oxal 	s->2	
oxala	 ->1	
oxalt	 ->2	
oxid 	i->1	o->3	
oxidu	t->1	
oxin 	o->1	
oxink	r->1	
oxisk	a->1	
oxnin	g->1	
oyal 	U->1	
oyds 	i->1	
oyola	 ->2	
oämne	n->1	
oändl	i->4	
oäng 	g->1	
oäng.	D->1	
oängs	y->2	
oängt	e->8	
oår f	ö->1	
oönsk	a->1	
oöver	l->1	s->5	
p (kr	i->2	
p , m	e->1	
p - o	c->2	
p - s	o->1	
p Cad	o->1	
p Eur	o->1	
p Jör	g->1	
p Tib	e->1	
p all	a->2	t->3	v->2	
p ans	e->2	v->1	
p ant	a->1	
p anv	ä->1	
p att	 ->11	
p av 	5->1	E->1	T->1	a->5	b->6	d->6	e->5	f->9	g->2	i->3	k->1	l->4	m->3	n->2	o->5	p->3	r->4	s->9	u->2	v->1	å->2	ö->1	
p avs	a->1	
p beg	ä->1	
p bet	a->1	r->1	
p bid	r->1	
p båd	e->1	
p bör	 ->2	
p de 	c->1	h->1	m->1	o->3	p->1	r->1	s->2	v->1	
p deb	a->2	
p dem	 ->2	
p den	 ->9	n->5	
p des	s->3	
p det	 ->7	.->1	:->1	t->3	
p dom	e->1	
p där	 ->3	
p eft	e->3	
p ell	e->3	
p en 	a->2	b->2	f->1	k->2	l->1	r->1	s->2	
p enl	i->1	
p ett	 ->6	
p exp	e->1	
p for	t->1	
p fra	m->2	
p frå	g->9	n->4	
p ful	l->1	
p fåt	t->1	
p för	 ->18	e->1	h->1	s->1	
p gen	o->2	
p gru	n->1	
p grä	n->1	
p had	e->1	
p har	 ->6	
p hel	a->1	
p huv	u->1	
p hän	d->2	
p här	 ->1	
p hög	e->1	
p i E	u->1	
p i S	v->1	
p i b	e->1	i->1	
p i d	a->1	e->5	
p i e	k->1	r->1	
p i f	ö->2	
p i h	a->1	
p i k	l->1	
p i m	a->1	i->2	
p i p	a->2	
p i r	e->1	å->2	
p i s	i->2	
p i t	a->1	i->1	
p i u	n->1	
p i v	å->2	
p i ä	g->1	
p idé	n->1	
p ige	n->4	
p inl	e->2	
p ino	m->2	
p int	e->6	
p kan	 ->1	
p kom	m->6	
p kon	f->1	
p lag	f->1	
p liv	s->1	
p läg	g->1	
p läm	n->1	
p län	g->1	
p man	 ->1	
p med	 ->7	.->1	
p mel	l->3	
p mot	 ->4	
p mås	t->2	
p nat	u->1	
p ni 	h->1	
p nya	 ->1	
p när	 ->1	
p någ	r->3	
p och	 ->23	
p olj	e->1	
p om 	d->4	i->1	m->1	s->1	v->1	
p ord	e->2	
p per	s->1	
p pos	i->1	
p pri	o->1	
p pro	b->2	
p på 	a->2	b->1	d->2	n->1	r->2	s->3	
p på.	J->1	V->1	
p ref	o->1	
p reg	i->1	
p räc	k->1	
p rät	t->2	
p råd	e->1	
p rös	t->1	
p sad	e->1	
p sig	 ->1	
p sin	a->1	
p sit	t->1	
p sjö	n->1	
p ska	l->4	p->1	
p sku	l->1	
p sky	d->1	
p som	 ->21	
p stä	l->2	
p sär	s->1	
p sät	t->1	
p såv	i->1	ä->1	
p til	l->18	
p tog	 ->1	
p tre	 ->1	
p två	 ->1	
p tyd	l->1	
p tyv	ä->1	
p und	e->3	
p upp	b->1	
p uta	n->2	
p utg	i->1	
p utt	a->2	j->1	
p utv	e->2	
p vad	 ->4	
p vid	 ->2	
p vil	l->2	
p väl	k->2	
p än 	e->1	
p änd	r->1	
p änn	u->1	
p är 	a->2	d->2	e->1	r->1	ä->1	ö->1	
p är,	 ->1	
p äre	n->2	
p äve	n->1	
p öns	k->1	
p öve	r->1	
p" fr	a->1	
p"!I 	d->1	
p", a	l->1	
p", v	i->1	
p, Ar	i->3	
p, ED	D->1	
p, an	s->1	
p, av	s->1	
p, bl	a->1	
p, de	 ->1	c->1	t->1	
p, dä	r->1	
p, då	 ->1	
p, ef	t->3	
p, en	 ->5	
p, fo	r->1	
p, få	r->1	
p, fö	r->1	
p, ge	 ->1	
p, ha	n->1	
p, he	r->2	
p, i 	b->1	
p, in	t->1	
p, ju	s->1	
p, li	k->1	
p, me	d->1	n->2	
p, mi	n->1	
p, nu	 ->1	
p, oc	h->6	
p, om	 ->1	
p, på	 ->1	
p, ri	k->1	
p, so	m->2	
p, sä	r->1	
p, ut	a->1	
p, va	r->1	
p, vi	l->2	
p, äv	e->1	
p-sho	p->1	
p. Sk	ä->1	
p. sä	k->1	
p. tr	a->1	
p..(F	R->1	
p.Ahe	r->1	
p.Dag	e->1	
p.De 	f->1	
p.Den	 ->2	
p.Det	 ->10	t->2	
p.Eft	e->1	
p.Eur	o->1	
p.Fak	t->1	
p.Här	 ->1	
p.I a	p->1	
p.I d	e->1	
p.I o	c->1	
p.Inr	e->1	
p.Jag	 ->12	
p.Men	 ->1	
p.På 	s->1	
p.Sjä	l->1	
p.Slu	t->1	
p.Som	 ->1	
p.Til	l->1	
p.Vi 	f->1	h->2	i->1	s->1	ö->1	
p.Vil	j->1	
p.Vis	s->1	
p.g.a	.->1	
p.Änd	å->1	
p.Äve	n->1	
p: Ko	n->1	
p?Hur	 ->1	
pa - 	d->1	k->1	m->1	
pa OL	A->1	
pa Wa	l->1	
pa al	l->3	
pa an	d->1	s->1	t->1	v->1	
pa ar	b->5	t->2	
pa at	t->7	
pa av	 ->1	
pa be	d->3	s->4	
pa bä	t->1	
pa da	t->1	
pa de	 ->5	m->5	n->6	s->2	t->9	
pa di	s->2	
pa dr	i->1	
pa dä	r->2	
pa ef	f->1	t->1	
pa ek	o->1	
pa el	l->1	
pa en	 ->26	e->1	i->1	l->1	
pa er	f->1	
pa et	t->14	
pa eu	r->2	
pa ex	t->2	
pa fi	n->1	
pa fl	e->2	
pa fo	r->2	
pa fr	e->2	ä->1	
pa få	 ->1	
pa fö	d->1	r->19	
pa ge	m->3	n->1	
pa gl	ö->1	
pa ha	d->1	r->10	
pa he	n->1	
pa ho	n->1	
pa hå	l->1	
pa hö	g->1	j->1	
pa i 	d->4	e->1	f->2	s->2	ö->1	
pa ih	o->1	
pa im	p->1	
pa in	 ->5	c->1	d->1	f->1	s->1	t->2	
pa jä	m->1	
pa ka	n->5	
pa kl	a->1	
pa ko	m->5	n->5	
pa kr	i->3	
pa ku	l->1	n->1	
pa kv	a->2	
pa la	n->1	
pa lu	g->1	
pa ma	r->1	
pa me	d->10	
pa mi	g->1	n->2	s->1	t->2	
pa mo	t->1	
pa mä	n->5	
pa må	s->4	
pa mö	d->1	t->1	
pa na	r->1	
pa ny	a->5	
pa nä	r->1	
pa nå	g->5	
pa oc	h->20	k->2	
pa of	f->2	
pa ol	i->1	
pa om	r->1	
pa or	i->1	
pa os	s->2	
pa pa	r->1	
pa pe	n->1	r->1	
pa pl	a->1	
pa po	l->1	
pa pr	i->2	
pa på	 ->4	
pa re	d->1	g->1	l->1	s->2	
pa rä	t->3	
pa si	n->2	
pa sk	a->5	i->1	
pa sn	a->2	
pa so	m->20	
pa sp	e->1	ä->1	
pa st	i->1	r->2	
pa su	b->1	
pa sy	m->1	s->5	
pa så	 ->2	s->1	
pa ta	g->2	r->1	
pa te	r->1	x->1	
pa ti	l->12	
pa tr	o->3	y->1	
pa tv	i->1	å->1	
pa ty	c->1	d->1	
pa un	d->2	g->1	i->1	
pa ur	 ->1	v->1	
pa ut	 ->1	a->1	
pa va	r->1	
pa ve	r->1	
pa vi	k->1	l->1	s->2	
pa vä	r->1	x->1	
pa vå	r->2	
pa yt	t->1	
pa än	n->1	
pa är	 ->11	
pa åt	e->1	
pa öv	e->1	
pa!Av	 ->1	
pa!Fr	u->1	
pa".J	u->1	
pa, K	v->1	
pa, S	c->1	
pa, b	l->1	
pa, d	e->3	v->1	ö->1	
pa, e	f->1	t->2	
pa, f	ö->1	
pa, h	a->1	
pa, i	 ->1	
pa, n	å->1	
pa, o	a->1	c->10	m->1	
pa, p	a->1	
pa, s	o->3	t->1	
pa, t	.->1	r->1	
pa, v	a->1	i->2	
pa, ä	r->2	
pa.. 	T->1	
pa..(	E->1	
pa.18	 ->1	
pa.De	n->3	s->1	t->11	
pa.Ef	t->1	
pa.En	 ->1	
pa.Et	t->1	
pa.Fr	u->2	
pa.Fö	r->1	
pa.He	r->6	
pa.I 	f->1	s->1	
pa.Ja	g->8	
pa.Ko	m->1	
pa.Ma	n->1	
pa.Me	n->1	
pa.Må	n->1	
pa.Nä	r->1	
pa.Oc	h->1	
pa.Pr	o->1	
pa.Re	g->1	
pa.Tr	o->1	
pa.Ty	 ->1	
pa.Un	d->1	
pa.Va	d->1	
pa.Vi	 ->8	d->1	
pa.Äv	e->1	
pa; e	n->1	
pa?He	r->1	
pa?Va	d->1	
pa?Vi	 ->1	
paNäs	t->1	
pacit	e->5	
packn	i->5	
pad a	n->1	
pad b	i->1	
pad k	o->1	
pade 	d->1	e->1	g->2	k->1	m->2	o->2	s->2	t->2	
padem	o->2	
pades	 ->9	
pagan	d->3	
pager	a->1	
pagne	-->1	
pagru	p->1	
paket	 ->3	.->1	e->3	
pakon	v->1	
pakt 	s->1	
pakte	n->4	
pales	t->12	
pamin	i->1	
pan e	l->1	
pan o	c->1	
pan, 	K->1	
pande	 ->36	r->5	t->23	
panel	e->1	
panie	n->7	
paniv	å->1	
panj 	f->2	m->1	
panj.	D->1	
panje	n->1	r->1	
panjo	r->1	
pansi	o->1	
pansk	 ->2	a->6	t->3	
pante	n->1	
papar	l->166	
pappe	r->5	
par -	 ->1	
par a	l->1	n->1	r->1	t->1	v->2	
par b	e->1	ä->1	
par d	e->8	i->1	ä->1	
par e	f->1	n->5	t->2	
par f	a->1	ö->3	
par g	å->1	
par h	ä->1	
par i	 ->1	d->1	n->1	
par j	a->1	
par k	o->1	
par m	a->1	e->1	i->5	ö->1	
par n	å->1	
par o	c->3	r->1	s->1	
par p	e->1	u->3	å->1	
par r	å->1	
par s	i->1	n->1	v->2	y->1	å->1	
par u	r->1	
par v	i->3	ä->1	å->1	
par å	r->2	
par ö	s->1	v->1	
par.A	t->1	
par.D	e->1	
par.I	n->1	
para 	d->1	e->1	i->1	o->1	
parab	l->1	
parad	o->6	
parag	r->2	
paral	l->5	
param	e->2	
parar	 ->3	
parat	 ->1	e->1	i->1	
parco	u->1	
pare 	E->1	a->2	f->1	o->1	
pare,	 ->1	
pare.	E->1	
parer	a->4	
paric	i->1	
parin	g->3	
park 	i->1	o->1	t->1	v->1	
parka	r->1	s->2	
parke	n->4	r->3	
parla	m->558	
parna	.->1	
parsa	m->1	
part 	t->1	
part.	Ä->1	
parte	m->9	n->1	r->21	
parti	 ->23	,->7	.->4	e->42	i->1	k->1	l->1	p->2	s->5	
partn	e->28	
parts	m->1	
paråd	e->1	
pas -	 ->2	
pas a	t->51	v->9	
pas b	e->2	i->1	l->1	
pas c	e->1	
pas d	e->3	j->1	
pas e	f->1	k->1	n->3	
pas f	i->1	o->2	r->2	u->1	å->2	ö->10	
pas g	a->1	e->2	
pas h	i->1	j->1	
pas i	 ->8	g->1	n->3	
pas j	a->10	
pas k	o->6	u->2	
pas l	e->1	i->2	
pas m	e->9	
pas n	a->3	i->1	o->1	ä->1	
pas o	c->8	l->1	
pas p	o->1	å->9	
pas r	u->1	ä->1	
pas s	a->2	j->1	k->6	l->1	o->1	t->1	v->1	y->1	å->1	
pas t	r->1	u->1	
pas u	n->1	
pas v	a->2	e->7	i->2	ä->2	
pas å	t->1	
pas, 	a->1	m->1	s->3	
pas.-	 ->1	
pas.D	e->3	ä->1	
pas.J	a->1	
pas.K	o->1	
pas.P	a->1	
pas.V	a->1	i->1	
pas: 	a->1	
pas?S	k->1	
pass 	f->1	o->1	t->1	v->1	
passa	 ->6	d->3	g->1	n->2	r->1	s->5	
passe	r->3	
passi	o->2	v->1	
passn	i->4	
passu	s->1	
past 	e->2	h->1	k->1	n->1	o->1	r->1	ä->2	
paste	 ->2	
pat -	 ->1	
pat d	e->1	
pat e	n->2	t->1	
pat f	ö->1	
pat m	o->1	
pat n	å->2	
pat s	t->1	ä->2	å->1	
pat t	i->1	
pat.F	P->1	
pat: 	"->1	
patet	i->1	
pati 	f->3	m->1	
patie	n->4	r->1	
patio	n->1	
patis	e->2	k->1	
patjä	n->1	
patri	o->1	
pats 	a->2	g->1	i->2	o->1	p->1	v->1	
pats.	D->1	
paval	e->3	
payan	n->2	
pback	n->1	
pbrin	g->3	
pbygg	a->6	d->1	n->12	t->1	
pbära	 ->1	
pbåda	 ->1	
pdate	r->3	
pdeln	i->3	
pdrag	 ->17	.->1	e->4	
pe i 	h->1	
pe på	 ->1	
peanu	t->1	
peau"	,->1	
pecia	l->14	
pecie	l->42	
pecif	i->29	
pedag	o->1	
pedit	i->1	
pedof	i->1	
pegla	 ->2	r->7	s->2	
pegli	n->1	
pegna	 ->1	
pehål	l->13	
peise	r->2	
peisk	 ->102	.->1	a->585	e->2	t->20	
peka 	B->1	a->7	d->2	f->3	p->6	v->1	
peka,	 ->1	
pekad	e->10	
pekan	d->9	
pekar	 ->11	,->1	
pekas	 ->3	,->1	
pekat	 ->9	,->4	.->1	
pekt 	a->3	f->18	h->1	m->1	s->3	v->1	
pekt:	 ->1	
pekta	b->3	k->3	
pekte	n->17	r->51	
pekti	o->6	v->32	
pektr	u->2	
pektö	r->6	
pekul	a->4	
pel -	 ->2	
pel B	a->1	
pel N	y->1	
pel R	i->1	
pel a	t->1	v->1	
pel b	e->1	l->1	
pel d	e->1	
pel e	t->1	
pel f	a->1	r->1	ö->9	
pel g	e->2	
pel h	a->3	j->1	ä->2	
pel i	 ->4	n->2	
pel m	e->1	
pel n	i->1	ä->1	
pel o	c->2	m->2	
pel p	å->20	
pel r	i->1	
pel s	e->1	k->3	o->1	ä->2	
pel t	i->1	r->1	
pel u	n->1	
pel v	i->1	
pel ä	n->1	r->1	
pel, 	a->1	e->2	l->1	m->2	v->1	
pel.D	e->1	
pel.I	 ->1	
pel.J	a->1	
pel.M	e->1	
pel.V	i->1	
pel: 	E->1	F->1	d->1	
pel; 	i->1	
pela 	d->1	e->8	i->3	o->1	v->1	
pela?	A->1	
pelad	e->1	
pelar	 ->12	e->9	n->3	
pelas	 ->1	
pelat	 ->5	
pelen	.->1	
pelet	 ->1	
pell 	g->1	
pelni	n->1	
pelpl	a->1	
pelre	g->4	
pelru	m->1	
pelvi	s->28	
pen "	T->2	d->1	
pen (	1->1	K->1	
pen -	 ->1	
pen D	e->4	
pen E	u->2	
pen N	a->2	
pen T	o->1	
pen U	n->2	
pen a	l->1	n->1	t->6	v->16	
pen b	a->1	e->3	ö->2	
pen d	ä->1	
pen e	g->1	l->1	r->1	t->1	
pen f	i->1	r->1	ä->1	ö->7	
pen g	a->1	o->2	ä->2	
pen h	a->11	o->1	
pen i	 ->8	n->6	
pen k	a->3	o->3	r->2	
pen m	a->2	e->4	o->12	å->1	
pen n	ä->5	å->1	
pen o	c->12	m->25	n->1	
pen p	å->4	
pen s	k->6	o->8	t->1	y->1	
pen t	i->4	
pen u	n->1	t->3	
pen v	a->2	e->1	i->3	o->1	
pen ä	n->2	r->14	
pen å	 ->2	t->1	
pen, 	b->2	d->1	e->3	f->1	k->2	m->3	o->5	p->1	s->3	u->1	v->2	ä->2	
pen. 	F->1	
pen..	 ->1	
pen.D	e->6	
pen.E	n->1	
pen.H	e->3	
pen.J	a->7	
pen.K	o->1	
pen.M	a->1	o->1	
pen.N	i->1	u->1	ä->1	
pen.P	r->1	
pen.S	a->1	o->2	
pen.T	a->1	i->1	
pen.V	i->1	
pen.Ä	n->1	
pen: 	J->1	m->1	
pen?.	 ->1	
penNä	s->1	
penba	r->36	
pence	r->1	
pende	r->5	
pendi	e->1	
penga	r->55	
penha	m->1	n->1	
penhe	t->60	
penin	d->1	
pennd	r->1	
penni	n->10	
pens 	B->2	b->6	d->3	e->4	f->7	g->2	h->1	i->4	j->1	k->6	l->4	m->5	n->1	r->19	s->6	t->1	v->6	y->3	ä->1	å->2	
pensa	t->3	
pense	r->8	
pensi	o->13	v->1	
pensp	r->1	
pente	k->1	
penut	v->1	
per E	U->1	
per a	n->1	v->5	
per b	i->2	l->1	
per c	a->10	
per d	e->5	o->1	
per e	l->3	n->3	
per f	r->4	å->1	ö->3	
per h	a->4	
per i	 ->4	n->6	
per j	ä->1	
per k	a->1	o->1	u->1	
per l	a->1	ö->1	
per m	a->1	e->2	o->1	ö->1	
per n	i->1	
per o	c->8	m->4	s->1	
per p	r->2	
per r	i->3	
per s	e->1	k->1	o->13	å->1	
per t	i->3	
per u	p->1	t->5	
per v	i->2	
per ä	n->1	r->4	
per å	r->3	
per, 	a->1	f->1	i->1	n->1	o->2	s->1	u->1	v->1	
per.A	l->1	
per.E	n->2	
per.F	ö->3	
per.G	e->1	
per.I	 ->1	
per.N	ä->1	
per.O	m->1	
per.V	i->2	
per: 	d->1	v->1	
pera 	o->1	
perad	e->2	
perah	u->1	
peras	 ->1	
perat	 ->2	i->9	u->4	ö->2	
perer	a->1	
peret	 ->1	
perfe	k->7	
perif	e->6	
perin	g->2	
perio	d->86	
perli	g->1	
perma	n->8	
pern 	h->1	
perna	 ->30	,->7	.->6	s->6	
peron	i->1	
perro	n->1	
pers 	s->1	
persl	u->1	
perso	n->104	
persp	e->17	
perte	r->20	
pertg	r->3	
perti	s->3	
pertk	o->17	
pertr	a->1	e->1	
pertu	t->1	
pes e	l->1	
pes r	e->1	
peskå	l->1	
pessi	m->2	
pest 	o->1	
peste	n->4	
pet "	e->2	k->1	
pet (	t->1	
pet -	 ->2	
pet a	t->1	v->2	
pet b	e->2	
pet d	e->3	
pet e	l->1	x->1	
pet f	r->2	ö->7	
pet g	j->1	
pet h	a->3	
pet i	 ->3	n->2	
pet j	u->1	
pet k	a->4	o->8	v->1	
pet l	i->1	y->1	
pet m	e->1	o->1	å->5	
pet n	o->1	ä->1	
pet o	c->16	
pet p	l->1	o->1	r->1	å->3	
pet r	e->1	
pet s	a->1	e->2	k->1	o->3	y->1	ä->2	
pet t	a->1	i->2	r->1	
pet v	a->1	i->2	ä->1	
pet ä	v->1	
pet ö	p->1	
pet) 	h->1	
pet, 	a->1	b->1	d->2	f->4	k->1	n->1	o->3	s->2	v->1	ä->2	
pet.H	e->1	
pet.J	a->1	
pet.M	a->1	i->1	
pet.N	u->1	
pet.O	c->1	
pet.P	a->1	
pet?R	I->1	
peten	s->7	t->4	
petit	i->1	
pets 	"->1	a->1	f->2	i->2	l->1	m->1	n->1	p->2	s->1	u->1	v->1	å->1	
pets.	E->1	
petsf	ö->1	
pfall	 ->1	
pfann	s->1	
pfatt	a->13	n->38	
pfyll	a->31	d->1	e->19	s->2	t->1	
pfödn	i->1	
pfölj	n->10	
pföra	 ->1	n->11	
pförs	 ->1	
pgick	 ->3	
pgift	 ->21	!->1	,->2	.->6	:->1	e->43	s->3	
pgodk	ä->1	
pgrad	e->1	
pgå t	i->1	
pgåen	d->7	
pgång	.->2	
pgår 	i->1	t->4	
pgöre	l->2	
pharm	a->1	
pherd	s->3	
phet 	a->1	f->1	
phet,	 ->1	
phets	a->1	
phov 	t->8	
phovs	m->5	
phtal	a->1	
phänt	a->1	
phäva	s->3	
phävs	.->2	
phål 	i->1	
phål:	 ->1	
phåle	n->1	
phöjs	 ->1	
phör 	a->2	e->1	
phöra	 ->3	.->2	
phört	.->1	
pia t	i->1	
pic B	r->1	
pice 	f->1	
piell	a->3	t->5	
pien 	o->1	
pien,	 ->2	
piera	 ->1	
pillo	l->1	
pilot	 ->1	e->1	p->2	
pin h	a->1	
pinio	n->4	
pionj	ä->1	
pirat	e->1	
pirer	a->3	
piska	 ->2	
pit o	m->1	
pit s	i->1	
pita 	h->1	i->2	o->1	v->1	ä->1	
pita,	 ->1	
pita.	D->1	M->1	S->1	
pital	 ->5	,->1	.->1	e->5	i->2	s->3	
pitel	 ->6	
pitul	e->2	
pjakt	 ->1	
pkay 	f->2	h->1	
pkay,	 ->3	
pkay.	V->1	
pkayD	e->1	
pkayb	e->1	
pkays	 ->2	
pkoll	e->1	
pkomm	e->6	
pkraf	t->1	
pla s	a->1	
place	r->17	
plade	 ->1	
plan 	e->1	f->7	k->1	m->2	o->2	r->1	s->3	u->2	
plan,	 ->2	
plan.	D->2	I->1	V->1	
plan:	 ->1	
planN	ä->1	
pland	 ->2	
plane	n->13	r->84	t->3	
plant	e->2	o->1	
plari	s->2	
plas 	b->1	t->1	
plast	 ->3	!->1	,->2	
plats	 ->17	,->7	.->1	e->19	
platt	a->1	
pleme	n->11	
plen 	m->2	v->1	
plena	r->4	
plenu	m->5	
plet 	V->1	f->1	k->1	
plett	 ->1	e->13	
pleva	 ->7	
plevd	e->1	
pleve	l->1	r->3	
plevs	 ->2	
plevt	 ->3	
plex 	f->1	
plex.	J->1	
plexa	,->1	
plext	 ->1	
plice	r->12	
plici	t->1	
plig 	e->1	h->1	i->5	k->1	n->2	o->1	p->1	r->2	s->1	u->1	y->1	å->1	
plig,	 ->2	
plig.	J->1	
pliga	 ->42	r->1	s->1	
pligh	e->4	
pligt	 ->32	,->1	.->2	
plikt	 ->5	.->2	a->4	e->17	i->5	
plima	n->3	
plime	n->1	
plims	o->1	
plin 	f->1	i->1	n->1	o->1	
plin,	 ->1	
pline	r->3	
plinf	r->1	
pling	 ->1	.->2	
plinr	å->1	
plinä	r->4	
plitt	r->4	
pliva	 ->1	
ploma	t->11	
plosi	o->1	v->1	
plund	r->1	
plura	l->1	
plus 	a->1	t->1	
plysa	 ->2	
plysn	i->2	
pläde	r->2	
plåde	r->11	
plåge	r->1	
plåna	n->1	
plånb	o->1	
plåni	n->1	
plösa	 ->1	
plöse	s->1	
plösn	i->1	
plöst	 ->1	
plöts	l->4	
pmana	 ->12	d->2	r->31	s->4	t->2	
pmani	n->7	
pmjuk	n->2	
pmunt	r->21	
pmärk	s->53	
pmätt	a->1	e->1	
pmöte	n->1	t->11	
pna d	e->1	
pna f	ö->2	
pna g	r->1	
pna m	a->1	
pna o	c->1	
pna p	a->1	r->1	
pna r	e->1	
pna, 	d->1	o->1	
pnade	 ->3	
pnar 	d->1	f->1	
pnare	 ->1	
pnas 	d->1	f->1	
pnen 	m->1	p->1	
pning	 ->47	,->4	.->12	a->8	e->33	s->15	
pnå d	a->1	e->10	
pnå e	k->2	n->14	t->5	
pnå f	a->1	r->1	
pnå g	e->1	
pnå m	e->2	å->1	
pnå n	å->1	
pnå p	å->2	
pnå r	e->1	
pnå s	i->1	
pnå v	å->4	
pnå y	t->1	
pnå ö	n->1	
pnå, 	n->1	
pnå. 	D->1	
pnå.F	r->1	
pnå.J	a->1	
pnå.S	l->1	
pnådd	a->3	e->3	
pnår 	d->4	e->4	m->3	s->1	v->1	
pnås 	b->1	e->1	g->1	i->2	
pnås.	F->1	L->1	
pnått	 ->6	,->1	.->1	s->5	
po, s	o->1	
poet 	a->1	
pok i	 ->1	
pok, 	m->1	
poken	 ->2	
pol a	t->1	v->1	
pol i	 ->1	n->1	
pol m	e->1	å->1	
pol o	c->6	
pol s	o->2	
pol t	i->1	
pol, 	i->1	o->1	p->1	
pol-f	ö->1	
pol.E	u->1	
pol.H	e->1	
pol; 	f->1	
polav	t->1	
pole 	p->1	
polem	i->1	
polfr	å->1	
polfö	r->2	
polic	y->4	
polin	t->1	
polis	,->1	.->1	;->1	a->1	e->8	i->1	m->2	s->2	v->1	
polit	a->1	i->533	
polko	n->1	
pols 	a->1	m->1	u->1	
polsi	t->1	
ponde	n->1	
ponen	t->5	
poner	a->7	
pons 	f->1	
ponsr	a->1	
ponta	n->4	
pool,	 ->1	
popul	a->1	i->4	ä->2	
por, 	s->1	
pordf	ö->1	
porno	g->2	
porsl	i->1	
port 	a->23	b->3	d->1	f->5	h->3	i->3	l->1	m->1	o->26	p->2	r->1	s->6	t->1	v->3	ä->2	ö->2	
port)	 ->1	
port,	 ->9	
port-	 ->1	s->2	
port.	N->1	U->1	V->1	
portN	ä->1	
porta	b->1	
portb	e->2	
portd	i->1	
porte	n->46	r->63	
portf	e->1	r->1	ö->1	
portg	r->1	
porti	o->9	
portk	o->2	
portm	a->1	o->1	
portn	ä->1	
porto	m->3	
portp	r->1	
ports	i->1	ä->7	
portu	g->70	n->2	t->1	
portv	i->1	
porär	 ->1	t->1	
pos b	e->1	
posit	i->87	
post 	a->1	f->2	o->1	t->1	u->1	v->1	
post.	N->1	
poste	n->1	r->5	
postv	e->1	
poten	t->6	
potes	e->1	
potet	i->1	
potis	m->5	
pots 	s->1	
poulo	s->5	
poäng	 ->1	.->1	s->2	t->8	
pp (k	r->2	
pp - 	o->1	s->1	
pp Eu	r->1	
pp Ti	b->1	
pp al	l->5	
pp an	s->3	t->1	v->1	
pp at	t->3	
pp av	 ->10	s->1	
pp be	g->1	t->1	
pp bi	d->1	
pp bå	d->1	
pp de	 ->9	b->2	m->2	n->13	s->3	t->11	
pp do	m->1	
pp dä	r->1	
pp ef	t->3	
pp el	l->1	
pp en	 ->10	
pp et	t->6	
pp ex	p->1	
pp fo	r->1	
pp fr	a->2	å->9	
pp fu	l->1	
pp fö	r->12	
pp ge	n->2	
pp gr	ä->1	
pp ha	d->1	r->5	
pp he	l->1	
pp hu	v->1	
pp hä	n->2	r->1	
pp hö	g->1	
pp i 	E->1	b->1	d->6	e->2	m->3	p->2	r->1	s->2	t->2	v->1	ä->1	
pp id	é->1	
pp ig	e->4	
pp in	l->1	o->1	t->1	
pp ka	n->1	
pp ko	m->5	n->1	
pp la	g->1	
pp li	v->1	
pp lä	g->1	m->1	n->1	
pp me	d->8	
pp må	s->1	
pp na	t->1	
pp ny	a->1	
pp nå	g->3	
pp oc	h->6	
pp ol	j->1	
pp om	 ->2	
pp or	d->2	
pp po	s->1	
pp pr	i->1	o->2	
pp på	 ->10	.->2	
pp re	f->1	g->1	
pp rä	c->1	t->2	
pp rö	s->1	
pp sa	d->1	
pp si	g->1	t->1	
pp sk	a->2	y->1	
pp so	m->7	
pp st	ä->2	
pp sä	r->1	t->1	
pp så	v->1	
pp ti	l->11	
pp to	g->1	
pp tr	e->1	
pp tv	å->1	
pp ty	d->1	v->1	
pp un	d->2	
pp ut	a->1	g->1	t->3	v->2	
pp va	d->3	
pp vi	l->2	
pp vä	l->2	
pp än	 ->1	d->1	
pp är	 ->4	,->1	e->2	
pp, E	D->1	
pp, a	n->1	v->1	
pp, b	l->1	
pp, d	e->1	
pp, e	f->3	n->1	
pp, f	å->1	
pp, h	e->2	
pp, i	 ->1	
pp, j	u->1	
pp, m	e->1	i->1	
pp, n	u->1	
pp, o	c->2	
pp, r	i->1	
pp, s	o->2	ä->1	
pp, v	i->1	
pp..(	F->1	
pp.Ah	e->1	
pp.De	n->2	t->3	
pp.Fa	k->1	
pp.Ja	g->7	
pp.Me	n->1	
pp.På	 ->1	
pp.Vi	 ->2	l->1	
pp.Än	d->1	
pp.Äv	e->1	
pp?Hu	r->1	
ppa a	n->1	
ppa e	n->1	u->1	
ppa i	 ->1	h->1	n->4	
ppa m	a->1	
ppa r	e->1	
ppa s	i->1	
ppa t	i->4	
ppa ö	v->1	
ppade	 ->3	s->5	
ppand	e->2	
ppar 	d->1	m->1	u->1	
ppara	t->1	
ppas 	-->2	a->51	f->3	i->2	j->10	k->3	n->3	o->4	p->4	s->3	v->10	å->1	
ppas,	 ->4	
ppast	 ->9	
ppbac	k->1	
ppbri	n->3	
ppbyg	g->20	
ppbär	a->1	
ppbåd	a->1	
ppdat	e->3	
ppdel	n->3	
ppdra	g->22	
ppe i	 ->1	
ppehå	l->13	
ppell	 ->1	
ppen 	"->2	D->4	E->2	N->2	T->1	U->2	a->7	b->1	d->1	f->4	g->2	h->3	i->3	k->5	m->2	n->2	o->3	p->1	s->5	t->2	u->1	v->4	ä->2	
ppen,	 ->4	
ppen.	H->1	J->2	N->1	
ppenb	a->36	
ppenh	e->60	
ppens	 ->13	
pper 	a->2	b->1	e->1	f->3	h->3	i->6	k->1	m->1	n->1	o->3	s->4	t->2	u->1	v->1	ä->2	
pper,	 ->4	
pper.	A->1	E->1	G->1	I->1	N->1	
pper:	 ->1	
ppera	s->1	
ppere	t->1	
pperi	n->2	
pperl	i->1	
ppern	a->21	
ppers	 ->1	l->1	
ppet 	"->3	a->2	e->1	f->3	i->1	j->1	k->2	l->1	m->2	o->8	p->1	s->4	t->1	v->1	ö->1	
ppet,	 ->2	
ppet.	O->1	
ppfan	n->1	
ppfat	t->51	
ppfyl	l->54	
ppföd	n->1	
ppföl	j->10	
ppför	a->12	s->1	
ppgic	k->3	
ppgif	t->77	
ppgra	d->1	
ppgå 	t->1	
ppgån	g->2	
ppgår	 ->5	
ppgör	e->2	
pphet	 ->2	,->1	s->1	
pphov	 ->8	s->5	
pphän	t->1	
pphäv	a->3	s->2	
pphöj	s->1	
pphör	 ->3	a->5	t->1	
ppjak	t->1	
ppkol	l->1	
ppkom	m->6	
ppla 	s->1	
pplad	e->1	
pplan	d->2	
pplas	 ->2	
pplev	a->7	d->1	e->4	s->2	t->3	
pplin	g->2	
ppliv	a->1	
pplys	a->2	n->2	
pplåd	e->11	
pplös	a->1	e->1	n->1	t->1	
ppman	a->51	i->7	
ppmju	k->2	
ppmun	t->21	
ppmär	k->53	
ppmät	t->2	
ppmöt	e->12	
ppna 	d->1	f->2	g->1	m->1	o->1	p->1	r->1	
ppna,	 ->2	
ppnad	e->1	
ppnar	 ->2	e->1	
ppnas	 ->2	
ppnin	g->17	
ppnå 	d->11	e->21	f->2	g->1	m->3	n->1	p->2	r->1	s->1	v->4	y->1	ö->1	
ppnå,	 ->1	
ppnå.	 ->1	F->1	J->1	S->1	
ppnåd	d->6	
ppnår	 ->13	
ppnås	 ->5	.->2	
ppnåt	t->13	
ppone	r->3	
ppord	f->1	
pport	 ->40	)->1	,->7	.->1	N->1	e->61	s->1	u->2	
pposi	t->2	
ppren	s->2	
pprep	a->51	n->1	
pprik	t->6	
pprop	 ->3	,->1	.->1	
pprus	t->1	
ppryc	k->1	
ppräc	k->2	
ppräk	n->1	
pprät	t->36	
pprör	a->3	d->2	
pps u	t->1	
pps v	ä->3	
ppsam	l->4	
ppsat	t->3	
ppsbr	o->1	
ppsby	g->1	
ppska	t->23	
ppskj	u->4	
ppsko	v->2	
ppspå	r->2	
ppsre	d->2	
ppsrä	t->1	
ppsst	ä->1	
ppssä	t->2	
ppsto	d->4	
ppstä	l->3	
ppstå	 ->3	:->1	n->1	r->16	t->11	
ppsva	r->2	
ppsäg	n->1	
ppsät	t->2	
ppt e	n->1	t->1	
ppt i	n->1	
ppt s	e->1	
ppt t	r->1	
pptag	a->3	e->2	n->2	
pptar	 ->1	
pptas	 ->1	.->1	
ppte 	l->1	
pptes	 ->2	
pptil	l->1	
pptog	s->2	
ppträ	d->9	t->1	
pptäc	k->11	
ppund	a->1	
ppver	k->2	
ppvig	l->1	
ppvis	.->1	a->4	
ppväg	a->1	
ppvär	d->1	
ppy e	n->1	
prack	a->1	
pragm	a->1	
prakt	i->33	
prana	t->1	
prat.	B->1	
prata	 ->3	r->1	
praxi	s->8	
preci	s->43	
prefe	r->3	
preju	d->4	
preli	m->3	
premi	ä->10	
prens	n->2	
prenö	r->3	
prepa	 ->15	,->1	d->8	r->15	s->7	t->5	
prepn	i->1	
prero	g->1	
prese	n->47	
presi	d->9	
press	 ->3	a->3	e->9	i->2	k->2	m->1	n->1	
prest	a->4	
prick	a->1	f->1	n->1	
prida	 ->2	n->1	s->1	
pride	r->5	
pridi	t->1	
pridn	i->8	
prids	 ->2	
prikt	i->6	
pril 	1->1	f->1	
pril.	J->1	
primi	t->1	
princ	i->194	
prini	p->1	
prior	i->38	
pris 	f->3	å->1	
pris.	S->1	
prisa	 ->1	
prise	r->10	s->2	t->7	
prisn	i->1	
priss	ä->1	
prisu	t->1	
priva	t->21	
privi	l->7	
probl	e->174	
proce	d->1	n->93	s->107	
produ	c->27	k->49	
profe	s->7	
profi	l->3	
progr	a->237	e->1	
proje	k->62	
prokl	a->1	
promi	s->22	
prona	z->1	
prop 	o->2	s->1	
prop,	 ->1	
prop.	S->1	
propa	g->4	
propo	r->9	
propå	 ->1	
prost	i->1	
prote	k->4	s->9	
proto	k->24	
prov 	p->9	
provi	n->3	s->2	
provk	a->1	
provs	k->2	t->1	
prung	 ->2	.->2	e->2	l->12	s->1	
prust	a->1	
pryck	n->1	
präck	n->2	
prägl	a->5	
präkn	i->1	
pränt	a->1	
prätt	a->27	h->9	
pråk 	f->1	p->3	t->1	
pråk.	 ->1	
pråka	 ->1	r->8	
pråke	t->3	
pråkl	i->3	
pråko	m->2	
pråkt	a->1	
prång	,->2	
pröra	 ->1	n->1	s->1	
prörd	a->1	h->1	
pröva	 ->4	r->1	s->4	
prövn	i->5	
prövo	å->1	
ps av	 ->1	
ps fa	k->1	
ps ut	t->1	
ps vä	g->3	
ps- o	c->1	
ps.Ju	s->1	
ps.Me	n->1	
psaml	i->4	
psatt	a->3	
psavt	a->2	
psbef	o->1	
psbeg	r->1	
psbes	l->1	t->1	
psbro	t->1	
psbyg	g->1	
psdir	e->1	
psfrå	g->1	
psini	t->7	
psinn	i->1	
psins	a->1	t->5	
psint	r->1	
psis 	n->1	
pskat	t->23	
pskhe	t->1	
pskju	t->4	
pskon	c->1	s->1	t->1	
pskov	 ->1	e->1	
pskäl	 ->1	.->1	
pslag	 ->2	n->1	s->2	
psmas	k->2	
psmed	b->1	
psmän	 ->10	n->6	
psmål	 ->1	
psniv	å->11	
pson 	h->1	
psorg	a->1	
pspel	a->2	
pspol	i->2	
pspro	d->1	g->2	
pspår	a->1	n->1	
psram	e->1	
psred	a->2	
psreg	i->1	l->8	
psrät	t->9	
psstr	a->1	
psstä	m->1	
psstö	d->2	
pssys	t->1	
pssät	t->2	
pstod	 ->4	
pstäl	l->3	
pstå 	f->1	n->1	o->1	
pstå:	 ->1	
pstån	d->1	
pstår	 ->13	,->1	.->2	
pståt	t->11	
psvar	v->2	
psyko	l->1	
psägn	i->1	
psätt	n->2	
psåtg	ä->2	
pt be	k->1	s->1	
pt de	n->1	
pt di	s->1	
pt en	s->1	
pt et	t->1	
pt fo	r->1	
pt i 	F->1	t->1	
pt in	l->1	
pt ko	m->1	
pt or	o->1	
pt se	x->1	
pt sk	a->1	
pt ti	l->1	
pt tr	e->1	
pt ut	,->2	.->3	
pt va	t->1	
pt öv	e->1	
pt.De	n->1	
pt.Ha	n->1	
pta k	r->1	
pta v	i->1	
pta.D	e->1	
ptabe	l->27	
ptabl	a->10	
ptaga	n->3	
ptage	n->2	
ptagn	a->2	
ptans	 ->3	,->2	e->2	
ptar 	a->1	
ptas 	s->1	
ptas.	V->1	
pte d	e->1	
pte f	r->1	
pte l	ö->1	
pte t	i->1	
pte u	t->2	
ptemb	e->15	
pten 	o->2	p->1	
pten,	 ->1	
ptera	 ->16	,->1	.->7	d->3	n->2	r->5	s->8	t->3	
ptes 	i->1	t->1	
ptet 	b->1	f->2	
ptike	r->3	
ptill	h->1	
ptima	l->3	
ptimi	s->4	
ption	 ->2	.->1	e->7	s->4	
ptisk	 ->2	,->1	a->1	t->1	
ptoga	m->2	
ptogs	 ->2	
ptom 	o->1	
pträd	a->5	e->4	
pträt	t->1	
ptäck	a->3	e->2	s->2	t->4	
publi	c->6	k->20	
pular	i->1	
pulis	m->1	t->3	
puls 	f->1	t->1	
pulse	r->4	
pulär	a->1	t->1	
pumpa	s->2	
pund 	e->1	f->1	
pund.	D->1	
punda	n->1	
punkt	 ->131	,->14	.->19	:->2	?->1	e->173	s->2	
purit	a->1	
pus j	u->5	
pverk	 ->1	,->1	
pvigl	a->1	
pvill	i->1	
pvis.	Ä->1	
pvisa	 ->1	r->1	s->1	t->1	
pväga	 ->1	
pvärd	e->1	
py en	d->1	
pyram	i->1	
pyrig	h->1	
pänna	 ->1	n->3	
pänni	n->7	
pärr 	n->1	
pärra	r->2	
på - 	a->1	m->1	o->2	s->1	
på 10	 ->1	
på 13	 ->2	
på 14	0->1	
på 20	 ->1	0->2	
på 22	,->1	
på 33	 ->1	
på 34	 ->1	
på 37	 ->1	
på 40	 ->1	
på 5 	m->1	
på 50	 ->1	-->1	
på 7,	2->1	
på 75	 ->1	
på 80	 ->2	
på 86	 ->1	
på 90	 ->1	
på 95	 ->1	
på Al	l->2	
på At	l->1	
på BS	E->1	
på Ba	l->5	
på Be	l->1	
på CE	N->1	
på CS	U->1	
på EG	-->3	
på EU	-->2	:->2	
på Er	i->1	
på Eu	r->10	
på Fö	r->1	
på Ge	n->1	
på Go	l->1	
på Ho	l->1	
på IS	P->1	
på In	t->6	
på Ir	l->1	
på Is	r->1	
på Ma	l->1	
på Ol	i->1	
på Pa	p->1	
på Ri	c->2	
på Ro	i->1	
på Ty	s->1	
på Vä	s->2	
på ac	c->1	
på ak	t->1	
på al	b->1	l->28	
på an	d->11	g->1	n->1	s->3	
på ar	b->6	g->1	t->4	
på as	y->1	
på at	t->145	
på av	f->1	
på ba	l->1	r->1	s->2	
på be	f->1	h->4	k->1	t->2	
på bi	l->5	
på bl	y->1	
på bo	r->2	s->1	
på br	e->3	i->1	o->3	
på bä	s->8	t->1	
på bå	d->3	
på ce	n->1	
på ci	v->1	
på cr	i->1	
på da	g->7	n->1	
på de	 ->48	b->2	f->1	l->1	m->7	n->95	r->3	s->9	t->126	
på di	r->2	
på dj	u->7	
på du	b->3	m->1	
på dy	l->1	
på ef	f->1	t->1	
på eg	e->3	
på ek	o->2	
på el	e->1	
på em	b->1	
på en	 ->51	d->1	g->1	h->1	s->1	
på er	 ->3	,->1	t->1	
på et	t->142	
på eu	r->12	
på ex	a->1	
på fa	m->1	r->2	
på fe	l->1	m->2	n->1	
på fi	s->2	
på fl	e->2	y->1	
på fr	a->3	e->1	i->1	å->7	
på fy	r->2	
på fä	l->5	r->1	
på fö	l->3	r->59	t->2	
på ga	t->1	
på ge	m->13	n->2	o->1	
på gl	o->1	
på go	d->1	t->1	
på gr	u->78	ä->1	
på gä	l->1	
på gå	n->4	r->1	
på gö	r->1	
på ha	t->1	v->4	
på he	m->1	
på hj	ä->1	
på hu	r->14	
på hä	n->1	
på hö	g->1	
på i 	d->1	f->3	
på ic	k->1	
på il	l->1	
på in	f->2	i->1	l->1	n->2	r->1	s->3	t->8	v->1	
på it	a->1	
på ja	k->1	
på jo	r->1	
på ju	s->2	
på jä	r->3	
på ka	m->2	n->1	t->2	
på kl	a->1	i->1	
på kn	u->1	
på ko	l->4	m->10	n->17	r->6	
på kr	a->1	
på ku	n->1	
på kv	a->1	
på kä	r->1	
på kö	r->1	
på la	g->2	n->10	
på li	k->1	s->2	
på lo	b->1	k->2	
på lä	m->3	n->3	
på lå	g->2	n->7	
på lö	r->1	
på ma	r->12	
på me	d->14	l->2	n->1	r->2	
på mi	g->2	l->10	n->15	t->1	
på mo	d->2	n->1	t->3	
på my	c->2	
på mä	n->1	
på må	l->1	n->4	
på mö	j->4	
på na	t->4	
på ne	d->1	
på no	r->3	t->1	
på ny	 ->2	a->3	t->21	
på nä	r->3	s->4	t->1	
på nå	g->21	
på ob	e->2	
på oc	h->3	k->1	
på ol	i->2	j->2	
på om	 ->4	k->1	r->14	
på on	s->2	
på or	d->2	
på os	s->5	
på pa	r->1	
på pe	n->1	r->2	
på pl	a->9	
på po	l->1	
på pr	i->5	o->4	
på ra	s->1	t->1	
på re	f->2	g->13	k->1	s->10	
på ri	k->1	s->1	
på ry	g->1	
på rä	d->1	t->10	
på rå	d->7	
på sa	k->1	m->21	
på se	d->1	k->3	m->1	n->5	r->1	
på si	f->1	g->7	k->7	n->10	s->1	t->5	
på sj	ä->1	
på sk	a->3	i->1	o->1	u->1	
på sl	u->1	
på sm	å->1	
på sn	a->1	
på so	c->1	
på sp	e->9	å->1	
på st	a->7	o->2	r->1	u->1	ö->2	
på su	b->2	
på sv	a->1	
på sy	d->1	s->3	
på sä	k->2	t->3	
på så	 ->14	d->2	
på ta	l->6	n->1	
på te	k->1	m->1	r->1	x->1	
på ti	d->5	l->5	
på tj	ä->1	
på to	p->1	r->9	
på tr	a->3	e->4	ö->3	
på tv	ä->1	å->6	
på tä	n->1	
på un	d->3	i->5	
på up	p->3	
på ut	f->1	s->1	v->3	
på va	d->9	l->2	r->4	t->1	
på ve	d->4	r->1	t->3	
på vi	d->1	l->13	s->2	
på vä	g->29	r->3	s->2	
på vå	r->16	
på yt	t->1	
på zi	g->1	
på Ös	t->2	
på än	d->4	n->2	
på är	 ->3	
på åh	ö->1	
på år	 ->1	
på åt	a->1	e->1	g->3	
på ök	a->1	
på ön	 ->1	
på öp	p->5	
på öv	e->1	
på, e	l->1	t->1	
på, f	ö->1	
på, h	u->1	
på, l	ö->1	
på, m	e->3	
på, n	ä->1	
på, o	c->4	m->1	
på, v	i->1	
på, ä	r->1	
på.Be	t->1	
på.De	t->3	
på.Do	c->1	
på.En	 ->1	
på.Eu	r->1	
på.Ja	g->3	
på.No	r->1	
på.Or	d->1	
på.Un	i->1	
på.Vi	 ->1	
på.Är	 ->2	
på: f	ö->2	
på: Ö	p->1	
på?. 	(->1	
på?Ja	g->1	
påbju	d->1	
påbör	j->11	
pådra	g->1	
påfre	s->1	
påföl	j->4	
pågic	k->3	
pågå 	i->1	
pågåe	n->6	
pågår	 ->7	.->3	
pågåt	t->1	
pålag	o->1	
pålen	 ->1	
pålit	l->1	
påläg	g->1	
påmin	d->1	n->29	
påpek	a->50	
pår a	v->1	
pår h	a->1	
pår i	 ->1	
pår t	a->1	
pår, 	d->1	o->1	
påra 	f->1	l->1	
påran	d->1	
påras	,->1	
påren	 ->1	
pårni	n->2	
påsky	n->7	
påstr	i->1	
påstå	 ->4	,->2	e->7	r->4	s->2	t->1	
påtag	l->4	
påtal	a->5	
påtry	c->3	
påtvi	n->4	
påver	k->37	
påvis	a->2	b->1	
pé oc	h->1	
péer 	a->1	i->1	m->1	s->1	
péer,	 ->2	
péern	a->3	
pérys	 ->1	
pöke 	d->1	
pöke.	M->1	
pöken	 ->1	
pökst	ä->1	
qal f	ö->1	
qal ä	r->1	
qua n	o->2	
qual 	D->1	h->1	s->2	v->1	ä->1	
qual"	 ->1	
qual,	 ->1	
que k	a->1	
que, 	s->1	
ques 	D->3	e->1	
ques"	.->1	
quier	d->1	
quins	 ->1	
quiol	a->1	
quisi	t->1	
quita	 ->1	
quo s	o->1	
quo, 	d->1	
quqal	 ->2	
r "Ku	l->1	
r "an	g->2	
r "fo	r->1	
r "in	l->1	
r "kr	o->1	
r "na	t->1	
r "öv	e->1	
r (C5	-->4	
r (FI	P->1	
r (ar	t->1	
r (i 	d->1	
r - 1	9->2	
r - a	n->2	r->1	t->6	v->2	
r - c	e->1	
r - d	e->11	o->1	
r - e	l->2	n->2	x->1	
r - f	ö->2	
r - g	ö->1	
r - h	a->2	u->1	
r - i	 ->2	d->1	n->5	
r - j	a->1	
r - k	o->4	
r - l	å->1	
r - m	e->2	
r - n	y->1	ä->1	
r - o	c->9	
r - s	e->1	i->1	k->1	n->1	o->3	t->1	å->2	
r - t	i->1	
r - u	t->1	
r - v	e->1	i->2	
r - ä	r->2	v->4	
r - ö	v->1	
r -, 	a->1	
r 1 4	0->1	
r 1 f	r->1	
r 1,2	 ->1	
r 1,4	 ->1	
r 1/3	 ->1	
r 10 	e->1	m->1	p->1	
r 100	 ->1	
r 12 	f->1	
r 124	4->1	
r 130	 ->1	
r 15 	a->1	p->1	
r 167	 ->1	
r 174	 ->1	
r 176	2->2	
r 192	3->1	
r 193	0->1	
r 197	6->1	
r 198	2->1	6->1	
r 199	0->1	1->1	2->1	4->1	6->9	7->13	8->9	9->32	
r 2 b	l->1	
r 20 	e->1	g->1	m->1	å->1	
r 200	 ->1	0->41	1->1	2->6	3->1	4->1	6->6	7->1	
r 201	0->1	2->1	
r 25 	g->1	
r 262	 ->1	
r 27 	p->2	
r 28 	f->1	
r 29 	d->1	f->1	l->1	
r 3 0	0->1	
r 3-4	 ->1	
r 30 	f->1	p->1	
r 31 	f->1	
r 32 	m->1	
r 32.	J->1	
r 33 	0->1	f->1	
r 332	,->1	
r 35 	f->1	m->1	
r 36 	f->1	
r 37 	f->1	
r 38 	f->1	
r 39 	f->1	
r 4 0	0->1	
r 40 	f->1	p->1	å->2	
r 41 	f->1	
r 42 	f->1	
r 43.	F->1	
r 44 	f->1	
r 45 	f->1	
r 46 	o->1	
r 5 f	r->1	
r 5 m	i->1	
r 5 å	r->1	
r 5,8	 ->1	
r 50 	0->1	p->1	
r 6 f	r->1	
r 60 	f->1	
r 7 g	r->1	
r 7 p	r->1	
r 7.F	r->1	
r 73,	9->1	
r 75 	m->1	
r 76 	p->1	
r 8 f	r->1	
r 80 	e->1	p->2	å->1	
r 81 	p->1	
r 9 f	r->1	
r 90 	d->1	p->1	
r 97.	S->1	
r 97/	9->1	
r Agr	i->1	
r Ala	v->1	
r Alb	e->1	
r Als	a->1	
r Alt	e->5	
r Amo	k->2	
r Ant	ó->1	
r Ara	f->1	
r Azo	r->1	
r BNI	 ->1	
r BNP	 ->1	
r BSE	-->1	
r Bar	a->2	n->10	ó->1	
r Bel	g->1	
r Ber	e->5	
r Bis	c->1	
r Bol	k->1	
r Bou	r->2	
r Bow	e->2	
r Bre	t->3	
r Bro	k->2	
r Bry	s->1	
r CEN	 ->1	
r CSU	:->1	
r Cen	t->2	
r Coc	a->1	
r Con	s->1	
r Cox	 ->1	!->1	,->1	
r Dan	m->3	
r Deu	t->1	
r Dor	i->1	
r Duh	a->1	
r ECH	O->1	
r EG-	d->2	k->3	
r EG.	V->1	
r EG:	s->1	
r EMU	,->1	:->1	
r EU 	i->2	
r EU,	 ->1	
r EU-	f->1	i->1	m->1	v->1	
r EU.	F->1	V->1	
r EU:	s->9	
r Egy	p->1	
r Ehu	d->1	
r Eko	n->1	
r Els	t->1	
r Eri	k->3	
r Eur	o->112	
r Eva	n->3	
r Exx	o->1	
r FN.	H->1	
r FN:	s->2	
r FPÖ	-->2	
r Far	o->1	
r Fin	l->1	
r Flo	r->1	
r FoU	,->1	
r Fol	k->1	
r Fra	s->1	
r Fru	t->1	
r För	e->6	
r GAS	P->1	
r Gam	a->2	
r Gen	è->1	
r Gol	a->1	f->1	l->1	
r Gom	e->1	
r Gra	ç->1	
r Gre	k->1	
r Gus	p->1	
r Gut	e->1	
r Hai	d->1	
r Hel	s->1	
r Him	a->1	
r Hän	s->2	
r I o	c->1	
r I-p	r->1	
r II 	i->1	
r II-	p->2	
r III	 ->1	
r IMO	.->1	
r INT	E->1	
r Int	e->2	
r Isr	a->5	
r Ita	l->1	
r Jap	a->1	
r Jon	c->2	
r Jos	p->1	
r Jör	g->2	
r Kan	t->3	
r Kin	a->1	n->10	
r Koc	h->1	
r Kos	o->1	
r Kou	c->1	
r Kul	t->2	
r Kum	a->1	
r Kvi	n->1	
r Kyo	t->1	
r Laa	n->7	
r Lan	g->3	
r Lei	n->1	
r Lis	s->1	
r Lot	h->2	
r Lux	e->1	
r Lyn	n->2	
r Maa	s->2	
r Mar	g->1	i->1	
r Mel	l->1	
r Mon	t->16	
r Mor	a->1	
r Nat	o->1	
r Ned	e->1	
r Nie	l->1	
r Nik	i->2	
r Nog	u->1	
r OFS	R->1	
r OLA	F->2	
r Ora	n->1	
r Osl	o->1	
r PPE	-->1	
r PVC	.->1	
r Pac	k->1	
r Pal	a->2	e->1	
r Pap	a->1	
r Pat	t->18	
r Poe	t->3	
r Poh	j->1	
r Pom	é->1	
r Pon	n->1	
r Poo	s->1	
r Por	t->3	
r Pre	u->1	
r Pro	d->1	
r REP	 ->1	
r Rap	k->1	
r Ras	c->1	
r Red	i->2	
r Rhô	n->1	
r Rot	h->1	
r Rus	h->1	
r Råd	e->1	
r Sav	e->2	
r Sch	r->3	ö->1	ü->2	
r Sea	t->1	
r Seg	n->1	u->1	
r Sei	x->2	
r Sha	r->1	
r Sko	t->1	
r Sol	a->1	b->1	
r Spe	r->1	
r Swo	b->1	
r Syr	i->2	
r São	 ->1	
r Tac	i->1	
r Tam	m->1	
r Tan	g->1	
r Tes	a->1	
r The	a->1	
r Tib	e->6	
r Tor	r->1	
r Tsa	t->2	
r Tur	k->4	
r UCL	A->1	
r UNM	I->1	
r USA	 ->1	
r USD	 ->1	
r Urq	u->1	
r Vit	o->5	
r Vol	k->1	
r WTO	?->1	
r Wal	e->2	l->1	
r Was	h->1	
r Wyn	n->1	
r [SE	K->1	
r abs	o->13	u->1	
r acc	e->6	
r adm	i->1	
r age	r->1	
r aid	s->1	
r akt	a->2	i->2	u->7	ö->1	
r ald	r->9	
r all	 ->5	a->92	d->11	i->2	m->13	o->1	r->1	t->145	v->12	
r amb	i->3	
r ame	r->1	
r ana	 ->1	l->3	m->4	
r anb	u->1	
r and	 ->1	e->2	r->22	
r anf	ö->2	
r ang	e->5	å->4	
r anh	ä->1	
r ank	l->1	
r anl	e->4	ö->1	
r anm	ä->3	
r ann	a->13	
r ano	n->2	r->1	
r ans	a->2	e->14	j->7	l->8	p->2	t->7	v->43	å->1	ö->1	
r ant	a->18	i->1	o->3	
r anv	ä->18	
r arb	e->35	
r arr	a->1	
r art	i->7	
r as"	.->1	
r asy	l->4	
r att	 ->1975	,->2	e->1	r->1	
r auc	t->1	
r av 	"->1	-->1	5->1	C->1	E->6	G->1	H->2	W->1	a->9	b->2	c->2	d->41	e->10	f->13	g->2	h->5	i->3	k->13	l->8	m->7	n->1	o->5	r->1	s->31	t->4	u->2	v->2	y->1	ö->1	
r av.	M->1	
r avb	r->2	
r avd	e->1	
r avf	a->4	
r avg	a->1	j->2	å->2	ö->9	
r avh	ä->1	
r avi	s->2	
r avl	a->1	ä->1	
r avs	a->3	e->8	i->16	k->2	l->5	t->5	ä->2	
r avt	a->2	
r avu	n->1	
r avv	e->2	i->2	
r bak	g->1	o->7	
r bal	a->1	
r ban	a->2	
r bar	a->29	b->1	
r bas	e->3	
r bea	k->5	
r bed	r->8	ö->5	
r bef	a->3	i->1	l->1	o->8	r->3	ä->1	
r beg	a->2	r->12	ä->8	å->2	
r beh	a->10	o->10	å->1	ö->11	
r bek	l->6	r->2	v->4	y->2	ä->2	
r bel	o->1	y->1	
r bem	ö->1	
r ber	 ->5	e->21	o->9	y->1	ä->9	ö->3	
r bes	k->4	l->21	t->14	v->1	ö->1	
r bet	a->9	e->2	o->3	r->6	y->19	ä->18	
r bev	a->4	i->9	
r bid	r->11	
r bif	a->1	
r bil	 ->1	.->1	a->14	d->5	e->1	i->2	l->1	p->1	t->2	
r bin	d->1	
r bis	t->6	
r bju	d->1	
r bl.	a->2	
r bla	m->1	n->5	
r bli	 ->6	,->1	r->8	v->16	
r blo	m->2	
r bly	,->1	g->1	
r bom	b->3	
r bor	 ->1	d->3	t->6	
r bos	a->2	t->1	
r bot	t->1	
r bov	e->1	
r bra	 ->10	!->1	,->6	.->4	
r bre	d->1	
r bri	s->13	t->2	
r bro	m->1	t->6	
r bru	k->1	t->1	
r bry	t->1	
r brå	d->4	
r brö	d->2	
r bud	g->20	s->1	
r bus	s->1	
r byg	g->6	
r byr	å->2	
r byx	f->1	
r bär	 ->1	
r bäs	t->3	
r bät	t->12	
r båd	a->2	e->9	
r böj	t->1	
r bör	 ->22	d->1	j->6	
r cap	i->10	
r cen	t->4	
r cho	c->1	k->1	
r cir	k->3	
r cit	a->1	e->1	
r civ	i->3	
r cop	y->1	
r cor	p->1	
r dag	,->1	.->1	e->4	o->1	s->8	
r dan	s->2	
r dat	u->1	
r de 	1->2	9->1	a->19	b->14	c->1	d->7	e->28	f->35	g->16	h->10	i->18	k->30	l->4	m->29	n->22	o->11	p->12	r->13	s->61	t->19	u->5	v->15	y->4	ä->5	å->10	ö->5	
r de,	 ->2	
r deb	a->32	
r dec	e->3	
r def	i->5	
r del	 ->16	a->9	e->3	s->1	t->9	
r dem	 ->30	,->4	.->9	?->1	a->1	o->13	
r den	 ->362	,->3	.->2	n->102	s->2	
r der	a->27	
r des	s->110	t->1	
r det	 ->913	!->1	,->7	.->17	a->6	s->1	t->124	
r dia	l->1	
r dip	l->1	
r dir	e->12	
r dis	c->2	k->21	p->1	t->1	
r dit	 ->2	
r div	e->1	
r dju	n->1	p->7	r->1	
r djä	r->1	
r doc	k->33	
r dok	u->2	
r dol	l->6	
r dom	a->2	s->5	
r dra	 ->1	b->7	g->1	m->2	r->1	s->1	
r dri	f->1	v->1	
r dro	g->1	
r du 	m->1	ä->1	
r dub	b->2	
r dug	a->1	
r dum	h->1	
r dyk	e->1	
r dyn	a->1	
r där	 ->23	!->1	,->1	.->3	e->3	f->71	h->1	i->1	m->1	
r då 	E->1	a->5	d->3	i->3	j->2	m->2	o->1	s->3	v->1	ö->1	
r dål	i->7	
r död	.->1	a->2	
r döl	j->2	
r dör	r->2	
r döt	t->1	
r ecu	 ->1	,->1	
r ed 	g->1	
r eff	e->12	
r eft	e->34	
r ege	n->16	
r egn	a->1	
r ego	i->1	
r ej 	a->1	b->1	i->1	k->1	n->1	
r ej,	 ->1	
r ej.	E->1	R->1	
r eko	l->1	n->26	s->1	
r ele	k->1	m->1	
r ell	e->59	
r elv	a->1	
r eme	l->28	
r emo	t->9	
r en 	"->1	R->1	a->35	b->20	c->3	d->29	e->30	f->59	g->36	h->14	i->11	j->2	k->35	l->14	m->57	n->19	o->23	p->12	r->28	s->66	t->14	u->17	v->36	y->1	ä->3	å->6	ö->15	
r en.	E->1	
r ena	d->1	t->1	
r enb	a->4	
r end	a->11	e->1	
r ene	r->15	
r eng	a->2	e->1	
r enh	e->4	ä->5	
r eni	g->2	
r enk	e->4	l->1	
r enl	i->20	
r eno	r->6	
r ens	 ->2	a->3	e->2	k->1	t->1	
r er 	-->1	a->8	b->1	d->3	e->2	f->2	i->1	l->1	o->4	p->1	r->1	s->2	t->4	u->1	v->2	
r er,	 ->10	
r er.	J->3	O->1	
r era	 ->7	
r erf	a->2	
r erh	å->2	
r eri	n->2	
r erk	ä->4	
r ers	a->1	ä->1	
r ert	 ->9	
r eta	b->4	
r etn	i->1	
r ett	 ->305	,->1	.->2	
r eur	o->31	
r evi	g->3	
r exa	k->1	m->1	
r exc	e->1	
r exe	m->7	
r exi	s->1	
r exp	e->7	
r ext	r->9	
r fac	k->1	
r fak	t->15	
r fal	l->21	s->1	
r fam	i->1	
r fan	t->1	
r far	a->3	l->9	t->7	
r fas	c->1	t->14	
r fat	t->7	
r fed	e->1	
r fel	 ->3	!->1	,->1	.->2	a->2	r->1	
r fem	 ->4	t->1	
r fic	k->2	
r fin	a->12	n->21	
r fis	k->7	
r fjo	r->1	
r fla	g->1	
r fle	r->16	x->1	
r fli	t->1	
r flo	d->2	
r fly	g->2	k->2	t->3	
r flä	k->1	
r fod	e->3	
r fol	k->7	
r fon	d->1	
r for	d->5	m->6	s->5	t->33	
r fra	k->1	m->95	n->3	
r fre	d->8	s->2	
r fri	 ->1	a->2	g->1	h->11	v->2	
r fru	k->1	
r frä	c->1	m->13	
r frå	g->68	n->87	
r ful	l->17	
r fun	d->2	g->3	k->1	n->3	
r fyl	l->1	
r fyr	a->2	
r fys	i->1	
r fär	r->1	
r fäs	t->1	
r få 	d->1	e->1	f->1	k->2	l->1	m->1	o->1	v->1	ä->1	
r få,	 ->2	
r få.	V->1	
r får	 ->12	
r fåt	t->28	
r fög	a->1	
r föl	j->14	
r för	 ->417	,->5	.->4	a->4	b->16	d->16	e->81	f->7	h->17	k->7	l->15	m->7	n->11	o->7	p->5	r->6	s->73	t->12	u->11	v->17	ä->3	å->1	ö->3	
r gag	n->3	
r gam	l->1	
r gan	s->7	
r gar	a->4	
r ge 	a->1	e->1	
r gem	e->30	
r gen	a->3	d->1	e->2	o->50	t->6	
r ger	 ->2	
r ges	 ->2	
r get	t->12	
r gil	t->1	
r giv	a->1	e->11	i->2	
r gjo	r->49	
r gla	d->12	
r glo	b->1	
r glä	d->2	
r glö	m->4	
r god	 ->3	.->1	a->1	k->11	s->1	t->10	
r gol	v->1	
r got	t->1	
r gra	n->8	t->3	
r gri	p->1	
r gru	n->20	p->17	
r grä	n->13	
r grå	z->1	
r gud	s->2	
r gyn	n->3	
r gäl	l->5	
r gär	n->3	
r gå 	i->1	
r gån	g->4	
r går	 ->10	,->1	d->1	
r gåt	t->11	
r göm	m->1	t->1	
r gör	 ->7	a->18	
r ha 	e->5	f->1	h->1	i->1	m->3	n->1	t->1	u->2	
r had	e->1	
r haf	t->16	
r hak	a->1	
r hal	v->6	
r ham	b->1	n->2	
r han	 ->18	d->10	s->32	t->2	
r har	 ->108	,->2	.->1	m->1	
r hav	e->1	s->1	
r hed	e->1	r->1	
r hel	a->40	h->3	i->1	l->3	t->57	
r hem	m->5	
r hen	n->10	
r her	r->1	
r het	s->1	
r hin	d->2	
r his	t->5	
r hit	 ->1	t->11	
r hjä	l->9	r->1	
r hom	o->2	
r hon	 ->6	o->9	
r hop	p->1	
r hor	i->1	
r hos	 ->7	
r hot	a->4	b->1	e->1	
r hum	a->1	
r hun	d->2	
r hur	 ->34	u->2	
r huv	u->12	
r hys	e->1	t->1	
r häl	f->1	s->2	
r häm	m->1	
r hän	d->3	g->4	s->4	t->4	v->2	
r här	 ->24	,->1	.->1	;->1	?->1	e->1	m->1	
r häs	t->1	
r häv	d->3	
r hål	l->12	
r hår	d->1	t->1	
r hög	 ->1	,->1	e->1	l->1	r->2	s->2	t->4	
r höj	a->1	
r hör	 ->2	a->1	d->1	t->11	
r i -	 ->1	
r i 2	0->1	
r i A	k->1	
r i B	e->1	i->1	r->2	
r i C	e->1	
r i D	a->1	u->1	
r i E	U->5	k->1	u->35	
r i F	r->2	ö->2	
r i I	r->2	t->1	
r i K	a->1	i->1	o->5	
r i L	o->1	
r i M	e->1	
r i O	L->1	
r i P	a->1	
r i S	c->1	k->1	t->3	
r i T	V->1	
r i U	S->2	
r i W	a->1	
r i a	i->1	l->8	n->9	r->5	t->4	v->1	
r i b	a->1	e->3	i->4	u->2	
r i d	a->47	e->72	i->1	r->1	
r i e	f->2	k->1	n->16	r->1	t->10	
r i f	j->2	o->6	r->13	ä->1	ö->23	
r i g	e->3	o->2	r->3	ä->1	å->3	
r i h	a->1	e->3	j->1	u->2	ä->1	
r i i	n->2	t->1	
r i j	o->1	u->1	
r i k	a->9	o->6	r->6	v->1	
r i l	a->1	i->1	
r i m	e->7	i->5	j->1	o->4	ä->1	å->5	
r i n	i->2	o->1	u->1	å->2	
r i o	c->3	f->3	m->4	r->2	u->1	
r i p	a->13	l->2	o->3	r->6	u->1	
r i r	a->1	e->5	i->1	u->1	ä->3	å->3	
r i s	a->5	i->19	j->5	k->2	l->2	m->1	t->16	y->2	
r i t	o->1	r->3	v->1	ä->2	
r i u	n->4	p->3	t->6	
r i v	a->5	e->2	i->8	ä->4	å->5	
r i Ö	V->1	s->6	
r i ä	k->1	
r i å	r->1	
r i ö	s->1	v->4	
r i.A	n->1	
r ian	s->1	
r ibl	a->3	
r ick	e->2	
r ide	a->1	n->4	
r idé	 ->1	n->1	
r ifr	å->6	
r ige	n->12	
r ign	o->1	
r iho	p->4	
r ikr	a->1	
r ill	a->1	e->2	o->1	
r imm	i->1	
r in 	2->1	F->1	d->1	i->5	k->1	o->1	s->1	
r inb	j->1	l->2	
r inc	i->2	
r ind	e->1	i->2	u->11	
r inf	l->1	o->2	r->2	ö->32	
r ing	a->12	e->35	i->2	å->10	
r ini	f->1	t->5	
r ink	l->1	o->3	ö->1	
r inl	e->9	ä->1	
r inn	a->5	e->15	o->1	
r ino	m->56	
r inr	e->6	i->3	y->1	ä->5	
r ins	a->3	e->4	i->1	k->2	l->1	t->11	
r int	a->4	e->414	o->1	r->23	y->1	
r inv	a->1	e->2	o->5	å->5	
r irl	ä->1	
r isc	e->1	
r isr	a->1	
r itu	 ->6	
r ivä	g->1	
r ja,	 ->1	
r jag	 ->278	,->6	
r jor	d->17	
r ju 	E->1	a->7	b->1	d->4	e->2	f->1	h->1	i->6	o->4	p->2	r->2	s->3	
r ju,	 ->2	
r jud	a->1	
r jul	f->1	
r jur	i->5	
r jus	t->16	
r jäm	f->2	l->1	s->2	
r jär	n->3	
r kal	l->5	
r kam	m->4	p->4	
r kan	 ->53	d->2	s->5	
r kap	i->1	
r kar	a->1	t->2	
r kat	a->10	e->2	
r kem	i->1	
r kla	r->28	
r kli	m->2	
r klo	c->1	k->4	
r kly	f->1	
r kna	p->5	
r knu	t->3	
r koa	l->1	
r kol	l->9	
r kom	 ->2	m->326	p->4	
r kon	c->4	f->4	k->44	s->28	t->16	v->2	
r kor	r->6	t->8	
r kos	t->14	
r kra	f->6	v->8	
r kre	t->1	
r kri	g->1	m->1	n->6	s->2	t->2	
r kry	s->1	
r krä	n->2	v->9	
r kub	i->1	
r kul	o->1	t->26	
r kun	n->15	s->1	
r kur	s->1	
r kus	t->3	
r kva	l->2	n->1	r->3	
r kve	s->2	
r kvi	n->10	
r kvä	l->2	
r käm	p->2	
r kän	d->2	n->2	s->3	t->6	
r kär	n->8	
r köl	d->1	
r kör	t->2	
r lag	e->3	l->5	s->9	t->36	
r lan	d->7	
r las	t->3	
r le 	p->1	
r led	a->25	e->2	n->2	s->3	
r leg	a->3	i->3	
r let	t->7	
r lev	e->2	n->1	
r lid	i->3	
r lig	g->7	
r lik	a->15	n->2	s->6	t->1	v->5	
r lis	t->2	
r lit	e->16	t->3	
r liv	 ->1	e->1	s->20	
r lob	b->1	
r log	i->2	
r lok	a->4	
r lot	t->1	
r lov	a->4	v->1	
r luf	t->1	
r lug	n->2	
r lur	a->1	
r lyc	k->17	
r lyf	t->1	
r lys	a->1	s->4	
r läc	k->1	
r läg	e->3	g->7	r->1	
r läk	a->1	
r läm	n->10	p->10	
r län	d->8	g->14	
r lär	t->1	
r läs	b->1	f->1	k->1	t->1	
r lät	t->9	
r lån	g->32	
r lås	t->1	
r låt	a->3	i->1	
r löj	e->2	
r lön	e->1	s->2	t->2	
r löp	t->4	
r lös	a->1	t->3	
r mai	n->3	
r maj	o->4	
r mak	t->1	
r mal	t->2	
r man	 ->167	,->3	a->1	d->3	l->1	
r mar	g->1	k->8	
r mas	s->1	t->1	
r mat	e->3	t->1	
r med	 ->199	b->35	d->6	e->3	g->2	h->1	i->2	k->1	l->34	v->10	
r mek	a->1	
r mel	l->18	
r men	 ->7	a->2	i->12	
r mer	 ->27	.->1	a->1	g->1	p->1	
r mes	t->3	
r met	a->2	o->2	
r mig	 ->87	!->1	,->9	.->2	
r mil	i->1	j->45	
r min	 ->23	a->9	d->12	i->7	n->2	o->1	s->9	u->3	
r mis	s->5	
r mit	t->10	
r mob	i->1	
r mod	e->3	i->2	
r mog	e->1	
r mon	o->1	
r mor	a->1	g->1	s->5	
r mot	 ->23	g->1	o->2	s->8	t->5	
r mun	t->1	
r mut	o->1	
r myc	k->104	
r myn	d->5	
r män	 ->3	g->3	n->23	s->3	
r mål	 ->5	e->3	s->1	
r mån	 ->1	a->4	d->1	g->34	
r mår	.->1	
r mås	t->45	
r möj	l->44	
r möt	e->2	
r nak	n->1	
r nam	n->1	
r nar	k->1	
r nat	i->14	u->30	
r ned	 ->4	m->1	s->1	
r neg	a->2	
r nej	,->2	.->1	
r nek	a->1	
r ner	 ->2	e->2	
r ni 	a->18	b->2	d->3	e->2	f->2	g->1	h->1	i->3	j->1	k->5	l->1	n->1	o->3	r->2	s->3	u->2	ä->1	
r ni,	 ->3	
r niv	å->2	
r nog	 ->2	a->1	
r nor	m->10	
r not	e->7	
r nu 	a->3	b->1	d->3	e->7	f->3	i->3	k->2	m->2	n->1	o->3	p->2	s->3	t->4	u->1	v->2	
r nu,	 ->2	
r nu.	J->1	L->1	
r nu:	 ->1	
r num	e->1	
r ny 	f->1	h->1	p->1	
r nya	 ->13	;->1	n->2	
r nyc	k->1	
r nyh	e->1	
r nyl	i->2	
r nyt	t->4	
r näm	l->2	n->11	
r när	 ->37	a->4	i->4	m->2	s->1	v->37	
r näs	t->12	
r någ	o->74	r->32	
r nåt	t->4	
r nöd	i->1	v->37	
r nöj	a->1	d->3	e->3	
r oac	c->7	
r oav	b->1	s->1	
r oba	l->1	
r obe	r->4	s->1	
r obs	e->1	
r och	 ->570	
r ock	s->161	u->1	
r oen	s->2	
r oer	h->5	s->1	
r oet	i->1	
r off	e->6	r->3	
r ofr	å->1	
r oft	a->23	
r ofu	l->2	
r ofö	r->4	
r ojä	m->1	
r okl	a->3	
r oku	n->1	
r ola	g->1	
r oli	k->9	
r olj	e->4	
r oly	c->4	
r olö	s->1	
r om 	-->1	3->1	A->2	G->2	H->1	K->1	a->44	b->9	d->40	e->31	f->16	g->1	h->12	i->7	j->1	k->9	l->5	m->12	n->5	o->3	p->3	r->7	s->18	t->4	u->3	v->9	ä->2	å->4	
r om,	 ->5	
r om.	D->1	E->1	I->1	O->1	S->2	
r omb	e->1	
r omf	a->8	l->1	o->1	å->1	
r omk	r->9	
r oml	a->1	
r omp	r->1	
r omr	å->9	ö->4	
r oms	o->1	t->1	
r omv	a->1	
r omö	j->3	
r onö	d->2	
r opi	n->1	
r ord	 ->2	.->1	:->1	e->8	f->13	n->3	
r ori	m->1	
r oro	 ->6	,->1	.->3	a->1	n->1	v->1	
r ors	a->5	
r orä	t->4	
r oss	 ->117	,->6	.->8	:->1	
r ost	r->1	
r osä	k->1	
r oså	r->1	
r oti	l->3	
r otr	o->1	
r otå	l->1	
r oum	b->1	
r oun	d->2	
r out	h->2	
r ova	n->1	
r ovä	d->1	
r oöv	e->1	
r pap	p->1	
r par	a->2	l->52	t->4	
r pas	s->3	
r pek	a->3	
r pen	g->9	n->2	
r per	 ->2	f->2	i->17	s->12	
r pes	s->1	
r pla	c->1	n->8	t->1	
r ple	n->2	
r pli	k->2	
r plu	s->1	
r pol	i->23	
r pos	i->9	
r pot	e->1	
r poä	n->1	
r pra	c->1	k->2	
r pre	c->9	s->7	
r pri	n->6	o->1	s->2	v->1	
r pro	b->22	c->3	d->10	g->14	j->4	t->2	v->1	
r prä	g->1	
r prö	v->2	
r pun	d->1	k->9	
r på 	-->3	2->2	9->1	A->1	B->1	E->2	H->1	P->1	R->1	a->47	b->8	c->1	d->52	e->28	f->11	g->12	h->4	i->5	k->15	l->5	m->8	n->7	o->10	p->6	r->7	s->31	t->7	u->5	v->17	y->1	Ö->1	ä->1	
r på,	 ->3	
r på.	E->1	J->1	N->1	
r påb	j->1	ö->3	
r påf	ö->1	
r pål	a->1	
r påm	i->2	
r påp	e->7	
r pås	t->1	
r påt	a->3	r->1	
r påv	e->4	i->2	
r rad	i->2	
r rak	a->2	
r ram	a->1	
r rap	p->4	
r ras	i->3	
r rat	i->5	
r rea	g->1	k->2	l->3	
r rec	y->1	
r red	a->34	o->1	
r ref	e->1	o->12	
r reg	e->37	i->29	l->5	
r reh	a->1	
r rej	ä->2	
r rek	o->7	
r rel	a->3	e->2	i->1	
r ren	a->1	t->3	
r rep	r->3	u->1	
r res	a->1	e->1	o->9	p->4	t->1	u->7	
r ret	r->2	
r rev	i->4	
r rig	o->1	
r rik	a->1	t->10	
r rim	l->4	
r rin	g->1	
r ris	k->13	
r rol	i->1	l->4	
r rop	e->1	
r ros	e->1	t->1	
r rui	n->1	
r rum	 ->2	
r run	t->1	
r rus	t->1	
r rut	t->1	
r ryc	k->1	
r räd	d->4	
r räk	e->1	n->6	
r rät	t->66	
r råd	?->1	a->1	e->33	g->1	s->14	
r rör	 ->1	a->6	e->1	l->2	t->1	
r rös	t->15	
r sad	e->2	
r sag	t->20	
r sak	,->1	e->3	n->5	
r sam	a->5	b->2	f->2	h->4	l->2	m->32	o->4	r->1	t->23	
r san	n->1	t->8	
r sat	s->2	t->4	
r se 	e->1	h->1	o->1	s->1	t->3	ö->1	
r sed	a->29	
r seg	l->2	r->1	
r sek	r->1	t->2	u->1	
r sen	a->10	s->1	t->3	
r ser	 ->5	i->1	
r ses	 ->1	
r set	t->9	
r sex	 ->3	t->1	
r sid	a->2	
r sig	 ->118	,->3	.->5	
r sik	t->1	
r sin	 ->30	a->26	n->1	s->1	
r sis	t->5	
r sit	t->16	u->10	
r sju	 ->1	k->1	n->1	
r sjä	l->28	t->1	
r sjö	f->1	
r ska	d->9	l->59	m->1	p->12	r->1	t->2	
r ske	p->1	t->5	
r ski	c->3	l->6	
r skj	u->5	
r sko	g->5	
r skr	i->6	o->7	ä->1	
r sku	l->23	t->1	
r sky	d->8	l->9	m->1	
r skä	l->4	r->1	
r skö	r->1	t->1	
r sla	g->3	
r slu	k->1	s->1	t->11	
r slä	p->3	
r smu	t->1	
r små	 ->6	,->1	f->1	
r sna	b->6	r->6	
r sne	d->2	
r snä	v->1	
r soc	i->4	
r sol	i->3	
r som	 ->632	,->3	l->1	
r sov	j->1	
r spa	n->3	
r spe	c->8	l->7	n->3	
r spi	l->1	
r spo	n->1	
r spr	i->4	
r spä	n->1	r->1	
r spå	r->1	
r sta	b->4	d->2	n->2	r->8	t->28	
r ste	g->2	l->1	n->1	
r sti	c->1	m->1	
r sto	d->1	l->3	p->3	r->49	
r str	a->4	i->3	u->9	y->2	ä->6	
r stu	d->1	m->1	n->1	
r sty	r->4	
r stä	l->12	n->1	
r stå	 ->2	e->1	l->5	n->6	r->5	t->3	
r stö	d->23	r->9	t->6	
r sub	s->5	
r sun	d->1	
r sva	g->5	r->6	
r svå	r->19	
r syd	ö->1	
r syf	t->4	
r sym	b->3	p->1	
r syn	 ->1	e->2	l->3	n->1	p->1	
r sys	s->24	t->2	
r säg	a->3	e->1	
r säk	e->46	r->2	
r säl	l->1	
r säm	r->1	
r sän	k->1	
r sär	k->1	s->36	
r sät	t->3	
r så 	a->15	b->1	e->1	f->2	i->1	k->5	l->4	m->7	n->3	p->1	s->12	t->1	u->1	v->4	ä->3	
r så,	 ->3	
r såd	a->10	
r sål	e->16	u->3	
r sås	o->4	
r såv	ä->7	
r söd	r->1	
r sön	d->3	
r t.e	x->3	
r ta 	d->3	e->1	h->4	m->1	
r tac	k->1	
r tag	i->26	
r tal	a->17	m->321	
r tan	k->4	
r tar	 ->2	
r tas	 ->2	
r tek	n->6	
r tem	p->2	
r ten	d->1	
r tex	t->2	
r tib	e->2	
r tid	 ->2	e->5	i->9	s->1	t->1	
r til	l->413	
r tio	 ->1	t->3	
r tit	e->1	t->1	
r tju	g->1	
r tjä	n->14	
r tob	a->1	
r tog	 ->1	s->1	
r tol	e->1	k->4	
r ton	 ->2	
r top	p->1	
r tor	d->1	k->1	v->1	
r tot	a->3	
r tra	f->2	n->23	s->1	
r tre	 ->6	d->6	m->1	t->2	
r tro	 ->1	.->1	l->2	n->1	r->5	t->5	
r try	c->2	g->1	
r trä	 ->1	d->2	f->2	p->1	t->2	
r trå	k->2	
r trö	t->1	
r tun	g->1	n->1	
r tur	i->3	
r tus	e->2	
r tve	k->2	t->1	
r tvi	n->5	v->3	
r tvu	n->5	
r tvä	r->3	
r två	 ->20	h->1	
r tyc	k->1	
r tyd	e->1	l->14	
r tyn	g->2	
r typ	e->11	
r tyv	ä->7	
r tän	k->6	
r tär	t->1	
r tät	a->1	
r tåg	o->1	
r und	a->7	e->57	r->3	
r ung	a->1	d->4	e->4	
r uni	o->44	v->1	
r upp	 ->17	.->2	b->1	e->22	f->12	g->7	h->10	k->1	l->3	m->17	n->8	r->14	s->9	t->5	v->1	
r ur 	b->1	d->1	e->2	i->1	m->2	
r urs	p->1	ä->1	
r urv	a->1	
r ut 	T->1	a->1	f->2	m->1	n->1	o->2	p->8	s->4	t->2	ö->2	
r ut,	 ->3	
r ut.	F->1	S->1	Ä->1	
r ut?	.->1	
r uta	n->50	r->1	
r utb	i->5	r->1	y->2	
r ute	 ->4	l->1	s->3	
r utf	a->1	o->1	r->3	ä->6	ö->9	
r utg	i->3	å->2	ö->3	
r uti	f->4	
r utk	o->1	r->1	
r utl	o->1	ö->1	
r utm	a->2	
r utn	y->4	
r uto	m->3	
r utp	r->1	
r utr	e->1	i->4	o->1	y->1	ä->1	
r uts	a->1	k->26	t->10	
r utt	a->4	j->1	o->1	r->3	ö->2	
r utv	e->34	i->8	ä->1	
r utö	k->1	v->6	
r vad	 ->36	
r vag	a->1	
r vak	a->1	s->3	u->1	
r val	 ->1	d->2	e->1	t->6	
r van	 ->5	
r var	 ->11	a->42	d->2	e->1	f->2	i->27	j->17	m->5	o->1	s->7	t->1	
r vat	t->2	
r vec	k->2	
r ved	e->1	
r vek	h->1	
r vel	a->1	
r vem	 ->1	
r ver	k->46	
r vet	 ->6	,->1	a->4	e->12	
r vi 	-->1	E->2	L->1	P->1	a->52	b->17	d->28	e->23	f->28	g->8	h->30	i->55	j->1	k->23	l->5	m->12	n->12	o->18	p->9	r->9	s->38	t->22	u->7	v->15	ä->8	ö->1	
r vi,	 ->5	
r vid	 ->21	a->3	h->1	s->1	t->5	
r vig	v->1	
r vik	t->64	
r vil	a->1	j->10	k->16	l->22	s->1	
r vin	s->1	
r vir	k->1	
r vis	a->16	e->1	i->1	s->25	t->1	
r vit	b->8	t->1	
r vol	u->1	
r von	 ->1	
r vot	e->1	
r vun	n->2	
r vux	n->1	
r väc	k->5	
r väg	 ->3	b->1	n->1	
r väl	 ->13	d->9	f->1	j->2	k->8	m->1	s->3	t->2	
r vän	l->1	s->1	t->5	
r vär	d->11	r->1	t->3	
r väs	e->3	t->1	
r väx	l->1	t->1	
r vål	l->1	
r vår	 ->36	a->33	t->20	
r yng	r->1	
r ypp	a->1	
r yrk	a->1	e->1	
r ytt	e->15	r->1	
r ÖVP	 ->1	
r Öst	e->7	
r ägn	a->5	
r ägt	 ->3	
r äld	r->4	
r ämn	a->3	
r än 	1->4	3->1	F->1	a->3	b->1	d->5	e->12	f->3	g->1	h->1	k->1	l->1	m->3	n->3	o->1	p->1	r->1	s->3	t->4	v->9	
r änd	a->1	r->21	å->16	
r äng	s->1	
r änn	u->17	
r är 	E->1	F->1	a->11	b->5	c->1	d->37	e->10	f->9	g->1	h->3	i->7	j->2	k->1	l->3	m->5	n->10	o->9	p->1	r->1	s->12	t->3	u->3	v->8	ö->1	
r ära	n->2	
r äre	n->1	
r ärl	i->2	
r äve	n->35	
r å a	n->1	
r å e	n->1	
r åkl	a->1	
r åla	g->1	
r år 	1->12	2->11	a->1	f->1	s->2	
r år,	 ->1	
r åre	n->5	t->2	
r årt	u->1	
r åsa	m->1	
r åsi	k->3	
r åsk	å->1	
r åst	a->1	
r åt 	a->1	d->3	e->1	r->2	s->1	
r åta	 ->1	g->2	l->1	
r åte	r->33	
r åtf	ö->1	
r åtg	ä->6	
r åtm	i->3	
r åts	k->2	
r ått	a->2	
r öar	n->1	
r öde	l->1	
r ögo	n->7	
r öka	d->6	r->1	t->6	
r öns	k->7	
r öpp	e->13	n->3	
r öre	g->2	
r öst	e->2	r->1	
r öva	t->1	
r öve	r->92	
r övr	i->29	
r! 19	9->1	
r! Av	s->1	
r! Be	r->1	
r! Bl	a->1	
r! Ce	n->1	
r! De	 ->2	n->5	t->12	
r! Di	r->1	
r! Ef	t->4	
r! Er	a->1	
r! Et	t->1	
r! Eu	r->4	
r! Fö	r->8	
r! Go	t->1	
r! Gr	u->1	
r! Hi	t->1	
r! I 	b->1	d->5	e->1	m->1	u->1	
r! Ja	,->1	g->24	
r! Jä	m->1	
r! Ka	r->1	
r! Lå	t->4	
r! Me	d->1	
r! Ni	 ->1	
r! Nä	r->2	
r! Nå	g->1	
r! Om	 ->1	
r! PP	E->1	
r! På	 ->1	
r! So	m->3	
r! Ta	c->2	
r! Ti	l->3	
r! Un	d->2	
r! Vi	 ->8	d->1	s->1	
r! Vå	r->1	
r! Äv	e->3	
r! År	l->1	
r!"De	t->1	
r!"Om	 ->1	
r!.He	r->1	
r!De 	a->1	f->1	s->1	
r!Det	 ->3	t->1	
r!Eft	e->1	
r!Eri	k->1	
r!Jag	 ->5	
r!Med	 ->1	
r!Min	 ->1	
r!Myc	k->1	
r!Til	l->1	
r!Vi 	f->1	s->1	
r" ha	r->1	
r" må	s->2	
r" oc	h->1	
r" so	m->2	
r"), 	v->1	
r", s	o->1	
r".De	t->1	
r".Ja	g->1	
r".Om	 ->1	
r) Bo	r->1	
r) Vi	 ->1	
r) oc	h->3	
r).)B	e->1	
r)? H	a->1	
r)Fru	 ->2	
r)Jag	 ->1	
r)Kon	r->1	
r)Tac	k->1	
r, "n	e->1	
r, (B	r->1	
r, 16	6->1	
r, Bu	s->1	
r, Eu	r->1	
r, Ga	r->1	
r, Ma	r->1	
r, Pa	l->1	
r, Th	y->1	
r, Ty	s->1	
r, Wa	f->1	
r, ac	c->1	
r, ad	m->1	
r, al	b->1	l->8	
r, an	f->1	s->4	t->1	
r, ar	b->1	
r, at	t->37	
r, av	 ->5	
r, ba	r->1	
r, be	r->4	s->1	
r, bi	l->1	
r, bl	.->3	a->2	i->1	
r, bo	r->1	
r, br	ö->1	
r, bä	s->3	
r, bå	d->3	
r, de	 ->3	l->1	n->1	t->14	
r, di	f->1	
r, dj	u->1	
r, dv	s->8	
r, dä	r->11	
r, då	 ->7	
r, dö	d->1	
r, ef	t->10	
r, el	e->1	l->4	
r, en	 ->11	d->1	l->5	
r, er	b->1	
r, et	t->3	
r, ex	e->1	i->1	
r, fi	n->2	
r, fo	r->1	
r, fr	a->3	u->8	å->5	
r, få	r->1	
r, fö	r->36	
r, ga	m->1	
r, ge	m->3	n->3	r->1	
r, gy	n->1	
r, gå	 ->1	
r, gö	r->2	
r, ha	m->1	n->1	r->8	
r, he	l->1	r->16	t->1	
r, ho	t->1	
r, hu	r->1	v->1	
r, hä	r->2	
r, hö	j->1	
r, i 	d->3	e->6	f->1	l->1	m->1	p->2	s->4	t->1	
r, ib	l->1	
r, ic	k->1	
r, in	b->2	d->1	f->1	g->1	k->5	n->2	o->1	r->1	s->1	t->14	
r, ja	g->10	
r, jä	r->2	
r, ka	d->1	n->6	
r, ko	l->5	m->13	s->1	
r, kr	a->1	o->1	ä->2	
r, ku	l->1	
r, kä	r->18	
r, la	d->1	
r, le	d->2	
r, li	k->7	v->1	
r, lo	k->1	
r, lä	m->1	s->1	
r, lå	n->2	
r, ma	k->1	n->1	t->1	
r, me	d->16	n->57	r->2	
r, mi	l->1	n->8	s->1	
r, mo	n->1	r->1	
r, my	c->1	n->1	
r, mä	n->5	
r, må	 ->1	s->5	
r, na	t->1	
r, ne	d->1	k->1	
r, ni	 ->2	
r, no	g->1	
r, ny	 ->1	a->1	
r, nä	m->2	r->8	s->1	
r, nå	g->6	
r, oa	v->1	
r, oc	h->110	k->1	
r, ol	y->1	
r, om	 ->17	
r, or	d->1	e->1	g->2	
r, pe	r->1	
r, pl	u->1	
r, pr	e->3	i->2	
r, på	 ->7	
r, re	g->1	k->2	
r, ro	m->1	
r, rä	k->1	t->2	
r, rå	d->1	
r, rö	s->1	
r, sa	d->1	k->1	m->6	
r, se	 ->1	
r, si	n->2	
r, sj	u->1	
r, sk	a->2	i->1	u->2	
r, sm	a->1	
r, sn	a->1	e->2	
r, so	l->1	m->68	
r, sp	e->1	
r, st	a->2	ö->1	
r, sv	a->2	
r, sä	k->1	r->6	
r, så	 ->14	s->2	v->4	
r, ta	k->1	l->1	
r, ti	l->16	t->1	
r, tj	ä->3	
r, tr	a->3	e->1	o->2	
r, tu	r->1	
r, ty	 ->1	v->1	
r, un	d->6	g->4	
r, up	p->4	
r, ut	a->23	b->3	r->1	v->2	
r, va	d->2	n->1	r->2	t->1	
r, ve	r->1	t->2	
r, vi	 ->7	l->25	
r, vä	c->1	r->3	
r, vå	r->1	
r, än	 ->1	d->2	
r, är	 ->16	a->10	
r, äv	e->8	
r, åt	 ->1	a->1	e->4	m->1	
r, öv	e->1	
r- oc	h->4	
r- so	m->1	
r-bil	a->1	
r-kom	m->1	
r-nat	i->1	
r-pro	g->11	
r-reg	i->1	
r. (F	R->1	
r. Al	l->1	
r. De	n->2	t->5	
r. Ef	t->1	
r. En	 ->3	
r. Eu	r->1	
r. Fr	ä->1	
r. He	r->1	
r. Ja	g->2	
r. Ma	n->1	
r. Me	n->2	
r. Ni	 ->1	
r. Sy	r->1	
r. Så	 ->1	
r. Ti	l->1	
r. Vi	 ->1	
r. Vå	r->1	
r. in	t->1	
r. Än	n->1	
r.(Ap	p->1	
r.(IT	)->1	
r.(Li	v->1	
r.) H	e->1	
r.)Sä	k->1	
r.- (	D->1	P->2	
r.- H	e->1	
r.. (	E->2	F->2	
r..(E	N->2	
r..(N	L->1	
r...(	T->1	
r...H	e->1	
r..He	r->1	
r..Vi	 ->1	
r.90 	p->1	
r.All	a->1	d->1	t->1	
r.Alt	e->1	
r.Ame	r->1	
r.Ant	a->1	
r.Att	 ->3	a->1	
r.Av 	a->2	d->2	
r.Bar	a->2	
r.Bed	r->1	ö->1	
r.Bef	o->1	
r.Bet	r->1	ä->3	
r.Bla	n->2	
r.Bos	ä->1	
r.Bre	t->1	
r.CSU	:->1	
r.Dag	e->1	
r.De 	a->4	d->1	f->5	g->1	h->2	k->3	m->1	n->2	s->6	t->1	u->1	v->2	ä->1	å->1	
r.Den	 ->34	n->8	
r.Des	s->8	
r.Det	 ->110	t->35	
r.Dir	e->1	
r.Dom	s->1	
r.Där	 ->2	e->3	f->7	i->1	u->1	
r.Då 	v->1	ä->1	
r.EU-	k->1	o->1	
r.Eft	e->5	
r.En 	a->1	d->2	r->2	s->3	v->2	
r.Enb	a->1	
r.Enl	i->3	
r.Erf	a->1	
r.Ett	 ->6	
r.Eur	o->7	
r.Exe	m->1	
r.FPÖ	:->1	
r.Fem	 ->1	
r.Fol	k->1	
r.Fra	m->1	
r.Fre	d->1	
r.Fri	h->1	
r.Fru	 ->7	
r.Frå	g->3	
r.Får	 ->1	
r.För	 ->34	e->1	h->2	m->1	p->1	s->3	t->1	
r.Gem	e->2	
r.Gen	o->5	
r.Gör	 ->1	
r.Han	s->1	
r.Her	r->25	
r.Hur	 ->2	
r.Huv	u->1	
r.Hän	d->2	
r.Här	 ->5	o->1	
r.I E	u->1	
r.I H	e->1	
r.I I	r->2	t->1	
r.I R	a->1	
r.I a	l->1	n->1	
r.I b	e->1	
r.I d	e->6	
r.I e	g->1	n->2	
r.I f	ö->1	
r.I g	å->1	
r.I j	u->1	
r.I m	å->1	
r.I r	e->2	ä->1	
r.I s	a->1	t->1	
r.I v	i->2	å->1	
r.Ind	u->1	
r.Ing	e->3	
r.Ino	m->3	
r.Inr	e->1	
r.Int	e->1	
r.Ita	l->1	
r.Jac	q->1	
r.Jag	 ->118	
r.Kan	s->2	
r.Kar	l->1	
r.Kin	n->1	
r.Kod	e->1	
r.Kom	m->21	
r.Kon	k->2	s->2	v->1	
r.Kra	v->1	
r.Kvi	n->1	
r.Kär	n->1	
r.Lan	g->1	
r.Lik	a->1	s->2	
r.Lyc	k->1	
r.Låt	 ->6	
r.Man	 ->5	
r.Mar	k->1	
r.Med	 ->5	a->1	l->1	
r.Mel	l->1	
r.Men	 ->20	
r.Mer	 ->1	
r.Min	 ->3	a->1	
r.Myl	l->1	
r.Män	n->1	
r.Nat	u->4	
r.Ni 	k->1	
r.Niv	å->1	
r.Nu 	h->1	
r.Nya	 ->1	
r.När	 ->10	
r.Någ	o->1	
r.Obe	r->1	
r.Och	 ->7	
r.Ock	s->1	
r.Om 	a->1	d->8	e->1	f->1	g->1	i->1	m->2	v->1	
r.Omr	ö->1	
r.Ord	f->1	
r.Oro	v->1	
r.Par	l->2	
r.Pla	s->1	
r.Pro	b->3	
r.Pun	k->1	
r.På 	m->1	s->2	
r.Ras	i->1	
r.Red	a->1	
r.Ref	o->1	
r.Ren	t->1	
r.Rev	i->2	
r.Ris	k->1	
r.Räk	n->1	
r.Råd	e->3	
r.Sam	h->1	m->2	t->2	
r.Sed	a->2	
r.Sku	l->1	
r.Slu	t->2	
r.Som	 ->6	l->1	
r.Sta	t->1	
r.Sto	r->1	
r.Str	u->1	
r.Stö	d->2	
r.Så 	b->1	d->1	
r.Såd	a->1	
r.Sål	e->2	
r.Tac	k->5	
r.Ter	r->1	
r.Til	l->15	
r.Tro	t->1	
r.Ty 	v->1	
r.Tyv	ä->2	
r.Und	e->6	
r.Uni	o->1	
r.Ute	s->1	
r.Vad	 ->8	
r.Val	e->1	
r.Var	 ->1	f->3	j->1	
r.Vem	 ->2	
r.Vi 	a->6	b->7	f->4	g->1	h->19	i->2	k->10	l->1	m->16	s->4	v->11	ä->4	
r.Vid	a->1	
r.Vis	s->2	
r.Vår	 ->3	t->2	
r.kom	m->1	
r.Änd	r->3	å->2	
r.Är 	d->3	
r.Äve	n->5	
r.Å a	n->2	
r.ÖVP	 ->1	
r: "J	a->1	
r: An	m->1	
r: De	s->1	t->2	
r: Fi	n->1	
r: Fr	i->1	
r: Fö	r->1	
r: In	g->1	
r: Kä	n->1	
r: Om	 ->1	
r: På	 ->1	
r: Vi	 ->2	
r: an	g->1	t->1	
r: at	t->2	
r: de	n->3	t->5	
r: en	 ->2	
r: fö	r->3	
r: hu	r->1	
r: in	o->1	
r: ko	m->1	
r: nu	 ->1	
r: om	 ->1	
r: op	e->1	
r: ti	l->1	
r: ut	n->1	
r: ve	m->1	
r: vi	 ->3	l->1	
r: Är	 ->1	
r; at	t->1	
r; de	s->2	t->1	
r; då	 ->1	
r; en	 ->1	
r; i 	F->1	
r; in	l->1	
r; ja	g->1	
r; me	n->1	
r; oc	h->2	
r; vi	 ->1	d->1	
r?, r	å->1	
r?- (	P->1	
r?. (	E->1	
r?Bor	d->1	
r?Det	 ->2	
r?Där	f->1	
r?Eur	o->1	
r?Fru	 ->1	
r?Frå	g->1	
r?Har	 ->2	
r?Her	r->3	
r?Hur	 ->1	
r?I e	r->1	
r?I m	e->1	
r?Jag	 ->3	
r?Kan	s->1	
r?Kom	m->2	
r?Men	 ->2	
r?Nat	u->1	
r?Ni 	k->1	
r?Näs	t->1	
r?På 	d->1	
r?Som	 ->1	
r?Tac	k->1	
r?Vem	 ->1	
r?Vi 	m->1	t->1	
r?Är 	d->2	
r?Äve	n->1	
rHerr	 ->1	
rJag 	g->1	
rMed 	d->1	
rNäst	a->2	
ra "b	a->1	
ra "u	t->1	
ra - 	g->1	k->1	l->1	o->3	
ra 1 	p->1	
ra 10	 ->1	
ra 15	 ->1	
ra 16	 ->1	
ra 2 	p->1	
ra 25	 ->1	
ra 5 	m->1	
ra 55	 ->1	
ra 70	 ->1	
ra At	l->1	
ra Ba	r->1	
ra Da	n->1	
ra EE	G->1	
ra EU	 ->3	-->1	
ra Eu	r->13	
ra FN	:->1	
ra Fr	a->1	
ra In	t->1	
ra Is	r->2	
ra Je	r->1	
ra Li	b->2	
ra Lo	u->1	
ra Ri	i->1	
ra Ro	m->1	
ra Ty	s->2	
ra ad	m->1	
ra af	f->2	
ra ag	g->1	
ra ak	t->2	
ra al	k->1	l->15	t->2	
ra am	b->3	
ra an	d->2	h->2	m->1	s->15	t->2	v->2	
ra ar	a->1	b->11	g->1	r->2	t->2	
ra as	p->4	y->1	
ra at	t->101	
ra au	t->1	
ra av	 ->45	g->1	s->5	t->2	
ra ba	k->1	l->1	n->3	r->1	s->2	
ra be	d->4	f->3	g->3	h->5	k->1	l->3	r->5	s->9	t->15	u->1	v->1	
ra bi	d->1	l->3	n->1	t->1	
ra bl	i->2	
ra bo	s->1	
ra br	a->3	i->1	o->1	ä->1	
ra bu	d->1	
ra by	r->1	
ra bä	r->1	s->2	t->4	
ra bå	d->1	t->1	
ra bö	r->2	
ra ce	n->4	
ra da	g->8	t->1	
ra de	 ->36	b->2	l->21	m->14	n->73	r->4	s->16	t->94	
ra di	a->1	e->1	k->1	p->1	r->2	s->3	
ra dj	u->2	
ra do	k->1	
ra dr	a->2	ö->1	
ra du	m->1	
ra dy	r->1	
ra dä	r->1	
ra dö	d->1	
ra ef	f->7	t->1	
ra eg	n->7	
ra ek	o->5	
ra el	l->5	
ra em	o->1	
ra en	 ->117	,->1	d->1	e->37	h->4	k->3	l->3	s->2	
ra er	 ->18	,->1	f->2	i->1	k->1	
ra et	n->2	t->67	
ra eu	r->11	
ra ex	a->1	e->5	i->1	t->1	
ra fa	k->2	l->9	r->5	s->2	t->4	
ra fe	l->2	m->2	n->1	
ra fi	n->1	
ra fl	e->5	ö->1	
ra fo	r->6	
ra fr	a->11	e->1	u->1	å->41	
ra fu	l->4	
ra fä	r->1	
ra få	 ->3	
ra fö	l->4	r->159	
ra ga	n->1	
ra ge	m->9	n->11	
ra gi	v->5	
ra gj	o->1	
ra gl	a->1	ä->1	
ra go	d->4	
ra gr	a->2	u->18	ä->4	
ra gä	l->7	
ra gå	n->12	r->1	
ra gö	r->3	
ra ha	m->1	n->7	r->5	
ra he	l->13	m->3	n->2	r->1	t->1	
ra hi	n->1	s->1	t->1	
ra ho	n->4	p->1	r->1	
ra hu	n->1	r->12	s->1	v->2	
ra hä	l->1	r->5	
ra hå	l->5	
ra hö	g->2	
ra i 	D->1	E->2	F->1	I->1	K->1	L->2	R->1	a->1	b->1	d->7	e->6	f->5	g->1	h->1	k->1	l->1	m->3	r->1	s->3	t->1	v->1	ö->1	
ra ia	k->1	
ra ic	k->1	
ra id	e->1	é->2	
ra if	r->1	
ra ig	å->2	
ra ih	o->1	
ra il	l->2	
ra in	 ->4	d->1	f->5	g->1	i->3	l->4	n->2	o->2	r->1	s->13	t->13	v->4	
ra ja	g->1	
ra jo	b->1	
ra ju	l->1	s->1	
ra jä	m->2	
ra ka	m->2	n->4	p->1	t->3	
ra ke	d->1	
ra ki	l->1	
ra kl	a->7	i->1	
ra kn	u->1	
ra ko	l->65	m->30	n->31	r->8	s->3	
ra kr	a->1	e->2	i->3	o->1	ä->1	
ra ku	l->2	n->1	r->1	s->1	
ra kv	a->2	i->3	o->1	
ra kä	l->1	n->1	r->2	
ra la	b->1	g->7	n->5	
ra le	d->6	k->1	
ra li	k->7	t->2	v->5	
ra lo	k->2	
ra lä	g->2	m->4	n->21	r->1	t->1	
ra lö	f->1	n->1	s->2	
ra ma	j->1	k->2	r->2	t->1	
ra me	d->80	l->2	n->2	r->7	s->1	
ra mi	g->6	l->9	n->19	s->3	t->4	
ra mo	d->2	m->1	t->6	
ra my	c->21	n->1	
ra mä	n->7	
ra må	l->6	n->11	s->12	t->1	
ra mö	j->10	
ra na	i->1	t->8	
ra ne	d->1	g->1	
ra nu	?->1	
ra ny	a->7	c->2	h->3	t->4	
ra nä	m->6	r->6	s->1	t->1	
ra nå	g->33	
ra nö	d->6	j->2	
ra ob	e->3	l->2	
ra oc	h->54	k->2	
ra of	f->2	ö->2	
ra ok	o->1	
ra ol	i->6	j->3	y->2	
ra om	 ->30	,->1	e->2	g->1	r->14	s->5	ö->1	
ra on	ö->1	
ra op	t->2	
ra or	d->22	e->1	g->1	o->2	s->3	
ra os	s->11	
ra ot	i->1	
ra pa	r->12	
ra pe	d->1	k->1	l->2	n->2	r->3	
ra pl	a->4	
ra po	l->14	r->1	s->3	
ra pr	a->3	e->1	i->7	o->26	
ra pu	b->1	n->12	
ra på	 ->41	.->1	p->1	s->1	
ra ra	p->10	
ra re	a->2	d->4	f->4	g->17	k->1	l->1	n->1	p->2	s->11	t->1	
ra ri	k->5	m->1	s->3	
ra ro	l->1	m->1	
ra ru	m->1	n->1	
ra rä	c->1	d->1	t->3	
ra rå	d->3	o->1	
ra rö	s->1	
ra sa	k->7	m->18	n->2	t->2	
ra se	k->7	n->2	
ra si	d->19	f->1	g->23	n->22	t->9	
ra sj	ä->2	
ra sk	a->7	i->5	o->1	r->3	u->3	y->1	ä->2	
ra sl	u->7	å->1	
ra sm	å->4	
ra sn	a->4	ä->1	
ra so	c->3	l->1	m->14	
ra sp	e->3	
ra st	a->8	e->1	o->11	r->6	u->2	ä->2	å->2	ö->7	
ra su	b->2	m->3	
ra sv	å->5	
ra sy	f->1	m->1	n->4	s->8	
ra sä	g->4	k->7	m->1	r->5	t->10	
ra så	 ->18	.->2	d->7	
ra ta	 ->1	c->3	l->2	n->4	
ra te	k->1	x->2	
ra ti	d->3	l->72	m->2	
ra tj	ä->4	
ra to	m->1	r->1	x->1	
ra tr	a->5	e->4	o->1	u->2	ä->1	
ra tu	r->1	
ra tv	i->1	å->11	
ra ty	d->2	n->1	
ra un	d->13	g->2	i->8	
ra up	p->17	
ra ur	 ->2	s->1	
ra ut	 ->2	.->2	a->2	b->3	e->1	f->2	g->1	i->1	m->2	r->2	t->2	v->6	
ra va	c->1	d->11	k->2	l->1	p->1	r->9	
ra ve	c->15	r->2	
ra vi	d->3	k->8	l->18	n->3	s->5	t->1	
ra vo	r->1	
ra vä	d->2	g->2	l->10	r->8	s->2	x->1	
ra vå	r->8	
ra yt	l->1	t->6	
ra Ös	t->3	
ra äg	d->1	n->1	
ra än	d->20	n->2	
ra är	 ->28	l->2	
ra å 	m->1	
ra år	 ->10	.->3	e->19	s->1	
ra åt	 ->1	a->2	e->2	g->14	
ra ög	o->3	
ra ök	a->1	
ra ön	s->1	
ra öp	p->1	
ra ör	o->1	
ra ös	t->2	
ra öv	e->19	
ra! D	e->1	
ra!Mä	n->1	
ra"..	 ->1	
ra".D	e->1	
ra, 1	6->1	
ra, a	d->1	n->2	t->6	
ra, b	o->1	
ra, d	e->5	
ra, e	f->1	
ra, f	ö->5	
ra, g	e->1	ö->1	
ra, h	a->2	e->1	j->1	
ra, i	 ->3	b->1	n->2	
ra, k	o->2	
ra, m	e->7	å->1	
ra, o	c->8	m->1	
ra, p	å->1	
ra, s	o->2	ä->1	å->2	
ra, u	n->1	p->1	t->2	
ra, v	a->2	i->3	
ra, ä	r->3	v->1	
ra, å	t->1	
ra. M	e->1	
ra.Al	l->1	
ra.Av	 ->1	
ra.Ba	k->1	
ra.De	s->1	t->12	
ra.Dä	r->3	
ra.EG	-->1	
ra.En	 ->3	l->2	
ra.Fö	r->2	
ra.He	r->2	
ra.Hä	r->1	
ra.I 	f->1	v->1	
ra.In	o->1	
ra.Ja	g->15	
ra.Lä	g->1	
ra.Lå	t->2	
ra.Me	d->1	n->2	
ra.Mi	n->1	
ra.Må	n->1	
ra.Na	t->1	
ra.Nu	 ->1	
ra.Nä	r->2	
ra.Oc	h->1	
ra.Pa	r->1	
ra.Pe	r->1	
ra.På	 ->2	
ra.So	m->1	
ra.Sä	g->1	
ra.Un	g->1	
ra.Va	d->1	
ra.Vi	 ->4	
ra: I	 ->1	
ra: V	a->1	
ra: g	e->1	
ra: r	ä->1	
ra: s	k->1	
ra: u	t->1	
ra: Ä	v->1	
ra; f	ö->2	
ra?An	s->1	
ra?De	t->1	
ra?Ja	g->1	
rabba	 ->1	d->27	r->3	s->7	t->12	
rabeh	a->5	
rabis	k->6	
rabla	"->1	
rabre	p->1	
rabst	a->2	
rabvä	r->1	
raca 	M->3	
racka	t->1	
raco-	a->1	
rad A	d->1	
rad a	n->2	r->1	t->2	v->9	
rad b	e->3	l->1	o->1	y->1	
rad d	e->1	o->2	
rad e	f->1	l->2	n->3	
rad f	o->2	r->3	ö->5	
rad g	e->1	r->1	
rad i	 ->7	m->1	n->6	
rad k	o->5	r->1	v->1	
rad m	a->6	e->1	i->1	
rad n	a->1	
rad o	c->3	l->2	
rad p	o->2	r->1	u->1	å->4	
rad r	e->1	ä->1	
rad s	a->2	e->1	i->2	k->1	m->1	o->3	y->1	
rad t	a->1	i->5	
rad u	n->1	t->1	
rad v	e->3	i->1	
rad y	r->1	
rad ä	n->1	r->1	
rad ö	v->9	
rad, 	i->1	s->1	t->1	
rad.D	e->1	
rad.H	e->1	
rad.K	o->1	
rad.M	e->2	å->1	
rad.U	t->1	
rad.V	e->1	
rade 	-->1	1->1	E->2	a->14	b->8	d->12	e->3	f->20	g->4	h->5	i->17	j->1	k->19	l->5	m->14	n->3	o->16	p->13	r->7	s->16	t->7	u->2	v->5	y->1	å->4	ö->1	
rade,	 ->6	
rade.	 ->1	A->1	D->3	F->2	H->1	M->1	S->1	V->1	
raden	 ->2	.->1	
rader	 ->4	.->2	;->1	a->3	n->2	
rades	 ->24	,->1	.->1	
radet	 ->2	.->1	
radik	a->16	
radio	l->2	
radit	i->19	
radox	,->1	a->5	
radvi	s->3	
rael 	a->4	b->1	d->1	f->2	h->1	i->1	m->1	o->10	v->1	
rael,	 ->4	
rael-	S->1	
rael.	D->2	S->1	
rael?	E->1	
raele	r->5	
raeli	s->15	
raelk	r->1	
raels	 ->6	
raf o	m->1	
rafat	s->1	
raff 	o->2	
raff,	 ->1	
raff-	 ->2	
raffa	 ->1	s->3	
raffb	e->1	
raffl	a->1	
raffp	r->2	
raffr	ä->28	
rafi 	p->1	
rafi.	D->1	V->1	
rafik	 ->2	-->1	.->2	e->3	l->1	
rafin	.->1	
rafis	k->10	
rafry	t->2	
raft 	2->1	a->3	b->1	d->3	e->1	f->4	h->1	i->3	k->1	m->1	n->2	o->3	p->2	s->7	t->2	u->1	v->2	
raft,	 ->9	
raft.	D->2	H->1	M->1	V->1	
raft?	 ->1	N->1	
rafte	n->17	r->9	
raftf	u->12	
rafti	g->34	
rafts	a->4	o->1	p->2	r->1	s->1	v->1	
raftt	a->1	r->4	
raftv	e->8	
rag -	 ->1	
rag a	t->5	v->1	
rag d	e->2	
rag e	f->1	
rag f	r->5	ö->1	
rag h	a->1	
rag i	 ->3	n->3	
rag k	o->2	
rag m	e->1	
rag o	c->1	m->2	
rag s	k->2	o->10	
rag t	i->14	
rag v	a->1	
rag ä	n->1	r->2	
rag å	t->2	
rag, 	h->1	i->1	
rag.B	e->1	
rag.D	e->1	
rag.H	e->1	
rag.R	e->1	
rag.V	i->2	
rag: 	j->1	
raga.	V->1	
ragan	d->114	
raged	i->4	
ragel	s->1	
ragen	 ->17	,->3	.->6	:->1	s->2	
raget	 ->67	)->4	,->14	.->20	;->1	?->1	s->14	
ragis	k->6	
ragit	 ->12	
ragma	t->1	
ragna	 ->1	
ragni	n->48	
ragra	f->3	
ragsa	n->1	r->1	
ragsf	ä->1	
ragsg	i->8	
ragsm	ä->1	
ragsn	a->1	
ragsr	e->2	
ragss	i->1	
ragst	e->2	
ragsä	n->3	
rahan	d->1	
rahus	 ->1	
raine	 ->1	,->1	
rak h	a->2	
rak i	n->1	
rak k	u->1	
rak l	o->1	
rak m	e->1	
rak s	e->1	o->1	
rak v	a->1	
rak ö	v->1	
rak, 	s->1	
rak.D	e->2	
rak.T	r->1	
rak?N	e->1	
raka 	m->2	
rakam	m->1	
rakas	s->1	
rakel	 ->1	
raket	 ->2	
rakis	k->1	
rakop	o->5	
rakry	g->1	
raks 	b->1	p->1	s->1	
rakt 	b->1	f->1	m->1	o->1	u->1	
rakt.	V->1	
rakt:	 ->1	
rakta	 ->6	n->2	r->18	s->8	t->1	
rakte	r->2	t->1	
raktf	a->1	
rakti	g->4	k->10	s->23	v->2	
raktä	r->9	
ral I	n->2	
ral b	e->1	
ral d	e->1	
ral f	r->1	
ral p	l->1	r->1	
ral r	o->2	
ral s	o->1	t->2	
ral å	k->1	
ral, 	d->1	
ral- 	o->6	
ral.F	ö->1	
ral.H	u->1	
rala 	a->1	b->4	d->1	e->1	f->2	g->4	i->3	k->2	l->2	m->1	o->3	p->9	s->1	u->1	v->1	
rala,	 ->2	
ralas	i->6	
ralat	l->1	
ralba	n->8	
ralde	m->1	
raldi	r->17	
ralen	 ->1	?->1	
raler	 ->2	.->1	
raleu	r->1	
ralfö	r->1	
ralib	e->1	
ralis	e->23	k->5	m->5	t->10	
ralle	l->5	
rallt	 ->8	.->2	
ralse	k->2	
ralt 	E->1	i->1	o->2	p->2	s->2	v->1	ä->1	
ralt,	 ->1	
ram "	K->1	
ram -	 ->4	
ram 8	0->1	
ram D	e->1	
ram a	l->1	v->5	
ram b	e->2	l->1	
ram d	e->19	
ram e	f->1	m->17	n->15	t->23	
ram f	l->1	ö->40	
ram g	e->1	ö->1	
ram h	a->4	ä->4	
ram i	 ->13	n->2	
ram k	a->1	o->2	v->1	
ram l	a->1	ä->1	ö->1	
ram m	e->7	o->1	y->1	å->4	
ram n	i->1	o->1	u->1	ä->1	å->2	
ram o	c->7	m->3	
ram p	r->1	å->5	
ram r	e->4	i->1	
ram s	a->1	i->3	k->3	l->1	o->11	p->1	t->2	y->2	å->2	
ram t	a->1	i->44	r->2	
ram u	n->1	t->1	
ram v	a->2	i->3	å->2	
ram ä	n->2	r->1	v->1	
ram å	s->1	
ram ö	v->2	
ram, 	K->1	a->1	b->1	d->3	f->2	i->1	j->1	m->2	o->5	p->1	r->1	s->6	u->2	v->1	
ram..	(->1	
ram.D	e->5	
ram.F	r->3	ö->1	
ram.G	e->1	ö->1	
ram.H	e->1	u->1	
ram.J	a->2	
ram.K	o->1	u->1	
ram.M	e->2	
ram.N	a->1	
ram.O	m->1	
ram.R	e->1	
ram.S	l->1	t->1	y->1	
ram.T	i->1	
ram.V	i->2	
ram?J	a->1	
ram?V	i->1	
raman	s->1	
ramar	 ->2	,->3	.->1	n->2	
ramat	i->6	
ramav	t->3	
ramen	 ->57	,->3	
ramet	e->1	r->1	
ramfa	r->1	
ramfö	r->145	
ramgi	c->1	
ramgå	 ->1	n->38	r->12	t->1	
ramhä	r->1	v->4	
ramhå	l->17	
ramhö	l->2	
ramid	i->1	
ramka	s->1	
ramko	m->10	
ramla	d->1	g->12	
ramlä	g->8	
ramme	 ->1	n->35	t->73	
ramni	n->2	
ramp 	J->1	i->1	
rampe	r->3	
rampl	a->8	
rampr	o->12	
ramru	n->1	
ramsk	j->1	r->1	
ramst	e->32	ä->10	å->5	ö->1	
ramt 	f->1	
ramta	g->5	
ramti	d->107	
ramtr	ä->2	
ramtv	i->2	
ramut	f->1	
ramve	r->1	
ramvi	l->3	
ramåt	 ->12	,->3	.->7	
ramöv	e->2	
ran H	a->1	
ran a	n->1	t->9	
ran f	r->3	ö->2	
ran g	j->1	
ran h	a->1	
ran i	 ->1	
ran j	a->1	
ran m	e->1	
ran o	c->2	f->1	m->5	
ran s	k->1	o->1	
ran t	i->3	
ran u	n->1	
ran v	a->1	
ran ö	v->1	
ran, 	s->2	t->1	u->1	
ran- 	o->1	
ran.)	 ->1	
ran.D	e->2	
ran.F	r->1	
ran.N	i->1	ä->1	
ran?F	r->1	
ran?O	m->1	
ranat	i->1	
ranbi	l->8	
ranc,	 ->1	
ranca	s->1	
rance	,->1	.->1	
ranci	s->1	
rand 	b->1	f->1	i->1	s->1	
rand.	J->1	
randa	 ->1	,->1	
rande	 ->429	!->6	,->37	.->19	:->1	?->1	b->2	f->1	k->9	l->3	n->61	r->3	s->114	t->91	
randi	g->2	
randm	ä->1	
rando	m->14	
randr	a->10	
rands	 ->1	
range	m->4	r->2	
ranin	v->1	
raniu	m->2	
rankr	a->4	i->39	
ranle	d->2	
ranna	 ->2	n->1	r->2	
rannh	e->1	
rannl	a->1	ä->1	
ranns	a->1	k->1	
ranoi	s->1	
rans 	g->1	m->1	o->2	
rans,	 ->3	
rans.	D->2	E->1	
ransc	h->7	
ranse	n->1	u->1	
ransi	t->7	
ransk	 ->2	a->62	n->23	t->2	u->1	
ransl	a->1	u->1	
ransm	ä->5	
ransp	o->108	
ransv	a->6	
rant 	f->2	h->2	i->1	p->1	s->2	t->1	ö->1	
rant.	D->1	S->1	
rante	r->59	
ranti	 ->9	,->1	.->1	e->15	f->2	n->3	s->3	
rantö	r->3	
ranva	p->4	
ranvä	n->18	
ranz 	F->3	
ranço	i->1	
raord	i->1	
raper	i->1	
rappo	r->109	
rapro	d->1	
rar -	 ->1	
rar 1	5->1	
rar 3	-->1	
rar E	u->3	
rar I	n->1	
rar P	r->1	
rar R	h->1	
rar S	e->1	
rar a	l->7	n->1	r->1	t->30	v->3	
rar b	a->2	e->1	u->1	ä->1	
rar d	e->66	i->1	o->1	ä->1	å->1	
rar e	l->1	n->10	r->5	t->7	x->2	
rar f	a->3	ö->17	
rar g	e->1	r->1	
rar h	a->1	e->5	o->3	u->1	ä->6	
rar i	 ->21	.->1	n->20	
rar j	a->14	u->1	
rar k	l->1	o->6	r->3	v->1	
rar l	ä->1	ö->1	
rar m	a->7	e->7	i->7	o->4	y->1	ä->1	
rar n	a->1	e->1	i->2	u->1	y->4	ä->1	å->2	
rar o	c->13	l->1	m->4	s->6	
rar p	a->5	e->3	r->2	å->7	
rar r	e->1	å->3	
rar s	a->2	i->12	k->1	o->5	u->1	v->1	ä->2	
rar t	e->1	i->25	j->1	y->1	
rar u	n->1	p->1	t->3	
rar v	a->2	e->1	i->11	ä->1	å->5	
rar y	t->1	
rar ä	l->1	n->1	r->1	v->3	
rar å	t->1	
rar ö	p->1	v->3	
rar! 	A->1	B->1	D->2	E->1	F->2	H->1	J->4	N->1	P->1	S->2	T->1	V->1	
rar!J	a->1	
rar!M	i->1	
rar!T	i->1	
rar, 	W->1	a->1	d->1	f->1	h->1	i->1	j->3	k->7	m->1	o->4	p->2	s->3	t->1	u->1	v->1	ä->2	
rar..	.->1	
rar.A	m->1	
rar.D	e->1	
rar.F	ö->3	
rar.H	ä->1	
rar.J	a->1	
rar.N	a->1	
rar.R	ä->1	
rar.S	k->1	
rar.V	i->2	
rar: 	D->1	
rar; 	m->1	
rara 	l->1	
rarbe	t->2	
rare 	a->3	b->2	d->1	e->1	f->2	h->1	i->4	n->1	o->6	p->2	s->4	t->4	ä->6	ö->1	
rare,	 ->4	
rare.	D->1	I->1	V->1	
raren	 ->1	
rares	 ->1	
rarki	.->1	n->2	s->1	
rarlä	k->1	
rarna	 ->9	,->4	s->4	
rars 	u->1	
rart,	 ->1	
rarte	r->1	
rartr	a->1	
rarv 	o->1	
rarv,	 ->2	
rarv.	E->1	
rarve	t->1	
ras 4	0->1	
ras E	u->1	
ras a	n->11	r->1	t->6	u->1	v->28	
ras b	e->2	l->1	r->1	ä->1	ö->1	
ras c	e->2	
ras d	a->1	e->4	i->2	ö->1	
ras e	f->1	g->2	k->3	l->3	n->2	v->1	x->2	
ras f	a->2	l->1	o->1	r->4	u->2	ö->22	
ras g	e->8	
ras h	a->1	j->1	u->2	y->1	
ras i	 ->30	n->9	
ras j	u->2	
ras k	a->1	o->6	
ras l	a->1	e->2	i->2	
ras m	e->16	i->1	o->1	ö->1	
ras n	a->3	u->1	ä->4	å->1	
ras o	b->1	c->14	f->2	l->2	m->3	r->2	v->1	
ras p	r->1	å->13	
ras r	a->2	e->1	i->1	u->1	ä->4	
ras s	a->3	e->2	k->2	n->3	o->7	t->5	v->1	ä->3	å->4	
ras t	a->1	i->12	r->1	v->1	
ras u	n->5	p->4	t->3	
ras v	a->1	e->1	i->3	ä->2	
ras y	t->1	
ras ä	n->1	r->1	v->1	
ras å	r->1	t->2	
ras ö	d->1	n->1	v->3	
ras!D	e->1	
ras!G	e->1	
ras, 	M->1	e->3	f->1	g->1	i->1	k->1	o->5	s->5	u->4	v->1	
ras. 	D->1	M->1	
ras.A	t->1	
ras.B	e->1	
ras.D	e->10	
ras.E	k->1	t->1	
ras.F	r->3	ö->1	
ras.G	e->1	r->1	
ras.I	 ->4	
ras.J	a->3	
ras.M	a->1	e->2	
ras.N	i->1	
ras.P	a->1	r->1	
ras.S	a->1	l->1	n->1	
ras.U	n->1	
ras.V	i->7	å->1	
ras.Y	t->1	
ras; 	e->1	
rasad	e->2	
rasas	 ->1	
rasat	 ->1	
rasbo	u->5	
rasch	e->3	
raser	,->1	
rasha	t->1	
rasil	i->1	
rasis	m->14	t->12	
raska	d->1	
rasma	t->1	
rassl	a->1	
rasso	n->1	
rasst	 ->1	
rast 	a->1	e->1	f->2	h->1	k->1	m->1	p->1	u->1	v->1	å->2	
rast.	V->1	
raste	 ->5	n->1	r->1	
rasti	s->3	
rastr	u->15	
rat -	 ->2	,->1	
rat A	d->1	
rat E	r->1	u->1	
rat F	l->1	
rat S	j->1	
rat a	l->1	t->8	v->1	
rat b	e->3	i->1	r->1	
rat d	e->12	i->1	o->1	
rat e	n->5	r->2	t->2	
rat f	l->1	r->2	ö->7	
rat g	e->1	
rat h	i->1	o->1	u->2	å->1	ö->1	
rat i	 ->6	n->2	
rat k	l->1	o->4	
rat l	i->2	
rat m	e->2	i->2	y->1	å->1	
rat n	u->1	å->2	
rat o	c->3	m->4	s->2	
rat p	r->2	å->1	
rat r	ä->1	
rat s	e->1	i->9	o->3	y->1	ä->1	
rat t	i->2	r->1	ä->1	
rat v	a->1	i->1	ä->1	å->3	
rat å	t->1	
rat, 	a->1	b->1	e->2	f->1	i->1	n->1	o->4	p->1	v->1	ä->1	
rat. 	H->1	
rat..	H->1	
rat.B	i->1	
rat.D	e->3	
rat.E	n->1	
rat.H	e->1	
rat.J	a->3	
rat.K	u->1	
rat.T	i->1	
rat.V	a->1	
rat; 	a->1	
rata 	f->1	o->2	
ratal	 ->1	s->5	
ratar	 ->1	
rateg	i->63	
raten	 ->1	.->1	
rater	 ->12	)->2	.->1	n->9	
rates	-->1	
ratet	 ->11	,->1	
rati 	d->1	i->1	k->1	o->9	s->1	u->1	
rati"	 ->1	
rati,	 ->3	
rati.	D->2	E->2	F->1	H->1	I->1	K->1	M->1	
ratie	r->3	
ratif	i->13	r->1	
ratin	 ->11	,->1	.->4	o->4	s->4	
ratio	n->69	
ratir	e->1	
ratis	 ->4	k->91	
rativ	 ->2	a->17	t->5	
ratog	e->2	
ratom	 ->3	)->1	
rator	i->3	
rats 	-->2	a->5	e->1	f->3	g->1	h->2	i->7	m->2	o->3	p->2	t->3	v->2	
rats,	 ->6	
rats.	D->3	H->1	M->1	
rats?	F->1	
ratta	s->1	
rattr	e->1	
ratul	a->6	e->31	
ratur	 ->2	,->1	e->8	f->2	
ratus	e->3	
ratör	e->2	
rauma	t->1	
rav -	 ->1	
rav 4	0->1	
rav 8	 ->1	
rav b	e->1	
rav d	e->2	
rav e	t->1	
rav f	r->3	ö->2	
rav g	ö->1	
rav i	 ->1	
rav l	e->1	
rav n	ä->1	
rav o	c->2	m->1	
rav p	å->17	
rav s	k->2	o->7	
rav t	i->1	
rav u	p->1	
rav v	i->1	
rav, 	d->1	e->1	f->1	m->1	
rav.(	S->1	
rav..	 ->1	
rav.D	e->2	
rav.E	r->1	
rav.R	å->1	
rav?V	i->1	
rava 	g->1	
raval	l->1	
ravar	 ->1	
raven	 ->23	.->3	:->1	
raver	a->4	y->1	
ravet	 ->13	.->3	
ravt 	s->1	
rax a	v->1	
rax e	f->1	
rax i	n->1	
raxis	 ->5	.->2	e->1	
ray, 	h->1	
raça 	M->5	
rb, e	n->1	
rba-,	 ->1	
rbala	 ->1	
rban"	 ->1	
rband	 ->2	
rbani	s->1	
rbar 	k->2	m->1	
rbar.	D->1	
rbara	 ->6	,->1	.->1	
rbarh	e->1	
rbari	e->1	s->1	
rbarm	a->1	
rbart	 ->2	,->1	.->1	
rbast	i->1	
rbaye	r->1	
rbedö	m->1	
rbegr	i->1	
rbehå	l->6	
rbela	s->3	
rbema	n->1	
rber 	o->2	
rber,	 ->3	
rbera	d->1	
rbere	d->25	t->2	
rbern	a->2	
rbest	ä->2	
rbeta	 ->64	,->1	.->3	?->1	d->2	l->1	n->11	r->35	s->2	t->14	
rbete	 ->112	,->11	.->28	?->3	n->9	t->51	
rbets	-->2	a->5	b->6	d->4	f->2	g->13	i->2	k->6	l->46	m->15	n->3	o->11	p->14	r->4	t->83	v->5	
rbett	 ->1	
rbetä	n->6	
rbi d	e->1	
rbifa	r->2	
rbigå	 ->1	e->4	s->1	
rbiha	n->1	
rbild	a->1	
rbind	a->1	e->21	
rbise	e->1	
rbisk	 ->1	a->5	
rbjud	a->19	e->13	i->1	
rbjöd	s->1	
rblev	 ->1	
rbli 	-->1	b->1	e->3	l->1	s->1	v->1	
rblic	k->1	
rblir	 ->6	
rblås	e->2	
rbrin	g->1	
rbrit	a->14	
rbrot	t->1	
rbruk	n->1	
rbryg	g->3	
rbryt	e->2	
rbrän	n->2	
rbud 	f->1	m->9	o->1	
rbud,	 ->2	
rbud.	D->2	V->1	
rbude	t->8	
rbuds	f->1	p->1	
rbund	e->1	i->3	s->8	
rbätt	r->78	
rböld	 ->1	
rböra	n->1	
rbörl	i->10	
rce b	ö->1	
rcelo	n->2	
rcent	r->1	
rcour	s->1	
rcykl	a->4	
rd - 	a->1	
rd 2 	i->1	
rd Co	r->1	
rd In	g->2	
rd Ko	u->1	
rd an	s->1	
rd ar	b->1	
rd at	t->4	
rd av	 ->3	s->2	
rd bl	a->1	
rd br	ä->1	
rd de	l->1	
rd dä	r->1	
rd ef	t->1	
rd ek	o->1	
rd el	l->1	
rd en	 ->1	
rd eu	r->1	
rd fr	å->1	
rd fö	r->9	
rd gr	a->1	
rd i 	F->1	S->1	d->1	h->1	
rd in	g->1	t->1	
rd iv	e->1	
rd ja	g->1	
rd ka	m->1	t->1	
rd ko	m->2	
rd kr	a->1	
rd ku	l->1	
rd ma	k->1	
rd me	d->2	
rd mi	l->1	n->1	
rd nä	r->1	
rd oc	h->16	
rd om	 ->3	
rd pr	ö->1	
rd på	 ->1	
rd si	t->1	
rd sj	u->1	
rd sk	a->1	
rd so	m->9	
rd ta	 ->1	
rd te	r->1	
rd ti	d->1	l->2	
rd ur	v->1	
rd va	d->1	r->1	
rd vi	 ->3	l->1	
rd), 	r->1	
rd, b	l->1	
rd, d	ä->1	å->1	
rd, h	y->1	
rd, m	e->2	
rd, o	c->5	
rd, s	a->1	o->2	å->1	
rd, t	i->1	r->1	
rd, ä	r->1	
rd-af	f->1	
rd-fö	r->1	
rd.Be	d->1	
rd.De	 ->1	s->1	t->3	
rd.Dä	r->1	
rd.Eu	r->1	
rd.He	r->1	
rd.I 	s->1	
rd.Ja	g->1	
rd.Un	d->1	
rd.Vi	 ->2	
rd: "	D->1	O->1	
rd; d	e->1	
rd; i	n->2	
rda a	k->1	r->3	t->1	v->1	
rda d	e->2	
rda e	f->1	l->2	n->1	u->1	
rda f	o->1	r->1	ö->1	
rda g	a->1	
rda h	i->1	ä->1	
rda k	a->1	o->5	r->1	u->1	
rda l	a->1	ä->1	
rda m	e->3	
rda n	y->1	ä->1	ö->1	
rda o	c->2	
rda p	a->1	e->3	o->3	
rda r	e->3	å->1	
rda s	k->1	m->1	o->2	t->1	u->1	y->1	
rda t	r->1	å->1	
rda u	t->2	
rda v	e->1	i->1	ä->1	å->1	
rda ä	r->1	
rda, 	f->1	i->1	n->1	r->1	s->1	
rda.D	e->1	
rda.H	a->1	e->1	
rda.O	c->1	
rda?D	e->1	
rdad.	S->1	
rdade	 ->1	s->1	
rdag 	k->1	
rdag,	 ->1	
rdage	n->3	
rdagl	i->2	
rdala	g->4	
rdaly	d->2	
rdam 	-->1	1->1	i->1	o->1	p->1	s->1	t->1	v->1	ä->1	
rdam,	 ->3	
rdam.	N->1	
rdame	r->4	
rdamf	ö->27	
rdamr	e->1	
rdan 	a->1	b->1	i->1	m->1	s->1	
rdan.	A->1	D->1	J->1	
rdand	e->7	
rdani	e->1	
rdans	 ->1	
rdar 	d->2	m->1	r->1	s->1	
rdar,	 ->1	
rdare	 ->3	.->1	
rdas 	n->1	
rdas.	H->1	
rdast	 ->1	.->1	
rdat 	a->1	f->1	n->1	
rdats	 ->1	
rdbru	k->56	
rdbrä	n->1	
rdbäv	n->10	
rde K	o->1	
rde a	n->1	t->2	v->1	
rde b	e->1	l->3	ö->1	
rde d	e->10	o->1	å->1	
rde e	f->1	g->1	n->4	t->2	
rde f	i->1	r->1	å->2	ö->3	
rde g	e->2	ö->1	
rde h	a->8	y->1	
rde i	 ->8	n->6	
rde j	a->1	u->2	
rde k	a->2	l->1	o->4	u->2	
rde m	a->2	e->2	i->2	å->1	
rde n	ä->2	å->1	
rde o	c->2	s->1	
rde p	a->1	e->1	l->1	o->1	u->1	å->2	
rde r	e->5	i->1	ä->1	å->1	
rde s	e->1	k->4	o->2	t->2	
rde t	a->1	i->3	ä->1	
rde u	n->1	p->1	t->4	
rde v	a->10	i->4	
rde, 	a->1	n->1	t->1	
rde- 	o->1	
rde-l	ä->1	
rde.D	e->2	
rde.G	e->1	
rde.J	a->2	
rde.L	å->1	
rde.N	ä->1	
rde.T	a->1	
rdeau	x->1	
rdede	l->2	
rdefu	l->7	
rdege	m->3	
rdel 	f->1	m->2	
rdel,	 ->2	
rdel.	M->2	
rdela	 ->2	d->1	k->2	r->5	s->3	t->2	
rdele	n->1	
rdeln	i->23	
rdelö	s->1	
rdemo	n->1	
rden 	"->1	a->3	d->1	h->1	i->3	m->1	o->2	p->3	s->6	t->2	
rden,	 ->3	
rden.	D->2	H->1	J->1	R->1	
rdena	 ->3	.->1	
rdenn	e->1	
rdens	 ->3	
rdent	l->25	
rder 	-->1	U->1	a->5	b->4	d->3	e->10	f->32	g->3	h->3	i->11	k->4	m->10	n->3	o->8	p->6	s->49	t->6	u->1	v->4	ä->3	
rder,	 ->13	
rder.	A->1	D->7	E->1	F->4	I->1	J->2	M->1	T->1	U->1	V->1	Ä->1	
rder?	.->1	
rdera	 ->10	d->4	r->2	s->4	t->1	
rderi	n->44	
rderl	i->5	
rdern	a->22	
rdes 	a->3	d->2	e->1	f->1	i->2	o->1	t->2	u->1	v->1	
rdes,	 ->1	
rdes.	D->1	
rdess	k->1	t->1	
rdet 	"->1	a->3	e->1	f->3	g->1	i->2	k->1	o->3	t->9	ä->1	
rdet.	H->1	J->1	
rdeur	o->1	
rdför	a->223	
rdhet	 ->1	
rdig 	l->2	m->2	o->2	
rdig.	P->1	
rdiga	 ->5	,->1	n->1	r->3	t->1	
rdigh	e->18	
rdigs	t->1	
rdigt	 ->4	
rdinä	r->1	
rdirl	ä->2	
rdise	r->9	
rdisk	 ->2	a->2	
rdita	l->1	
rdjup	a->6	n->5	
rdkus	t->1	
rdlad	e->1	
rdlig	a->6	t->1	
rdlis	t->1	
rdmån	 ->1	
rdna 	d->1	e->1	f->1	g->1	l->1	u->1	v->1	
rdnac	k->2	
rdnad	 ->6	e->4	
rdnan	d->2	
rdnar	 ->1	e->3	n->1	
rdnas	 ->2	
rdnat	 ->2	s->1	
rdnin	g->155	
rdo R	o->1	
rdom 	a->4	f->1	n->1	
rdom,	 ->1	
rdoma	r->1	
rdoml	i->1	
rdoms	f->1	h->1	
rdon 	(->2	-->1	b->1	e->1	f->1	i->3	k->1	m->1	o->3	p->3	s->13	u->1	ä->1	
rdon,	 ->8	
rdon.	D->3	J->3	L->1	M->1	V->1	
rdon?	V->1	
rdonN	ä->1	
rdone	n->6	t->1	
rdons	i->1	p->1	t->3	ä->1	å->1	
rdor 	s->1	
rdorn	a->1	
rdra 	d->2	e->1	
rdrag	 ->9	.->2	e->141	s->12	
rdran	 ->5	,->1	.->1	
rdrar	 ->2	
rdras	 ->4	.->1	
rdrat	 ->1	
rdre 	p->1	
rdrif	t->3	
rdrik	t->2	
rdrin	g->1	
rdriv	a->1	e->11	n->1	
rdröj	a->1	
rds r	e->1	
rds- 	o->1	
rdsbu	s->1	
rdska	l->1	
rdsli	s->1	
rdslö	s->2	
rdsmy	n->1	
rdsmå	l->1	
rdsom	r->1	
rdspa	k->2	
rdspl	a->3	
rdspr	o->1	
rdspu	n->1	
rdssk	i->1	
rdsst	a->2	
rdsto	w->3	
rdsut	v->1	
rdsvi	n->1	
rdtid	.->1	
rdtys	k->1	
rdubb	l->2	
rdunk	l->1	
rdvrä	n->1	
rdvän	d->1	
rdväs	t->1	
rdärv	a->2	b->1	l->1	
rdöma	 ->7	n->6	
rdöme	r->5	
rdömt	 ->2	
rdörr	e->1	
re - 	,->1	j->1	n->1	o->1	u->1	
re 11	5->1	
re 15	 ->1	
re 20	0->1	
re 21	 ->1	
re 35	 ->1	
re 4,	 ->1	
re Am	s->1	
re BN	P->1	
re De	 ->1	
re Di	r->1	
re Eu	r->2	
re Hi	t->1	
re Ki	n->1	
re ad	 ->1	
re ak	t->1	
re al	l->3	t->1	
re am	b->1	
re an	 ->1	a->1	d->1	g->2	l->2	s->9	t->1	
re ar	b->1	
re at	t->28	
re av	 ->8	f->1	g->1	r->1	
re ba	l->1	s->1	
re be	d->1	f->3	g->2	h->1	k->1	r->1	s->11	t->6	v->1	
re bi	f->1	l->2	
re bl	i->4	
re bo	r->1	
re br	a->1	
re by	r->4	
re bä	t->1	
re bå	t->1	
re bö	r->2	
re ch	e->1	
re da	g->2	
re de	 ->2	b->2	l->4	m->1	n->5	t->6	
re di	s->3	
re do	m->1	
re du	s->1	
re dy	k->1	
re dä	r->1	
re då	 ->1	
re ef	f->1	t->1	
re ek	o->3	
re el	-->1	l->6	
re em	o->1	
re en	 ->9	e->1	g->1	h->1	l->1	
re et	t->6	
re eu	r->4	
re ex	a->1	e->1	
re fa	l->2	n->3	r->1	t->1	
re fe	m->1	
re fi	n->4	
re fj	ä->1	
re fl	e->1	
re fo	r->2	
re fr	a->6	i->2	å->29	
re fu	n->1	
re fy	r->2	
re få	 ->2	r->2	
re fö	r->67	
re ge	m->1	n->5	
re gj	o->1	
re go	d->2	
re gr	a->4	u->1	ä->3	
re gå	 ->1	n->2	
re gö	r->1	
re ha	d->1	f->2	n->1	r->20	
re he	l->2	
re hi	n->1	t->1	
re ho	s->1	
re hu	r->2	
re hä	n->1	
re hå	l->1	
re hö	r->2	
re i 	D->1	E->3	K->2	T->1	a->2	b->1	d->13	e->2	m->3	p->1	s->1	t->1	u->2	v->3	å->4	
re id	é->1	
re in	f->3	n->2	o->2	r->1	s->3	t->5	v->1	
re it	a->1	
re jo	r->1	
re jä	m->2	
re ka	m->1	n->15	t->2	
re kl	a->1	
re ko	l->4	m->15	n->9	r->1	
re kr	e->1	i->1	ä->3	
re ku	n->5	
re kv	i->1	
re kä	n->2	
re la	g->2	s->1	
re le	g->1	
re li	k->1	
re lä	m->2	n->2	r->1	
re lö	s->1	
re ma	k->2	r->69	
re me	d->12	k->1	l->1	n->1	r->3	s->1	
re mi	g->1	l->3	n->2	
re mo	t->4	
re my	c->2	n->1	
re må	n->11	s->5	
re mö	j->2	
re ni	o->1	v->3	
re nu	 ->1	
re nä	m->3	r->3	s->3	
re nå	g->4	
re oc	h->45	k->3	
re ol	y->1	ä->1	
re om	 ->8	r->7	ö->1	
re or	d->2	o->2	ä->1	
re os	s->1	
re ov	a->1	e->1	
re pa	r->2	
re pe	k->1	n->1	r->4	
re pl	a->2	
re po	l->2	
re pr	e->4	i->2	o->4	
re pu	b->1	n->1	
re på	 ->18	
re re	f->1	g->4	k->1	s->6	
re ri	k->1	s->1	
re ro	l->2	t->1	
re rä	c->1	k->1	t->2	
re sa	d->1	g->1	k->1	m->5	n->1	
re se	 ->1	d->2	n->1	r->2	
re si	g->13	k->1	t->2	
re sj	ä->1	
re sk	a->10	e->1	u->3	y->1	å->2	
re sl	u->1	
re sm	å->1	
re sn	a->1	
re so	c->1	m->37	
re sp	r->1	å->1	
re st	a->4	e->1	o->3	r->3	ä->1	å->3	ö->1	
re su	m->1	
re sy	f->1	s->3	
re sä	k->4	t->8	
re så	 ->2	
re ta	 ->1	k->1	l->6	
re ti	d->7	l->20	o->2	
re tj	ä->4	
re to	l->3	
re tr	o->1	
re tv	ä->2	å->1	
re ty	c->1	d->1	n->1	
re un	d->2	
re up	p->8	
re ut	 ->1	a->1	b->2	g->4	n->1	r->2	s->5	v->7	
re va	c->1	d->2	l->2	r->5	t->8	
re ve	c->3	l->1	t->1	
re vi	 ->1	d->1	k->6	l->4	n->1	r->1	
re vo	l->1	
re vä	s->2	
re än	 ->44	d->3	t->1	
re är	 ->10	
re år	 ->1	.->3	e->2	
re åt	e->2	g->1	
re ök	a->1	n->1	
re ön	s->2	
re öp	p->6	
re öv	e->1	
re!Sk	a->1	
re" s	k->1	o->1	
re", 	o->1	
re, A	l->1	
re, D	a->1	
re, F	ö->1	
re, H	a->1	
re, a	r->1	t->2	
re, b	e->1	r->1	ä->1	å->2	
re, d	e->2	
re, e	n->1	t->1	
re, f	i->1	ö->2	
re, h	a->3	e->2	
re, i	 ->3	n->2	
re, j	a->1	
re, k	a->1	o->1	
re, m	e->8	u->1	y->1	
re, n	ä->3	
re, o	a->1	c->8	s->2	
re, p	r->3	å->2	
re, s	a->1	k->1	o->7	ä->1	å->1	
re, u	n->1	t->2	
re, v	i->5	ä->1	å->1	
re, ä	r->4	
re, å	t->2	
re-At	l->1	
re. D	e->1	
re. O	m->1	
re. Ä	n->1	
re.Al	l->1	
re.At	t->1	
re.Bå	d->1	
re.De	n->1	r->1	s->2	t->15	
re.Dä	r->2	
re.Då	 ->2	
re.Ef	t->2	
re.En	 ->1	
re.Eu	r->2	
re.Fö	r->3	
re.He	r->1	
re.I 	d->2	o->1	s->1	
re.Im	m->1	
re.Ja	g->8	
re.Ko	m->2	
re.Ma	n->2	
re.Me	d->1	n->3	
re.Mi	n->2	
re.Nu	 ->1	
re.Nä	r->1	
re.Pr	o->1	
re.På	 ->1	
re.Ro	t->1	
re.Rå	d->1	
re.So	m->3	
re.Ti	l->2	
re.Tr	o->1	
re.Ur	 ->1	
re.Va	d->1	
re.Vi	 ->5	
re.Vå	r->1	
re.Än	d->2	
re.Är	 ->1	
re.Äv	e->2	
re: b	e->1	
re: d	e->1	
re?De	t->1	
re?Ka	n->1	
re?Oc	h->1	
re?Vi	 ->1	
rea b	e->1	
rea o	c->3	
reage	r->16	
reakt	i->11	o->10	
real 	p->1	
real,	 ->1	
reali	s->9	t->7	
reami	n->8	
reati	v->2	
reatö	r->1	
rebef	o->2	
rebeh	a->1	
rebil	d->1	
reboa	r->1	
rebrå	s->2	
rebyg	g->23	
recir	k->1	
recis	 ->36	a->1	e->11	t->1	
reck 	ä->1	
recov	e->1	
rectn	e->1	
recyc	l->1	
red b	a->1	
red d	a->1	
red e	x->1	
red i	 ->6	
red l	a->1	
red m	e->1	
red o	c->7	
red v	i->1	
red, 	f->1	
red.D	ä->1	
red.H	e->1	u->1	
red.I	 ->1	
reda 	E->1	a->1	d->1	e->1	h->1	m->1	p->3	s->2	u->3	å->1	
reda,	 ->2	
redak	t->1	
redan	 ->155	d->3	
redar	e->6	n->3	
redas	 ->1	t->1	
redd 	a->16	t->3	u->1	ä->1	
redda	 ->13	
redde	 ->1	,->1	n->2	
redel	s->5	
reden	 ->1	s->1	
reder	 ->8	i->2	
redga	t->1	
redie	n->2	
redit	e->2	
redje	 ->56	,->4	:->1	d->6	l->6	
redli	g->10	
redni	n->8	
redo 	a->3	
redog	j->1	ö->9	
redov	i->4	
redra	 ->3	g->160	r->2	
redro	g->1	
reds 	m->1	s->1	
reds,	 ->1	
reds.	J->1	
redsa	n->1	v->3	
redsb	e->2	
redsf	ö->3	
redsk	a->2	
redsp	a->1	r->22	
redss	a->4	t->24	
redsu	p->1	
reduc	e->4	
redöm	l->2	
ree-f	ö->1	
ree-l	o->1	
ree.D	e->1	
reell	 ->1	.->1	a->2	
refal	l->20	
refer	e->7	
refle	k->7	
refor	m->134	
refte	r->13	
refus	e->1	
reföl	l->1	
regel	 ->3	b->16	m->2	n->6	r->2	s->2	v->19	
reger	a->1	i->281	
regi,	 ->1	
regic	k->1	
regim	e->3	
regio	n->251	
regis	t->20	
regle	r->126	
regri	p->1	
regåe	n->15	
regån	g->2	
rehab	i->1	
rehav	a->1	
reisk	a->1	
rejud	i->4	
rejäl	t->3	
reker	n->1	
rekis	k->6	
rekla	m->2	n->15	
rekom	 ->1	m->65	s->1	
rekon	o->3	s->3	
rekor	d->2	
rekry	t->1	
rekt 	a->5	b->6	d->1	e->3	f->3	g->1	h->1	i->1	k->3	l->1	m->2	n->1	o->3	p->1	s->8	t->8	u->2	
rekt,	 ->2	
rekt.	D->3	F->2	J->1	M->1	U->1	
rekt;	 ->1	
rekta	 ->9	.->1	
rekti	n->1	v->193	
rekto	r->18	
rektö	r->1	
rekve	n->1	
rela 	S->1	
relat	e->4	i->22	
releg	a->1	
relev	a->9	
relig	g->26	i->4	
relik	e->1	
relim	i->3	
rell 	b->3	f->1	l->1	m->2	o->1	r->1	s->1	t->1	v->2	
rella	 ->28	
rellt	 ->14	,->1	
relse	 ->6	,->2	.->3	h->1	n->10	r->6	
reläg	g->2	
rema 	f->1	h->1	
remen	,->1	
remhö	g->14	
remis	m->5	s->1	t->5	
remiä	r->10	
remot	 ->19	
rems-	 ->1	
remsa	n->2	
remt 	h->2	r->1	s->1	
remål	 ->13	
remån	a->1	
ren -	 ->2	
ren 2	0->1	
ren H	a->1	
ren K	a->1	
ren V	i->1	
ren a	n->3	t->6	v->1	
ren b	a->1	e->4	i->1	
ren d	u->1	ä->2	ö->1	
ren e	f->1	l->2	n->4	r->1	v->1	
ren f	a->1	i->2	r->2	å->1	ö->33	
ren g	e->1	j->1	ä->1	
ren h	a->13	e->1	o->1	
ren i	 ->12	f->1	n->5	
ren j	ä->1	
ren k	a->3	r->2	
ren l	o->1	
ren m	e->3	å->3	
ren n	a->1	ä->1	
ren o	c->28	m->7	
ren p	e->1	l->1	å->5	
ren r	e->2	
ren s	a->4	e->3	k->8	o->5	t->2	å->1	
ren t	i->4	ä->1	
ren u	p->1	t->3	
ren v	a->2	i->3	
ren ä	n->1	r->11	
ren å	r->1	
ren ö	v->1	
ren).	H->1	
ren)J	a->1	
ren, 	A->1	T->1	a->2	d->2	e->3	f->5	i->1	m->3	n->1	o->8	p->1	r->1	s->5	t->3	u->1	v->3	
ren.)	.->1	F->3	H->1	
ren..	 ->1	
ren.A	t->1	
ren.D	e->7	ä->1	
ren.E	u->1	
ren.F	ö->1	
ren.H	e->1	u->1	
ren.I	 ->3	
ren.J	a->5	
ren.K	o->1	
ren.M	a->1	e->1	
ren.O	m->2	
ren.R	i->1	
ren.T	i->1	v->1	
ren.V	i->3	
ren.Ö	v->1	
ren; 	e->1	
ren?I	 ->1	
ren?V	i->1	
ren?Ä	r->1	
rena 	a->1	d->3	f->2	g->1	m->1	s->2	v->1	
renad	e->16	
renan	d->5	
renar	 ->7	,->1	.->1	e->4	n->2	
renas	 ->1	
rend 	f->1	i->1	j->1	o->1	u->1	
rend!	 ->2	
rend,	 ->2	
rend-	 ->1	
renda	 ->2	i->1	
rendb	e->1	
rende	 ->4	,->2	.->2	n->8	t->5	
rends	 ->2	
rendt	 ->6	,->1	
rengu	e->2	
rengö	r->3	
renhe	t->24	
renin	g->22	
renkl	a->7	i->1	
renli	g->9	
renov	e->3	
rens 	a->2	b->1	d->1	e->3	f->6	g->2	h->1	i->7	k->3	l->1	m->13	n->1	o->34	p->2	r->3	s->12	t->2	u->2	v->1	ä->5	
rens!	V->1	
rens,	 ->12	
rens-	 ->2	
rens.	D->5	F->1	J->1	M->1	O->1	S->1	
rens/	d->1	
rens:	 ->1	
rens?	E->1	J->1	
rensa	 ->2	r->1	v->1	
rensb	e->9	
rensd	e->2	o->1	u->2	
rense	n->162	r->6	
rensf	r->5	ö->3	
rensh	i->2	ä->2	
rensi	n->2	
rensk	o->18	r->37	u->5	
rensm	e->1	i->1	y->8	å->1	
rensn	a->2	i->7	
renso	m->2	r->1	
rensp	o->76	r->4	
rensr	a->1	e->10	ä->9	
renss	i->1	k->3	t->21	v->1	y->1	
rensu	t->2	
rensv	e->1	i->9	ä->1	
rensä	r->2	
rent 	a->9	f->2	g->1	h->2	i->2	k->2	r->1	t->2	u->1	
renta	 ->28	v->1	
rente	r->1	
renti	e->5	
rents	 ->1	
renz 	b->1	e->1	f->2	o->7	t->1	
renz)	(->1	.->1	
renz,	 ->3	
renzF	r->1	
renzb	e->1	
renör	 ->1	s->2	
rep m	a->1	
repa 	a->1	d->6	m->4	n->2	p->1	v->1	
repa,	 ->1	
repad	e->8	
repar	 ->15	a->2	e->4	
repas	 ->5	.->2	
repat	 ->2	:->1	s->2	
repni	n->1	
repp 	a->1	i->4	o->1	p->3	s->1	
repp,	 ->1	
reppa	 ->1	
reppe	n->1	t->10	
repps	s->2	
repre	n->3	s->21	
repri	s->2	
repub	l->18	
rer -	 ->1	
rer a	t->1	v->4	
rer b	ö->1	
rer d	ä->1	
rer e	f->1	l->1	
rer f	ö->2	
rer g	ö->1	
rer h	a->1	ä->1	ö->1	
rer i	 ->7	n->1	
rer k	a->1	
rer m	e->1	i->1	
rer o	c->14	m->4	
rer p	å->1	
rer s	o->24	å->2	
rer u	n->1	
rer v	a->1	
rer ä	n->2	
rer å	t->1	
rer! 	F->1	
rer, 	a->2	e->2	f->1	i->2	m->1	n->1	o->2	s->1	t->2	u->1	ä->2	
rer.D	e->6	
rer.E	u->2	
rer.J	a->1	
rer.K	o->1	
rer.P	r->1	
rer.T	i->2	
rer.V	i->3	
rera 	a->1	d->12	e->1	f->2	g->1	i->1	j->1	k->2	m->8	o->3	p->1	s->5	t->1	v->1	
rerad	 ->8	e->5	
rerar	 ->12	
reras	 ->12	.->3	
rerat	 ->4	;->1	s->3	
rerin	g->19	
rerna	 ->23	,->6	.->5	;->1	s->6	
rerog	a->1	
rers 	f->1	
reröv	r->1	
res a	n->1	t->1	
res d	ö->1	
res e	l->1	
res f	ö->1	
res i	n->2	
res l	e->3	o->1	
res n	a->1	
res o	c->1	f->1	
res p	o->1	
res r	y->1	ä->1	ö->2	
res v	ä->1	
res å	t->1	
res ö	g->1	
res, 	W->1	j->1	o->1	
resa 	d->1	e->1	f->1	i->3	m->1	o->2	p->1	t->1	ö->1	
resa,	 ->2	
resa.	J->1	
resan	 ->1	
resat	s->6	
resen	t->48	
reser	 ->3	v->6	
resid	e->9	u->1	
reskr	e->1	i->27	
resla	g->24	
reslo	g->11	
reslå	 ->15	r->38	s->16	
resol	u->100	
reson	a->1	e->3	
resor	 ->1	
resp.	 ->2	
respe	g->1	k->80	
respo	,->1	n->2	s->1	
respr	å->9	
ress 	p->3	s->1	
ressa	d->1	n->22	r->1	
resse	 ->21	,->5	.->3	?->1	n->60	r->13	t->5	
ressi	o->1	v->3	
ressk	o->2	
ressm	e->1	
ressn	i->1	
rest 	a->1	t->1	
resta	n->1	s->1	t->3	u->1	
reste	l->3	n->3	r->6	
resti	e->1	
restn	i->1	
restr	i->4	
rests	.->1	
restä	l->9	
restå	e->6	
resul	t->111	
resur	s->50	
resät	t->1	
ret (	C->1	
ret -	 ->2	
ret 1	9->10	
ret a	t->4	v->2	
ret b	e->1	
ret e	x->1	
ret f	a->1	i->1	å->1	ö->27	
ret g	a->1	e->1	
ret h	a->2	o->1	
ret i	 ->7	n->2	
ret k	a->1	o->1	r->1	
ret l	i->1	ä->1	
ret o	c->13	
ret p	l->1	å->1	
ret r	e->1	ö->1	
ret s	k->3	l->1	o->1	ä->2	
ret t	i->6	
ret u	p->1	t->2	
ret v	a->1	
ret ä	n->1	r->5	v->1	
ret å	l->1	
ret ö	v->1	
ret, 	d->1	f->2	i->2	o->3	s->1	v->2	
ret. 	D->1	
ret.D	e->5	
ret.E	f->1	
ret.F	ö->1	
ret.I	 ->1	
ret.J	a->4	
ret.L	å->1	
ret.M	i->1	
ret.T	u->1	y->1	
ret.V	i->2	
ret: 	k->1	
reta 	a->2	b->1	d->1	e->1	f->10	h->1	i->1	k->1	o->1	p->5	r->4	t->1	u->1	å->6	
reta,	 ->2	
retag	 ->55	,->14	.->15	a->23	e->66	n->9	s->25	
retan	d->1	
retar	e->1	i->2	
reter	a->2	
retes	s->12	
retis	e->2	k->2	
retor	i->3	
retro	a->11	
reträ	d->73	t->1	
rets 	L->1	f->2	h->2	s->3	
rets,	 ->1	
retsa	r->3	
retse	n->2	
retsl	o->2	
rett 	a->4	m->1	o->1	p->1	s->1	u->2	
rett.	M->1	
retti	o->2	
retto	n->3	
retts	 ->1	
reuro	p->1	
reuss	a->1	
reutb	i->1	
reutv	e->3	
rev d	i->1	ä->1	
rev f	r->1	
rev i	n->1	
rev n	y->1	
rev o	m->1	
rev s	o->1	
rev t	i->2	
rev u	n->1	
rev.F	r->1	
revid	e->17	
revis	i->18	
revli	g->3	
revlå	d->1	
revol	u->1	
revs 	a->1	s->1	u->1	
rextr	e->6	
rey C	a->3	
reyer	 ->2	.->1	
rez, 	u->1	
rfall	 ->1	,->1	.->1	
rfals	k->1	
rfara	n->76	
rfare	n->25	
rfari	t->2	
rfarn	a->1	
rfart	y->1	
rfatt	a->6	n->1	
rfekt	 ->5	.->1	a->1	
rfini	n->1	
rfinn	a->1	s->2	
rfira	r->2	
rfisk	e->1	
rfjol	,->1	
rflut	e->1	n->13	
rflyt	t->6	
rflöd	i->1	
rfode	r->4	
rfoga	 ->1	n->11	r->6	
rfond	e->55	s->3	
rford	e->5	o->1	
rform	 ->1	
rfors	 ->12	,->5	.->4	b->1	
rfrys	n->1	
rfråg	a->11	n->1	o->1	
rfunn	a->1	e->1	
rfäkt	a->1	
rfära	n->1	
rfärg	,->1	
rfärl	i->1	
rfång	 ->1	
rfölj	a->5	e->3	
rföll	 ->2	
rför 	-->1	2->1	7->1	C->1	E->2	K->1	W->1	a->51	b->18	d->9	e->3	f->11	g->6	h->12	i->18	j->6	k->28	l->1	m->25	n->3	o->6	p->4	r->9	s->25	t->9	u->8	v->30	y->1	ä->23	å->2	ö->1	
rför,	 ->8	
rför.	.->1	
rför:	 ->2	
rför?	D->1	F->1	Ä->1	
rföra	 ->2	s->3	
rförd	e->1	
rföre	n->2	t->2	
rföri	n->12	
rförm	å->1	
rfört	e->2	s->1	
rförv	ä->1	
rg Ha	i->14	
rg av	 ->1	
rg fi	c->1	
rg fö	r->1	
rg gj	o->1	
rg i 	f->1	
rg kr	i->1	
rg me	d->2	
rg oc	h->1	
rg om	 ->7	
rg sa	t->1	
rg ti	l->1	
rg ut	t->1	
rg öp	p->1	
rg, B	r->1	
rg, I	l->1	
rg, f	a->1	
rg, j	u->1	
rg, k	l->1	
rg, s	o->1	
rg.De	t->1	
rg.Ja	g->1	
rg.Le	d->1	
rg.Vi	 ->1	
rga f	ö->1	
rgad 	m->1	
rgan 	a->1	f->1	g->1	i->2	k->1	m->1	p->1	s->7	
rgan"	,->1	
rgan,	 ->6	
rgan.	K->1	
rgane	n->5	t->4	
rgani	 ->1	,->4	s->61	
rgar 	f->1	
rgard	e->1	
rgare	 ->40	,->7	.->7	:->1	n->10	s->7	
rgari	n->1	
rgarn	a->89	
rgars	k->7	
rgavs	 ->2	
rge e	r->1	
rge o	m->1	
rge v	ä->1	å->1	
rge, 	d->1	
rgen 	t->1	
rgens	 ->2	,->1	e->2	k->1	
rger 	a->2	d->2	f->3	h->1	k->1	l->1	r->1	s->2	v->2	
rger,	 ->2	
rger.	 ->1	T->1	
rgerM	e->1	
rgerb	e->1	
rgeri	n->1	
rgerl	i->3	
rges 	i->2	
rges,	 ->1	
rgh.V	i->1	
rgi b	e->1	
rgi g	e->1	ö->1	
rgi h	a->1	
rgi l	e->1	
rgi m	e->1	
rgi o	c->4	
rgi s	o->3	
rgi, 	k->1	o->1	
rgi-,	 ->1	
rgi.A	l->1	
rgi.E	t->1	u->1	
rgi.F	o->1	
rgi.M	a->1	
rgiag	e->1	
rgian	v->6	
rgibe	s->3	
rgice	n->1	
rgief	f->4	
rgifo	r->1	
rgift	e->2	
rgifö	r->4	
rgiim	p->1	
rgika	p->1	
rgiko	n->1	
rgikä	l->37	
rgimi	x->1	
rgimy	n->1	
rgin 	f->1	o->1	u->1	
rgin,	 ->1	
rgina	l->6	
rgior	g->2	
rgipo	l->1	t->1	
rgipr	o->5	
rgise	k->4	
rgisk	t->1	
rgisn	å->1	
rgisä	k->7	
rgive	n->4	
rgivl	i->1	
rgivn	a->3	
rgizi	s->5	
rgiäk	e->1	
rgiåt	e->1	
rglig	a->2	t->1	
rglöm	m->2	
rgmäs	t->2	
rgne 	f->1	
rgo s	o->1	
rgon 	a->2	b->1	d->1	e->2	j->1	k->17	l->1	s->1	ä->1	
rgon,	 ->2	
rgon.	A->1	D->1	H->1	J->1	V->2	
rgond	a->2	
rgot 	W->1	
rgrip	a->14	
rgrun	d->3	
rgrup	p->1	
rgräv	a->3	e->1	
rgsfu	l->1	
rgume	n->17	
rgäll	n->1	
rgäve	s->1	
rgå t	i->1	
rgång	 ->1	a->1	e->2	s->8	
rgår 	j->1	l->1	m->1	n->1	o->1	t->1	
rgått	 ->1	
rgör 	m->1	v->1	
rgöra	 ->10	n->3	
rgörs	 ->2	
rhand	 ->8	,->1	.->1	e->1	l->79	s->8	
rhast	a->3	
rhave	r->1	
rhead	-->1	
rhet 	R->1	S->1	a->3	b->5	d->6	e->4	f->13	g->1	h->5	i->17	k->2	m->5	n->4	o->52	p->3	r->1	s->5	t->8	u->2	v->5	ä->2	
rhet,	 ->12	
rhet.	(->1	A->1	D->9	E->1	F->1	H->1	I->1	N->2	O->4	S->2	T->1	V->3	
rhet?	K->1	N->1	S->1	
rhetJ	a->1	
rhete	n->54	r->3	
rhets	 ->1	-->1	a->1	b->1	e->3	f->5	g->3	k->2	l->1	m->8	n->4	o->1	p->6	r->20	s->4	v->2	
rheug	e->2	
rhind	r->31	
rhist	o->1	
rholk	a->4	
rhopp	n->12	
rhund	r->7	
rhus 	o->1	
rhus,	 ->1	
rhuse	t->1	
rhämt	a->1	n->1	
rhän;	 ->1	
rhäng	a->2	
rhågo	r->2	
rhåll	 ->2	.->1	a->57	e->3	i->3	n->2	s->2	
rhögh	e->2	
rhöll	 ->4	
rhörd	 ->2	a->1	
rhört	 ->9	
ri - 	s->1	
ri 19	9->4	
ri 20	0->5	
ri 8 	b->1	o->1	
ri La	n->3	
ri Va	t->1	
ri av	s->1	
ri be	f->1	
ri di	r->1	
ri en	 ->1	
ri et	t->1	
ri fr	å->1	
ri fö	r->4	
ri i 	T->1	e->1	k->1	
ri in	l->3	t->1	
ri ko	n->2	s->1	
ri me	d->1	
ri mo	t->1	
ri må	n->1	
ri nä	r->2	
ri oc	h->11	
ri om	 ->1	
ri rö	r->8	
ri se	r->1	
ri sk	a->1	
ri so	m->6	
ri va	r->2	
ri är	 ->2	
ri ök	a->1	
ri öp	p->1	
ri!He	r->1	
ri, d	å->1	
ri, e	f->1	
ri, l	i->1	j->1	
ri, m	e->2	i->2	
ri, n	e->1	
ri, o	b->1	c->4	
ri, s	i->1	k->1	å->1	
ri, t	.->2	
ri, u	t->1	
ri, v	a->1	
ri- o	c->10	
ri.Bå	d->1	
ri.Hu	r->1	
ri.Ja	g->1	
ri.Li	k->1	
ri.Ma	n->1	
ri.Vi	d->1	
ria -	 ->1	
ria P	a->1	
ria a	l->1	t->1	
ria d	a->1	e->1	
ria f	r->1	u->1	
ria i	 ->1	n->1	
ria m	a->1	
ria o	c->2	m->1	
ria r	ö->10	
ria s	a->1	o->1	
ria t	i->1	
ria v	a->3	ä->1	
ria å	t->1	
ria, 	d->1	e->1	o->1	r->1	
ria.D	e->1	
ria.Ä	n->1	
rial 	-->1	f->2	i->1	k->1	n->1	o->2	s->3	t->1	
rial,	 ->2	
rial.	D->2	F->1	J->1	S->1	
riale	n->1	t->3	
riane	 ->2	,->1	
rias 	f->3	
riat 	f->1	h->1	
riat.	M->1	
riati	s->2	
ribek	ä->4	
ribla	n->6	
ribut	i->1	
richt	 ->2	.->1	f->3	
ricio	 ->1	
ricit	e->1	
ricka	,->1	
ricke	r->2	t->1	
rickf	r->1	
rickn	i->1	
ricks	v->1	
rid i	 ->1	
rid m	e->7	o->1	
rid s	t->1	
rid, 	h->1	
rid.E	n->1	
rida 	i->1	k->2	m->2	s->1	
ridan	d->13	
ridas	 ->1	
ridd 	m->1	ä->1	
riden	 ->2	
rider	 ->23	.->1	
ridig	a->1	
ridis	k->30	
ridit	s->1	
ridli	g->1	
ridni	n->15	
ridor	e->2	
rids 	m->1	p->1	t->1	u->1	
rie C	u->1	
rie-s	t->1	
riefi	n->1	
riell	 ->4	a->9	t->2	
riels	e->6	
rien 	a->2	b->1	e->1	h->4	i->1	n->1	o->3	s->5	t->1	ä->2	
rien,	 ->4	
rien.	D->1	F->1	H->1	O->1	S->1	U->1	
rienf	r->1	
riens	 ->3	
rient	e->6	
rier 	-->1	f->1	g->1	i->1	k->3	m->1	o->11	p->1	s->8	u->1	ö->1	
rier,	 ->5	
rier.	.->1	D->2	L->1	M->1	
riera	d->1	r->1	
riern	a->18	
riesm	i->1	
riet 	i->1	m->1	o->1	s->1	ä->1	
riet"	.->1	
riet,	 ->2	
riet.	D->1	M->1	V->1	
riets	 ->2	
rifer	a->4	i->1	t->1	
rifie	r->1	
rifin	-->1	
rifrå	g->4	n->2	
rift 	a->1	f->1	o->2	
rift.	 ->1	
rifte	n->1	r->12	
rifti	g->1	
riftl	i->8	
rifts	-->1	f->1	ä->1	
rig a	r->1	t->3	v->1	
rig b	l->1	
rig d	e->1	
rig f	å->2	ö->15	
rig h	a->2	ä->1	
rig i	 ->1	n->2	
rig k	a->2	o->3	
rig m	e->6	y->1	
rig o	c->1	m->1	
rig p	e->1	å->1	
rig r	u->1	
rig s	a->1	o->2	ä->1	
rig t	i->2	v->1	
rig v	a->2	i->1	
rig ä	r->1	
rig å	s->1	
rig".	E->1	
rig, 	a->1	d->1	m->1	o->1	
rig.J	a->1	
riga 	E->2	a->1	b->12	e->1	f->12	g->3	h->1	i->3	k->3	l->2	m->2	o->1	p->7	r->1	s->3	u->3	v->3	ä->4	
riga,	 ->3	
riga.	A->2	H->1	I->1	
rige 	i->1	o->3	p->1	s->1	
rige.	 ->1	J->1	
rigen	 ->17	,->2	o->19	
riger	a->1	
riget	 ->5	.->3	s->4	
righe	t->51	
right	 ->2	s->1	
rigin	a->1	e->1	
rigjo	r->1	
rigor	ö->4	
rigsh	e->1	
rigss	k->1	
rigt 	a->5	b->3	e->1	f->1	h->4	i->3	k->4	l->1	m->1	o->5	p->8	s->3	t->2	v->1	ö->1	
rigt,	 ->3	
rigt.	J->1	
rigör	a->4	s->1	
rihan	d->2	
rihet	 ->44	,->38	.->5	:->1	;->1	e->25	s->2	
rik e	t->1	
rik i	 ->2	n->1	
rik n	ä->2	
rik p	o->1	
rik, 	i->1	u->1	
rik.F	a->1	
rik.G	e->1	
rika 	b->2	d->4	e->2	f->2	g->2	h->2	i->1	m->3	o->5	r->3	s->2	t->2	u->1	v->2	ä->1	ö->2	
rika,	 ->8	
rika-	o->1	
rika.	J->2	P->1	V->2	
rikan	d->2	e->5	s->10	
rikar	 ->1	e->4	n->5	
rikas	 ->8	t->3	
rike 	(->1	-->3	a->3	b->3	d->1	e->4	f->2	g->2	h->2	i->4	k->3	m->4	n->1	o->10	s->7	t->1	v->2	ä->3	
rike,	 ->15	
rike.	 ->1	.->2	D->5	F->2	I->1	J->2	M->1	N->1	O->1	V->3	Ö->1	
rike:	 ->1	
rikeE	n->1	
rikeF	r->1	
rikeN	ä->1	
riked	o->10	
riker	 ->10	,->1	n->2	
rikes	 ->26	-->4	f->4	h->4	m->9	p->3	
riket	 ->6	,->3	.->2	s->6	
rikis	k->49	
rikli	g->2	
rikom	m->1	
rikon	v->1	
rikt 	b->1	e->2	f->1	h->1	k->1	l->1	o->3	r->1	s->4	
rikt,	 ->1	
rikt.	B->1	I->1	
rikta	 ->19	,->1	.->1	d->14	n->1	r->8	s->3	t->13	
rikti	g->45	o->4	v->1	
riktl	i->70	
riktn	i->50	
riktp	u->2	
ril 1	9->1	
ril f	ö->1	
ril u	t->1	
ril.J	a->1	
rilag	s->1	
rilan	k->1	
rilik	n->1	
riljo	n->1	
rilob	b->1	
rimin	a->4	e->23	
rimit	i->1	
rimli	g->23	
rimma	r->1	
rimsa	v->2	
rimsb	e->2	
rimsp	a->1	
rimsr	å->2	
rimså	t->1	
rimål	,->1	
rin a	b->1	t->2	
rin b	e->1	
rin e	n->1	t->1	
rin f	o->1	å->1	ö->3	
rin h	a->1	
rin i	 ->4	
rin k	o->2	r->1	
rin l	ö->1	
rin m	e->1	
rin o	c->6	
rin p	å->1	
rin s	j->1	k->2	o->3	p->1	t->1	å->1	
rin v	i->2	
rin ä	n->1	r->1	
rin!H	e->1	
rin, 	d->1	f->1	g->2	h->1	m->1	o->1	p->1	s->4	t->1	v->2	
rin. 	D->1	M->1	
rin.D	e->2	ä->1	
rin.H	e->1	
rin.I	n->1	
rin.J	a->2	
rin.N	ä->1	
rin.S	a->1	t->1	
rin.V	a->1	i->2	
rin: 	e->1	
rin?P	a->1	
rinci	p->194	
rindu	s->2	
rinfö	r->4	
ring 	-->4	2->2	6->1	8->2	E->1	F->1	a->106	b->3	d->1	e->7	f->20	g->4	h->3	i->28	k->6	l->3	m->9	o->34	p->10	r->2	s->27	t->8	u->2	v->6	ä->10	
ring!	J->1	
ring"	 ->2	
ring)	 ->1	
ring,	 ->39	
ring.	 ->2	A->1	D->10	E->2	F->4	H->2	I->3	J->4	K->1	L->1	M->3	N->4	O->2	P->2	S->1	T->2	V->6	Ä->1	
ring;	 ->2	
ring?	D->1	H->1	O->1	
ringa	 ->11	.->1	d->1	n->2	r->172	s->1	t->3	
ringe	n->142	
ringg	å->2	
rings	 ->2	-->2	a->4	b->15	c->8	d->2	f->210	i->1	k->152	l->10	m->5	n->1	o->4	p->13	r->1	s->23	t->1	v->4	
ringå	n->1	
rinho	 ->4	.->1	s->1	
rinip	e->1	
rinna	 ->1	
rino 	i->1	k->1	o->1	
rino,	 ->1	
rino.	J->1	O->1	
rinos	 ->1	
rinra	 ->11	r->1	s->1	
rinre	s->1	
rinrä	t->1	
rins 	a->2	d->1	i->2	j->1	k->1	s->2	
rinse	e->1	
rinst	i->8	
rinta	g->1	
rinte	l->5	
rinär	e->1	f->1	p->1	
rio f	ö->1	
rio u	t->1	
riod 	a->2	d->2	f->4	i->4	k->1	o->1	p->2	r->2	s->2	v->1	ä->2	
riod,	 ->5	
riod.	D->1	V->1	
riod?	-->1	
riode	n->39	r->2	
riodi	s->14	
rior.	D->1	
riori	 ->3	t->36	
riot 	i->1	s->1	
rioti	s->1	
ripa 	a->1	d->3	e->2	i->3	m->1	o->2	p->1	t->2	
ripa,	 ->1	
ripa.	K->1	
ripan	d->19	
ripas	 ->1	
ripen	.->1	
riper	 ->15	
ripet	 ->2	,->1	
ripit	 ->2	
ripli	g->6	
ripna	 ->1	
ripol	i->3	
rips 	a->1	
rirra	 ->1	
ris (	P->1	
ris P	a->1	
ris f	ö->3	
ris h	a->1	ä->1	
ris i	 ->1	n->1	
ris k	o->2	
ris l	a->1	
ris m	å->1	
ris o	c->1	
ris s	o->2	
ris u	p->1	
ris v	a->1	
ris ä	n->1	r->1	
ris å	t->1	
ris, 	i->1	o->1	
ris.J	a->1	
ris.S	a->1	
ris: 	f->1	
ris?Ä	r->1	
risa 	d->1	
risdi	k->5	
risek	t->2	
risen	 ->3	.->3	
riser	 ->6	,->1	.->2	a->4	i->3	n->4	
rises	 ->2	
riset	 ->6	.->1	
risfö	r->1	
risk 	-->1	a->3	b->1	d->2	e->1	f->3	j->1	k->1	l->1	m->2	o->1	p->1	s->3	u->3	
risk,	 ->3	
risk.	V->1	
riska	 ->28	,->2	b->1	n->2	
riskb	e->4	
riske	 ->1	n->16	r->37	
riskf	a->1	r->1	y->1	ö->1	
riskh	a->6	
riskk	a->1	o->2	
riskn	i->1	
riskt	 ->9	
risku	p->1	
riskv	ä->3	
rislä	p->2	
rism 	m->1	o->8	s->1	u->1	
rism,	 ->4	
rism.	D->3	F->1	O->1	V->2	
risme	d->2	n->6	
risni	v->1	
risom	r->1	
rison	t->3	
rissi	t->1	
risst	y->1	
rissä	n->1	
rist 	f->3	p->19	s->1	u->1	ä->1	
rista	l->2	n->12	t->1	
ristd	e->11	
riste	n->12	r->33	
ristf	ä->8	
risth	a->1	
risti	g->1	n->1	s->2	
rists	e->2	
ristä	l->1	
ristå	e->1	
risut	v->1	
rit a	k->1	v->1	
rit b	i->1	ä->1	
rit d	ä->1	
rit e	f->1	n->10	t->2	
rit f	a->1	e->1	r->2	ö->3	
rit g	a->1	
rit h	a->1	ä->1	ö->1	
rit i	n->5	
rit k	o->2	ä->2	
rit l	e->1	å->1	
rit m	i->2	o->1	y->1	ä->1	ö->3	
rit n	å->1	ö->1	
rit o	c->1	e->1	
rit p	e->1	o->1	r->1	å->2	
rit r	i->2	
rit s	n->1	t->3	v->1	ä->1	å->3	
rit t	i->2	y->1	
rit u	n->1	
rit v	a->1	i->1	
ritan	,->1	n->14	s->1	
ritas	,->1	
ritat	i->1	
riter	.->1	a->20	i->36	
ritet	 ->45	,->13	.->10	:->1	?->2	e->32	s->25	
ritik	 ->10	,->1	.->1	e->4	
ritim	a->1	t->2	
ritis	e->10	h->1	k->22	
ritle	k->1	
ritor	i->17	
ritre	a->1	
ritt 	i->2	k->1	
ritt,	 ->1	
ritt.	M->1	
ritte	r->2	
ritti	n->1	s->16	
rium 	a->1	m->1	s->2	
rium,	 ->3	
rium.	A->1	D->1	H->1	P->1	R->1	
riuts	k->1	
riva 	b->1	d->9	e->7	g->1	h->1	i->2	k->3	n->1	p->2	s->1	t->1	u->1	
rivan	d->3	
rivas	 ->2	.->1	
rivat	 ->1	.->1	a->16	e->1	i->2	
rivbo	r->1	
rivel	s->5	
riven	 ->9	
river	 ->20	,->1	.->1	
rivet	 ->7	
rivil	e->6	i->1	l->12	
rivit	 ->5	s->3	
rivkr	a->3	
rivna	 ->4	
rivni	n->5	
rivs 	a->2	e->2	g->1	i->6	s->1	ö->1	
rivs,	 ->1	
rivs.	D->1	
riäre	r->3	
riärp	l->1	
rière	 ->1	
riös 	o->1	
riösa	 ->2	,->1	
riöst	 ->4	
rja a	n->2	r->3	t->2	
rja d	e->1	
rja e	f->1	t->1	
rja f	u->1	ö->7	
rja k	l->1	o->1	
rja m	e->35	i->2	
rja o	m->1	
rja p	å->3	
rja r	e->1	
rja s	i->1	
rja t	i->2	ä->1	
rja u	t->1	
rja å	t->1	
rjade	 ->9	s->1	
rjan 	a->6	d->1	e->2	h->2	i->2	p->2	t->1	u->1	
rjan,	 ->2	
rjar 	b->3	d->1	f->1	g->1	m->3	n->1	o->2	p->1	s->2	t->1	
rjar.	D->1	
rjat 	-->1	f->1	j->1	l->1	s->3	t->1	v->1	
rjat.	I->1	J->1	
rjats	,->1	
rjde 	a->1	
rje 1	0->1	
rje E	U->1	
rje a	n->2	v->1	
rje b	e->1	i->1	o->1	
rje d	a->7	e->1	i->1	
rje e	n->5	u->2	
rje f	a->6	o->6	r->1	ö->2	
rje g	e->1	å->4	
rje h	a->2	
rje i	n->3	
rje k	o->1	u->1	
rje l	a->9	
rje m	e->9	å->2	
rje o	a->1	
rje r	e->2	ä->1	
rje s	a->1	o->1	t->3	u->1	
rje å	r->9	t->1	
rjer 	f->2	
rjnin	g->4	
rk - 	d->1	o->1	
rk at	t->1	
rk be	t->1	
rk by	g->1	
rk da	g->1	
rk el	l->2	
rk en	i->1	
rk fi	n->1	
rk få	r->1	
rk fö	r->3	
rk ge	n->1	
rk ha	r->1	
rk i 	A->1	T->1	d->1	f->1	g->1	m->1	
rk in	o->1	t->4	
rk ka	n->1	
rk ko	m->1	n->2	
rk kä	n->1	
rk ly	c->1	
rk me	d->2	
rk må	s->1	
rk oc	h->6	
rk of	f->1	
rk po	l->2	
rk på	 ->3	
rk se	n->1	
rk sk	a->2	
rk so	m->5	
rk så	d->1	
rk ti	l->2	
rk tr	o->1	
rk ut	v->1	
rk vi	d->1	l->1	n->1	t->1	
rk är	 ->2	
rk, d	å->1	
rk, g	o->1	å->1	
rk, m	e->1	
rk, o	c->1	
rk, s	o->1	
rk, ä	r->1	
rk-da	m->1	
rk.Be	t->1	
rk.De	t->2	
rk.Då	 ->1	
rk.Fr	å->1	
rk.Ja	g->1	
rk.Sy	r->1	
rk.Va	n->1	
rk?Re	g->1	
rka -	 ->2	
rka 1	7->1	
rka 2	5->1	
rka E	u->1	
rka a	l->1	r->1	v->1	
rka b	i->1	o->1	
rka d	e->7	i->1	
rka e	n->2	
rka f	ö->11	
rka h	e->1	u->1	
rka i	 ->6	n->3	
rka k	a->1	o->3	u->2	
rka l	o->1	
rka m	a->1	e->2	i->1	
rka n	ä->2	
rka o	c->4	r->2	
rka p	o->2	r->1	å->1	
rka r	e->2	i->1	
rka s	a->1	i->1	k->1	o->1	t->2	å->1	
rka t	e->1	i->6	r->2	
rka u	n->1	t->1	
rka v	e->1	å->2	
rka ä	r->1	
rka å	t->1	
rka, 	a->1	d->1	j->1	s->2	
rka.H	e->1	
rkade	 ->2	
rkan 	a->2	d->1	f->1	i->1	m->3	o->2	p->9	s->1	t->1	v->1	ä->1	
rkan,	 ->1	
rkan.	V->1	
rkand	e->3	
rkane	n->3	r->1	
rkans	 ->1	
rkant	 ->2	.->1	
rkapi	t->1	
rkar 	a->1	b->1	d->11	f->1	h->5	i->6	k->2	l->1	m->6	n->1	o->1	p->1	r->3	s->6	t->1	u->2	v->6	ä->1	ö->3	
rkar,	 ->1	
rkara	n->5	
rkare	 ->13	,->3	.->1	n->12	s->2	
rkarn	a->35	
rkas 	a->5	f->1	l->1	n->1	p->2	
rkas,	 ->1	
rkas.	I->1	
rkass	o->2	
rkast	 ->1	a->10	e->4	n->1	
rkat 	-->1	h->1	o->1	
rkat,	 ->1	
rkata	s->13	
rkate	g->2	
rkats	 ->3	.->1	?->1	
rkbar	 ->1	a->1	t->1	
rkbor	r->1	
rkdam	m->1	
rke i	 ->2	
rke m	a->1	
rke t	i->5	
rkefö	r->1	
rkel 	n->1	
rkels	e->5	
rken 	G->1	a->2	b->2	f->3	g->1	i->3	j->1	k->1	m->4	o->2	p->3	r->1	s->2	u->2	ä->1	
rken,	 ->1	
rken.	D->1	
rkepo	s->1	
rker 	a->1	d->4	n->1	v->1	
rkera	 ->2	d->1	r->2	t->2	
rkeri	n->3	
rkesa	r->1	
rkese	t->1	
rkesf	ö->1	
rkesk	a->1	v->1	
rkesl	a->2	i->2	
rkesm	ä->1	
rkesu	t->7	
rkesv	a->1	
rket 	G->1	b->2	e->1	f->4	g->1	h->3	i->3	k->1	l->1	m->1	o->2	p->1	s->4	t->1	u->3	v->2	ä->3	
rket,	 ->6	
rkets	 ->2	
rki.D	e->1	
rkiet	 ->27	,->2	.->2	s->4	
rkilt	 ->1	
rkin 	o->1	
rkin.	D->1	
rkisk	 ->1	a->5	e->1	
rkiv 	l->1	
rkive	r->1	
rkki 	L->2	
rklag	a->6	
rklar	 ->2	a->52	i->24	
rklas	s->1	
rklig	 ->10	a->38	e->126	h->20	t->16	
rklyv	e->1	
rkläg	g->1	
rkmen	i->2	
rknad	 ->8	,->6	.->2	e->146	s->29	
rknin	g->35	
rknip	p->3	
rkogå	r->1	
rkoll	e->1	
rkoma	n->1	
rkomm	a->5	e->1	
rkoms	t->1	
rkonf	e->1	
rkont	r->2	
rkop 	b->1	
rkor 	s->1	
rkor,	 ->1	
rkort	a->1	n->1	
rkoti	k->7	
rkov 	n->1	
rkran	s->1	
rkrom	a->1	
rkräv	a->1	
rks b	e->1	
rks g	e->1	
rks o	c->1	m->1	
rks t	i->1	
rks.D	ä->1	
rks.O	L->1	
rks.V	i->1	
rksam	 ->4	h->82	m->12	t->6	
rksan	l->1	
rkstä	l->19	
rkt E	u->3	
rkt a	r->2	v->1	
rkt b	e->5	i->1	
rkt c	h->1	
rkt d	e->1	o->1	
rkt e	x->1	
rkt f	r->1	ö->1	
rkt i	n->2	
rkt k	o->1	
rkt m	a->1	i->4	
rkt o	c->2	
rkt p	o->2	
rkt r	e->2	
rkt s	a->1	t->5	
rkt v	a->1	
rkt ö	v->3	
rkt, 	f->1	
rkt.D	e->2	
rkta 	a->2	b->8	e->1	i->2	k->1	p->2	r->2	
rkts 	u->1	
rktyg	 ->6	?->1	s->1	
rkula	t->1	
rkule	r->2	
rkunn	a->2	
rkurs	e->1	
rkänd	 ->3	a->1	e->1	
rkänn	a->22	e->11	s->2	
rkänt	 ->1	s->1	
rkött	s->1	
rl He	i->1	
rl oc	h->1	
rl vo	n->3	
rl-He	i->1	
rlag 	f->2	o->1	t->1	
rlag,	 ->1	
rlag.	B->1	J->1	
rlagd	,->1	
rlage	n->1	
rlago	r->2	
rlagt	 ->1	,->1	s->1	
rlame	n->600	
rland	 ->16	,->1	.->4	e->2	s->2	
rlang	e->6	
rld W	i->1	
rld s	o->1	
rld, 	d->1	s->1	
rld.J	a->1	
rlden	 ->19	,->9	.->3	:->1	?->1	s->4	
rldsd	e->1	
rldse	k->1	
rldsf	r->1	
rldsh	a->4	
rldsk	r->6	
rldsl	i->1	
rldsm	a->1	
rldsn	i->1	
rldso	m->1	
rleda	s->1	
rledi	g->1	
rlega	d->2	
rleke	n->2	
rleva	,->1	?->1	
rleve	r->3	
rlevn	a->4	
rlevs	 ->1	
rlig 	a->1	b->3	e->3	f->3	h->1	k->1	l->1	m->1	n->2	o->5	p->2	r->3	s->1	u->2	
rlig!	H->1	
rlig,	 ->4	
rlig.	D->1	G->1	
rlig:	 ->1	
rliga	 ->63	,->1	.->1	;->1	r->54	s->3	
rlige	n->56	
rligg	a->1	
rligh	e->26	
rligt	 ->76	,->2	.->4	v->95	
rlika	 ->1	r->1	
rlikn	i->44	
rlin 	1->1	f->1	o->1	u->1	
rlin,	 ->2	
rlin.	O->1	
rling	 ->1	.->1	
rlist	e->2	
rlita	 ->2	r->4	
rlitl	i->4	
rliv,	 ->1	
rliv.	V->1	
rliva	 ->2	d->1	n->7	s->5	t->4	
rlora	 ->3	d->5	r->4	t->8	
rlsru	h->2	
rlund	a->3	
rlust	 ->1	.->1	b->1	e->7	
rlyse	r->1	
rlyst	 ->1	
rlägg	a->3	n->6	
rlägs	e->2	
rläkt	a->1	
rlämn	a->18	
rländ	a->2	e->16	s->18	
rläng	a->1	n->3	
rlärl	i->1	
rlätt	a->18	
rlåta	 ->5	n->1	s->1	
rlåte	n->3	
rlåti	t->2	
rlåtl	i->2	
rlåts	 ->1	
rlöst	,->1	a->1	
rløn,	 ->2	
rm at	t->2	
rm av	 ->24	
rm be	s->1	
rm da	m->1	
rm dö	l->1	
rm el	-->4	l->1	
rm fö	r->3	
rm i 	s->3	
rm ju	s->1	
rm ka	n->1	
rm ko	m->1	n->1	s->1	
rm lö	p->1	
rm oc	h->3	
rm på	 ->1	
rm sk	a->2	
rm so	m->4	
rm sp	r->1	
rm vi	 ->1	d->1	
rm vä	c->1	
rm är	 ->1	
rm öv	e->1	
rm, e	f->1	n->1	
rm, f	ö->1	
rm, m	e->1	
rm, o	p->1	r->1	
rm, s	o->1	
rm, u	t->1	
rm, ä	r->1	
rm-el	-->1	
rm.De	t->1	
rm.EG	-->1	
rm.Me	n->1	
rm.Nu	 ->1	
rm.Sa	m->1	
rm.Vi	 ->1	
rm.Är	 ->1	
rm: e	n->1	
rma M	a->1	
rma b	e->1	i->1	ä->1	
rma d	e->2	i->1	
rma e	n->1	
rma f	ö->3	
rma k	l->1	o->3	
rma m	a->2	o->1	
rma p	r->1	
rma s	i->2	k->1	u->1	v->2	
rma u	t->1	
rma v	å->1	
rma å	r->1	
rma ö	v->1	
rma.O	r->1	
rmace	u->1	
rmade	 ->5	
rmajo	r->1	
rmako	l->1	
rmala	 ->2	
rmali	s->3	t->1	
rmalt	 ->3	.->2	
rman 	R->1	
rman.	K->1	
rmand	e->5	i->1	
rmane	n->8	
rmans	 ->1	t->1	
rmar 	i->2	n->1	o->4	p->1	s->3	ö->1	
rmarb	e->3	
rmare	 ->15	
rmarn	a->13	
rmas 	a->1	p->1	s->1	
rmast	 ->1	,->1	e->11	
rmat 	a->1	f->1	u->6	
rmate	r->1	
rmati	o->72	v->2	
rmats	 ->1	
rmed 	a->2	b->2	e->3	f->6	i->4	k->8	l->1	m->2	o->4	p->2	r->1	s->4	t->2	u->1	v->1	ä->1	ö->3	
rmed,	 ->2	
rmedl	a->3	
rmell	 ->1	a->4	t->11	
rmels	e->1	
rmen 	a->6	i->1	k->2	o->1	r->2	s->1	
rmen,	 ->2	
rmen.	F->1	J->2	
rmena	n->2	
rmeni	n->1	
rmens	 ->5	
rmer 	a->12	f->13	g->1	h->1	i->2	k->3	l->2	m->1	o->5	p->4	s->11	v->1	ä->1	
rmer,	 ->4	
rmer.	D->5	F->1	H->1	I->1	M->1	O->1	S->1	T->1	
rmera	 ->18	d->3	r->1	s->4	
rmeri	n->17	
rmern	a->18	
rmfäl	l->1	
rmför	s->2	
rmidd	a->12	
rmine	r->1	
rmini	s->10	
rminn	e->1	
rmis.	F->1	
rmist	i->1	
rmnin	g->31	
rmo, 	H->1	
rmod 	e->1	
rmodi	g->1	
rmodl	i->12	
rmonb	e->1	
rmoni	 ->1	s->17	
rmorg	o->1	
rmout	i->1	
rmpak	e->1	
rmpro	c->10	g->3	j->1	
rmrap	p->2	
rmsig	n->2	
rmsta	d->1	
rmstä	m->1	
rmt a	n->1	r->1	t->1	
rmt d	e->1	
rmt e	k->1	r->1	
rmt h	å->1	
rmt m	y->1	
rmt o	m->3	
rmt t	a->5	
rmt u	n->1	
rmt v	i->1	ä->1	
rmule	r->18	
rmynd	a->1	i->14	
rmäss	i->1	
rmå b	e->1	
rmå r	å->1	
rmåga	 ->19	,->2	.->2	n->8	
rmåli	g->1	
rmån 	f->11	
rmåne	r->2	
rmåns	p->1	
rmår.	L->1	
rmåtg	ä->1	
rmé o	c->1	
rmén 	o->1	
rmén.	W->1	
rmögn	a->1	
rmöte	 ->2	
rn (f	o->1	
rn - 	a->1	d->1	f->1	s->1	
rn Er	i->2	
rn bi	l->1	
rn bö	r->1	
rn de	b->1	
rn dä	r->1	
rn el	l->1	
rn en	 ->1	l->1	
rn fi	n->1	
rn fo	r->1	
rn fr	o->1	
rn fö	r->7	
rn gr	ä->1	
rn ha	f->1	r->2	
rn i 	E->2	d->2	
rn in	n->1	t->1	
rn ka	n->1	
rn ko	m->3	n->1	
rn li	b->1	v->1	
rn me	n->1	
rn ny	l->1	
rn oc	h->14	
rn om	 ->2	
rn på	 ->1	
rn re	m->1	
rn sa	m->2	
rn sk	a->2	u->1	
rn so	m->3	
rn st	y->1	
rn sä	r->1	
rn så	 ->2	
rn ta	l->1	
rn to	g->1	
rn un	d->2	
rn va	d->1	
rn vi	d->1	
rn är	 ->3	
rn).D	e->1	
rn, B	r->1	
rn, R	o->1	
rn, a	r->1	
rn, e	t->1	
rn, f	å->1	
rn, h	a->1	
rn, i	 ->1	n->4	
rn, j	a->1	
rn, m	a->1	e->2	u->1	
rn, o	c->2	f->1	
rn, s	a->1	o->1	å->1	
rn, v	i->2	
rn- o	c->2	
rn.) 	H->1	
rn.. 	D->1	
rn.De	t->7	
rn.Dä	r->1	
rn.Fö	r->3	
rn.He	r->2	
rn.Ja	g->1	
rn.Ju	s->1	
rn.Ko	r->1	
rn.Mi	n->1	
rn.Om	 ->1	
rn.Vi	s->1	
rn.Ög	o->1	
rn/No	r->2	
rn?An	s->1	
rna (	K->1	
rna -	 ->18	
rna 1	 ->2	2->1	3->1	6->1	
rna 3	3->1	
rna 6	 ->1	
rna 8	1->4	5->3	7->1	
rna A	z->1	
rna I	X->1	
rna P	r->1	
rna T	u->1	
rna a	b->1	d->1	l->1	n->10	r->1	t->35	v->46	
rna b	e->10	i->3	l->8	o->5	y->1	ö->6	
rna d	e->4	i->5	o->1	r->4	ä->11	å->3	
rna e	f->1	l->9	m->4	n->6	r->1	t->3	u->1	x->2	
rna f	a->2	i->3	o->5	r->33	å->12	ö->132	
rna g	e->11	i->1	j->3	r->3	ä->2	å->2	ö->8	
rna h	a->43	e->4	o->3	u->1	ä->3	å->2	ö->4	
rna i	 ->171	b->1	n->33	
rna j	u->2	ä->1	
rna k	a->14	l->1	n->1	o->21	r->3	u->5	ä->3	
rna l	a->1	e->2	i->3	j->1	ä->1	å->1	ö->1	
rna m	a->2	e->51	i->1	o->2	y->1	å->17	ö->1	
rna n	a->1	r->2	y->1	ä->8	å->2	
rna o	c->143	m->38	r->2	s->1	
rna p	a->2	e->1	o->1	r->1	u->1	å->28	
rna r	e->7	ä->3	ö->2	
rna s	a->3	e->10	i->1	j->5	k->42	l->2	n->1	o->48	p->2	t->6	v->1	y->1	ä->3	å->3	ö->1	
rna t	.->1	a->8	i->41	o->2	r->1	v->1	y->1	
rna u	n->10	p->14	r->1	t->14	
rna v	a->9	e->4	i->21	ä->1	
rna ä	m->1	n->7	r->43	v->2	
rna å	s->1	t->2	
rna ö	k->2	n->1	v->5	
rna!D	e->1	
rna!H	e->1	
rna!O	m->1	
rna".	D->1	K->1	
rna"i	n->1	
rna, 	S->1	a->12	b->4	d->14	e->12	f->8	g->1	h->9	i->17	j->3	k->3	l->5	m->21	n->5	o->29	p->1	r->3	s->37	t->9	u->9	v->16	ä->2	
rna. 	D->2	K->1	S->1	V->1	
rna.(	T->1	
rna.)	B->1	
rna.-	 ->1	
rna..	(->1	
rna.A	l->6	m->1	v->2	
rna.B	e->2	
rna.D	e->58	o->1	ä->4	
rna.E	f->2	m->1	n->1	t->4	u->3	
rna.F	a->2	r->1	ö->12	
rna.G	e->1	i->1	
rna.H	a->1	e->3	u->3	ä->2	
rna.I	 ->11	b->1	n->3	
rna.J	a->23	u->1	
rna.K	a->2	o->8	
rna.L	i->2	å->2	
rna.M	a->1	e->13	i->5	
rna.N	a->1	i->2	u->1	ä->3	
rna.O	c->1	m->3	r->1	
rna.P	r->1	å->4	
rna.R	e->1	
rna.S	e->1	k->1	l->2	o->3	t->1	y->1	å->2	
rna.T	a->2	i->1	r->1	
rna.U	p->1	r->1	t->3	
rna.V	a->3	e->1	i->28	ä->2	å->1	
rna.Ä	n->2	v->1	
rna.Å	 ->1	
rna/s	a->1	
rna: 	F->1	m->1	v->1	
rna; 	j->2	l->1	o->1	
rna?E	t->1	
rna?H	a->1	u->1	
rna?I	 ->1	
rna?J	a->1	o->1	
rna?M	a->1	
rna?V	a->2	i->2	
rna?Ä	r->1	
rnaHe	r->1	
rnade	s->1	
rnage	l->1	
rnali	s->2	
rnamn	,->1	
rnan 	f->1	i->5	
rnar 	d->1	f->2	o->1	
rnard	 ->1	
rnare	 ->1	
rnas 	E->7	a->23	b->4	c->1	d->3	e->5	f->26	g->3	h->3	i->13	k->14	l->6	m->6	n->4	o->19	p->11	r->13	s->28	t->6	u->6	v->9	y->1	ä->1	å->3	ö->1	
rnas,	 ->2	
rnas.	 ->1	
rnati	o->82	v->12	
rnbar	n->1	
rnd L	a->3	
rne o	c->1	
rne, 	E->1	
rnear	v->1	
rnedr	a->2	
rneka	 ->2	,->1	.->1	n->1	r->2	s->1	
rnene	r->8	
rner 	m->1	
rneri	n->2	
rnern	a->1	
rnet 	f->1	n->1	s->1	ä->1	
rnet,	 ->4	
rnet.	D->1	I->1	O->1	
rnfre	d->1	
rnfrå	g->2	
rnhil	l->1	
rnier	 ->11	,->1	s->2	
rning	 ->5	,->3	.->1	a->7	e->5	s->6	
rnise	r->24	
rniti	s->1	
rnivå	.->1	
rnié 	u->1	
rnkat	a->1	
rnkra	f->22	
rnogr	a->2	
rnpor	n->2	
rnpri	n->2	
rnpun	k->2	
rns a	l->1	
rns d	e->1	
rns f	r->2	ö->1	
rns h	i->1	
rns n	y->1	
rns o	c->1	r->1	
rns p	o->2	r->1	
rns s	a->1	i->2	p->1	
rns u	t->1	
rns v	ä->1	
rnste	n->1	
rnstr	å->1	
rnsäk	e->3	
rnt s	j->1	n->1	o->1	
rnt u	t->1	
rnt.S	å->1	
rntek	n->2	
rnten	.->1	
rntun	n->1	
rnuft	 ->1	.->1	e->1	i->11	
rnvap	e->8	
rnväg	 ->8	,->1	.->2	a->1	s->3	
rnya 	m->1	
rnyan	d->1	
rnyar	 ->1	
rnyas	 ->1	
rnyba	r->39	
rnyel	s->6	
rnäte	t->1	
rnödv	ä->1	
rnör,	 ->1	
ro - 	e->1	t->1	
ro 19	9->1	
ro Eu	r->1	
ro at	t->4	
ro be	a->1	
ro bl	a->1	
ro de	t->1	
ro di	s->1	
ro fu	l->1	
ro fö	r->10	
ro ha	r->1	
ro i 	e->1	f->2	h->1	m->1	n->1	
ro le	d->1	
ro me	l->1	
ro må	s->1	
ro nä	r->2	
ro nå	g->3	
ro oc	h->5	
ro om	 ->1	
ro pe	r->2	
ro på	 ->4	
ro so	m->12	
ro ti	l->2	
ro tr	e->1	
ro un	d->1	
ro va	r->1	
ro är	 ->3	
ro äv	e->1	
ro öv	e->1	
ro!Al	l->1	
ro, d	e->1	
ro, f	ö->2	
ro, h	u->1	
ro, k	o->1	
ro, o	c->2	r->1	
ro, s	a->1	o->2	t->1	
ro, t	i->1	
ro, v	i->1	
ro, ä	n->1	
ro-rå	d->1	
ro.At	t->1	
ro.Be	t->1	
ro.De	s->1	t->1	
ro.Dä	r->1	
ro.Fl	e->1	
ro.Fö	r->1	
ro.Hu	r->1	
ro.Ja	g->2	
ro.Kn	a->1	
ro.Nä	r->1	
ro.Om	 ->1	
ro.Se	d->1	
ro.Tr	o->1	
ro.Vi	 ->3	
roa f	ö->1	
roa o	s->1	
roa s	i->1	
road 	ö->3	
roade	 ->2	
roakt	i->12	
roand	e->9	
roans	t->1	
roar 	e->1	k->1	o->1	s->2	
roate	r->1	
roble	m->183	
roced	u->1	
rocen	t->94	
roces	s->109	
rocks	k->1	
rodac	 ->3	"->1	-->1	
rodas	 ->1	.->3	
rodda	.->1	
rodde	 ->8	
roder	s->2	
rodi 	a->3	b->1	h->2	i->1	l->2	o->5	s->1	t->2	
rodi,	 ->1	
rodi.	S->1	V->1	
rodi;	 ->1	
rodis	 ->7	
roduc	e->31	
roduk	t->53	
roedt	e->14	
roeko	n->5	
roend	e->127	
rof -	 ->1	
rof a	v->1	
rof e	l->1	x->1	
rof f	ö->5	
rof h	a->2	
rof i	 ->1	n->2	
rof k	u->1	
rof l	i->1	
rof o	c->2	
rof s	o->4	
rof u	t->1	
rof ä	g->1	
rof, 	h->1	m->1	o->1	s->1	
rof.D	e->1	ä->1	
rof.E	n->1	
rof.J	a->1	
rofal	a->1	
rofdr	a->1	
rofed	e->1	
rofen	 ->13	,->5	.->2	
rofer	 ->17	"->1	,->4	.->5	n->4	
rofes	s->7	
rofhj	ä->1	
rofil	 ->1	.->2	
rofin	a->1	
rofsi	t->1	
rofst	r->1	ö->2	
roför	e->1	
rog a	k->1	
rog f	ö->1	
rog s	i->1	
rog t	i->2	
rogan	s->1	t->1	
rogat	i->1	
rogbe	r->1	
rogen	 ->1	
roger	 ->1	
roget	 ->1	
rogku	l->1	
rogra	m->238	
rogre	s->1	
rogru	n->1	
rogs 	d->1	n->1	
roisk	 ->1	
rojek	t->64	
rojka	n->1	
rojus	t->6	
rok d	e->1	
rok f	ö->2	
rok g	j->1	
rok o	c->1	
rok s	a->1	
rok, 	f->1	k->1	s->1	
rokig	 ->1	t->1	
rokla	m->1	
rokre	d->2	
rol, 	d->1	
rol.M	e->1	
roleu	m->1	
rolig	 ->4	,->1	a->2	e->6	t->5	
roll 	-->1	E->1	a->21	d->2	f->7	g->2	i->17	k->2	m->1	n->3	o->6	p->1	s->10	u->1	v->4	ä->3	ö->5	
roll!	J->1	
roll,	 ->19	
roll-	 ->1	
roll.	D->4	E->1	F->2	H->1	I->2	J->2	K->2	M->1	P->2	S->2	T->2	U->1	V->3	
roll:	 ->1	
rolla	n->1	
rolle	n->26	r->60	
rollf	u->1	
rollm	a->1	y->1	ö->2	
rollo	m->1	r->1	
rolls	y->3	
rollu	t->14	
rollv	e->1	
roläm	p->2	
rom d	a->1	
rom g	ö->1	
rom, 	k->1	
romad	e->1	
romer	 ->1	,->3	a->4	n->1	
romet	 ->1	
romis	s->22	
rområ	d->3	
roms 	f->1	
romsa	 ->3	r->1	
romsv	ä->1	
ron -	 ->1	
ron a	t->1	v->3	
ron e	l->1	
ron f	ö->2	
ron o	c->1	
ron p	å->1	
ron s	k->1	
ron ä	r->1	
ron ö	v->1	
ron, 	h->1	i->1	s->1	
ron- 	o->1	
ronaz	i->1	
ronge	n->1	
roni.	(->1	
ronik	-->1	
ronis	e->1	k->9	
ronju	v->1	
ronmä	r->2	
ronod	l->3	
ronom	i->1	
rons 	s->1	t->1	v->1	
ronta	t->1	
ronte	n->3	
roomr	å->1	
rop o	c->1	m->1	
rop s	k->1	
rop, 	p->1	
rop.S	o->1	
ropa 	-->2	a->7	b->1	d->1	e->4	f->6	h->11	i->9	k->10	m->13	n->1	o->19	p->3	r->2	s->26	t->4	u->4	v->7	ä->11	
ropa!	A->1	F->1	
ropa"	.->1	
ropa,	 ->36	
ropa.	.->2	1->1	D->15	E->2	F->3	H->6	I->2	J->8	M->3	N->1	O->1	P->1	R->1	T->2	U->1	V->10	Ä->1	
ropa;	 ->1	
ropa?	H->1	V->2	
ropaN	ä->1	
ropad	e->2	
ropag	a->3	e->1	r->1	
ropak	o->1	
ropam	i->1	
ropan	i->1	
ropap	a->166	
ropar	 ->3	å->1	
ropas	 ->48	
ropat	j->1	
ropav	a->3	
ropei	s->712	
ropet	 ->1	
ropol	 ->7	,->2	.->1	;->1	a->1	k->1	s->3	
ropor	t->9	
roppe	 ->1	n->1	
ropro	j->1	
ropå 	b->1	
ropé 	o->1	
ropée	r->9	
ror -	 ->1	
ror a	t->80	v->1	
ror d	e->6	ä->2	
ror e	g->1	
ror f	a->1	ö->1	
ror g	ö->1	
ror i	n->14	
ror j	a->23	u->1	
ror k	a->2	
ror m	a->1	e->2	i->1	y->1	
ror n	i->4	o->1	
ror o	c->7	
ror p	e->1	å->10	
ror s	a->1	o->3	å->1	
ror t	i->2	
ror u	p->1	t->1	
ror v	i->3	
ror ä	n->1	r->2	v->1	
ror ö	v->1	
ror, 	g->1	h->1	p->1	t->1	
ror.J	a->1	
ror.N	y->1	
ror.S	a->1	
ror.V	i->2	
ror?H	a->1	
rorda	 ->1	r->1	
rordn	a->5	i->42	
roren	a->19	i->9	
roris	m->2	t->8	
rorna	 ->6	
rorsa	k->6	
ros f	ö->1	
ros m	e->1	
ros o	c->1	
ros s	t->1	
rosat	s->1	
rosen	r->1	
roske	p->3	
rosmo	l->1	m->3	
rossa	r->1	
rosse	t->2	
rosst	ê->1	
rosta	t->2	
rostb	i->1	
rosti	t->1	
rot.J	a->1	
rota 	d->1	h->1	k->1	
rotad	e->2	
rotar	 ->2	
rotas	 ->5	
rotat	i->1	
rotek	t->4	
rotes	t->9	
rotfä	r->1	
rothe	r->1	
rotni	n->17	
rotok	o->26	
rots 	a->34	d->20	e->1	i->1	k->1	m->1	p->1	r->1	s->1	t->1	v->1	
rotsy	s->1	
rott 	a->1	b->1	i->2	m->4	o->2	p->2	s->2	
rott,	 ->9	
rott.	D->1	I->1	J->1	O->1	Ä->1	
rotta	t->2	
rotte	t->4	
rottm	å->1	
rotts	 ->1	b->3	f->1	l->17	m->2	o->2	r->1	
rotul	l->1	
rotur	i->1	
rouk 	a->1	
roup 	,->1	
roux-	a->1	
rov f	ö->4	
rov o	c->2	
rov p	å->9	
rov s	å->1	
rov",	 ->1	
rov, 	ä->1	
rov. 	D->1	
rov.D	e->1	
rovan	,->1	.->1	s->1	
rover	s->4	
rovet	 ->1	,->2	
rovic	 ->1	
rovin	s->3	
rovis	o->2	
rovka	r->1	
rovko	n->1	
rovsi	d->1	
rovsk	o->2	
rovst	e->1	
roväc	k->3	
rovär	d->15	
rpa a	n->1	
rpa b	e->1	
rpa d	e->1	
rpa h	e->1	
rpa k	o->1	
rpa t	e->1	
rpack	n->5	
rparl	a->1	
rpart	e->1	i->1	
rpas 	o->1	
rpas?	S->1	
rpass	a->1	
rpegn	a->1	
rpers	o->1	
rpet 	i->1	ä->1	
rplan	e->1	
rplik	t->21	
rpnin	g->1	
rpol-	f->1	
rpoli	t->20	
rpopu	l->1	
rpost	e->2	
rpres	i->1	
rpris	e->1	
rprog	r->3	
rproj	e->1	
rpt d	e->1	
rpt f	o->1	
rpta 	k->1	v->1	
rpus 	j->5	
rpå k	o->1	
rpå t	i->1	
rquio	l->1	
rr Al	a->1	
rr Ba	r->2	
rr Be	r->5	
rr Bo	u->1	w->2	
rr Co	x->3	
rr Ev	a->2	
rr Fr	u->1	
rr Go	l->1	
rr Gr	a->1	
rr Hä	n->2	
rr Jo	n->1	
rr Ki	n->4	
rr Ko	c->1	u->1	
rr La	n->1	
rr Mo	n->1	
rr No	g->1	
rr Pa	p->1	t->2	
rr Po	e->3	h->1	o->1	
rr Ra	p->1	
rr Sc	h->2	
rr Se	g->1	i->1	
rr Sp	e->1	
rr Wy	n->1	
rr al	l->1	
rr ba	r->1	
rr bl	i->1	
rr bö	j->1	
rr de	n->1	t->2	
rr då	 ->1	
rr el	l->2	
rr fi	c->1	
rr fo	r->1	
rr fö	r->6	
rr ge	n->1	
rr gö	m->1	
rr ha	r->6	
rr i 	k->1	
rr in	t->4	
rr ka	n->2	
rr ko	l->2	m->80	n->1	
rr le	d->15	
rr mi	n->2	
rr nä	r->1	
rr oc	k->1	
rr of	t->1	
rr or	d->5	
rr pa	r->3	
rr rå	d->12	
rr sa	m->1	
rr se	t->1	
rr st	e->1	
rr sä	g->1	
rr ta	l->319	
rr tj	ä->1	
rr va	n->3	
rr än	n->1	
rr är	 ->3	
rr äv	e->1	
rr åt	e->1	
rr öp	p->1	
rr, i	n->2	
rr, m	e->1	
rr, ä	n->1	
rr.Vi	 ->1	
rr?Vi	 ->1	
rra T	y->1	
rra d	e->2	
rra k	o->6	
rra m	å->2	
rra o	c->1	
rra p	r->2	
rra r	e->1	
rra s	i->1	
rra v	e->13	
rra å	r->19	
rrad 	a->1	
rrade	 ->1	
rrain	e->2	
rrand	 ->1	e->1	s->1	
rrang	e->6	
rrar 	P->1	m->1	o->1	p->4	t->2	v->1	
rrar!	 ->18	J->1	M->1	
rrar,	 ->16	
rrar.	V->1	
rrar;	 ->1	
rrarn	a->2	
rras 	y->1	
rras,	 ->1	
rrask	a->1	
rrat.	D->1	
rrati	o->2	
rrats	,->1	
rre -	 ->2	
rre a	m->1	n->5	r->1	
rre b	e->3	i->1	
rre d	e->3	
rre e	n->1	u->1	
rre f	r->2	ö->2	
rre h	a->1	ä->1	
rre i	 ->1	d->1	n->1	
rre j	ä->2	
rre k	a->1	r->1	
rre l	a->2	
rre m	e->3	å->1	
rre o	c->3	l->1	r->2	
rre p	l->1	r->2	å->1	
rre r	e->1	i->1	o->2	
rre s	a->1	i->1	j->1	k->1	n->1	o->1	t->2	ä->2	
rre t	y->1	
rre u	p->3	t->5	
rre v	a->1	i->4	o->1	
rre ä	n->3	
rre ö	p->6	
rre, 	i->1	
rrect	n->1	
rrefo	r->1	
rrege	r->3	
rregl	e->3	
rrekt	 ->13	,->2	.->6	;->1	a->5	
rren 	f->2	
rren,	 ->3	
rrens	 ->21	!->1	,->4	-->2	.->3	:->1	a->1	b->9	d->5	e->39	f->8	h->4	i->2	k->42	m->11	n->2	o->3	p->80	r->19	s->6	u->2	v->11	ä->2	
rrent	 ->1	e->1	
rrepa	r->1	
rrepr	e->2	
rrera	 ->4	d->1	
rres 	r->1	
rresp	o->1	
rrest	e->4	
rrey 	C->3	
rrez,	 ->1	
rrgån	g->1	
rrgår	 ->3	
rrido	r->2	
rrika	r->7	
rrike	 ->32	,->7	.->19	E->1	F->1	N->1	s->13	
rriki	s->49	
rring	 ->3	,->1	.->3	a->1	e->1	
rris 	(->1	
rrita	t->1	
rrite	r->3	
rrito	r->17	
rriär	e->3	p->1	
rroga	n->2	
rrong	e->1	
rror.	S->1	
rrori	s->10	
rrump	e->2	
rrupt	i->7	
rrvar	r->1	
rräde	r->1	
rrän 	m->2	å->2	
rrätt	a->1	e->1	
rråd 	(->1	
rråd,	 ->1	
rråde	n->1	t->12	
rrón 	i->1	t->1	v->1	
rrör 	s->2	t->1	u->1	
rröst	a->1	
rs 19	9->1	
rs 20	0->1	
rs EG	-->1	
rs EU	-->1	
rs al	l->1	
rs an	a->1	h->1	s->6	
rs ar	b->3	
rs at	t->1	
rs av	 ->18	
rs ba	k->1	
rs be	f->1	h->1	s->3	t->8	
rs bi	l->1	
rs br	u->1	
rs bu	d->3	
rs by	g->1	
rs de	l->5	n->1	
rs du	 ->1	
rs dö	d->2	
rs ef	t->1	
rs ek	o->3	
rs en	 ->3	d->1	l->1	
rs er	f->1	s->1	
rs et	t->2	
rs fl	a->4	e->1	
rs fo	r->1	
rs fr	a->3	i->1	ä->2	å->1	
rs fu	l->4	
rs fö	r->8	
rs gi	l->1	
rs go	d->1	
rs gr	u->1	
rs ha	d->2	n->2	r->3	
rs hj	ä->1	
rs hä	l->4	
rs i 	2->1	K->1	b->1	d->2	e->1	f->1	g->1	k->1	p->1	r->2	s->1	v->2	å->1	
rs in	k->2	s->1	t->4	
rs ju	d->1	
rs ka	n->3	p->1	
rs ko	m->5	
rs le	d->1	g->1	
rs li	b->2	v->1	
rs lä	r->1	
rs lö	p->1	
rs me	d->3	
rs mo	t->1	
rs må	l->1	n->1	s->2	
rs na	t->2	
rs ne	d->1	
rs ni	v->1	
rs oa	n->1	
rs oc	h->7	
rs of	f->1	
rs ok	u->1	
rs ol	ä->1	
rs or	g->1	
rs pa	r->5	t->1	
rs pl	a->1	
rs po	l->1	
rs pr	i->1	o->1	
rs på	 ->5	
rs ra	s->1	
rs re	g->1	s->1	
rs ro	l->1	
rs rä	k->1	t->3	
rs sa	m->1	
rs si	d->1	k->1	
rs sk	u->3	ö->1	
rs so	c->1	l->1	m->2	
rs st	a->1	r->1	ö->1	
rs sy	f->1	
rs sä	k->1	r->1	
rs så	r->1	v->1	
rs ta	c->1	
rs ti	d->4	l->2	
rs to	g->1	
rs tr	o->1	
rs ty	p->1	
rs un	d->1	
rs up	p->2	
rs ut	b->1	f->1	g->1	m->1	t->4	
rs va	l->2	
rs vä	g->1	
rs yr	k->1	
rs äg	a->1	
rs är	 ->2	
rs ås	i->1	
rs åt	e->1	
rs ök	a->1	
rs öp	p->1	
rs öv	e->3	
rs, L	u->1	
rs, a	t->2	
rs, e	n->1	
rs, f	ö->2	
rs, i	n->1	
rs, k	o->2	
rs, m	e->1	o->1	
rs, o	c->5	m->1	
rs, p	å->1	
rs, s	å->1	
rs, ä	v->1	
rs-bi	l->1	
rs. E	u->1	
rs..(	F->1	
rs.De	n->2	s->1	t->6	
rs.He	r->1	
rs.Ja	g->3	
rs.Me	n->1	
rs.Nu	 ->1	
rs.On	ö->1	
rs.Ty	v->1	
rs.Ut	f->1	
rs.Vi	 ->3	
rs.Vå	r->1	
rsaft	o->1	
rsail	l->1	
rsak 	t->1	
rsak.	E->1	N->1	
rsaka	 ->5	d->2	r->3	s->2	t->6	
rsake	n->4	r->13	
rsalm	e->1	
rsaml	a->1	i->12	
rsamm	a->7	
rsamt	 ->1	
rsana	l->1	
rsatt	a->4	s->1	
rsavg	r->1	
rsbef	r->2	
rsbel	o->1	
rsber	ä->1	
rsbes	l->1	
rsbri	s->1	
rsbud	g->1	
rsche	r->1	
rsdag	 ->5	.->3	
rse d	o->1	
rse f	r->1	ö->1	
rse k	o->1	
rse o	c->1	l->1	
rse s	a->1	
rse, 	l->1	
rse.D	e->1	
rse.V	a->1	
rseil	l->1	
rsekt	o->5	
rsel!	 ->1	
rsell	 ->2	a->1	
rsen 	-->1	f->1	h->1	n->1	o->1	p->1	
rsen,	 ->1	
rsena	 ->2	d->10	r->1	s->1	
rseni	n->13	
rser 	a->3	d->1	f->4	h->1	i->2	k->1	o->7	p->1	s->6	t->2	
rser,	 ->3	
rser.	.->1	D->2	H->1	I->1	V->2	
rsern	a->17	
rses 	m->1	
rsfri	h->43	
rsfrå	g->4	
rsful	l->4	
rsför	d->4	h->1	
rship	 ->1	
rsiel	l->9	
rsifi	e->2	
rsikt	 ->6	,->2	e->11	i->65	s->1	
rsinr	i->1	
rsion	 ->1	)->2	e->10	
rskal	a->2	i->2	
rskap	 ->13	,->5	.->4	a->2	e->5	s->4	
rskar	e->4	n->1	
rskas	.->1	
rskil	d->32	j->2	l->1	t->126	
rskin	g->2	
rskju	t->1	
rskni	n->35	
rskon	a->1	
rskot	t->2	
rskri	d->18	f->1	
rskro	t->1	v->1	
rskrä	c->4	
rskt 	m->1	
rskul	d->1	t->1	
rskäm	d->1	
rskän	n->1	s->2	
rskåd	l->6	
rskår	,->1	
rslag	 ->295	,->31	.->35	;->1	?->3	e->125	n->3	s->1	
rslan	d->1	
rslin	s->1	
rslun	t->1	
rsmak	t->1	
rsmed	e->1	
rsmin	i->1	
rsmän	n->1	
rsmål	.->1	
rsom 	D->1	E->3	F->2	O->1	T->1	a->6	b->2	d->85	e->2	f->6	h->5	i->3	j->13	k->2	m->12	n->3	o->1	p->4	r->2	s->6	t->4	u->1	v->23	å->1	
rsom,	 ->1	
rsomr	å->7	
rson 	a->1	h->2	i->2	s->1	
rson,	 ->1	
rsona	l->23	n->1	
rsone	l->2	n->1	r->40	
rsoni	n->4	
rsonl	i->34	
rsons	 ->1	
rsord	n->1	
rsot 	s->1	
rspeg	l->3	
rspek	t->17	
rsper	i->3	
rspol	i->4	
rspor	t->1	
rspos	t->1	
rspro	g->1	
rspru	n->19	
rspår	n->1	
rsrap	p->2	
rsski	f->2	
rsslö	s->1	
rst a	l->1	v->8	
rst c	a->1	
rst d	å->3	
rst e	f->3	x->1	
rst f	å->1	
rst g	e->1	j->1	
rst h	a->2	
rst i	 ->4	n->1	
rst j	u->1	
rst k	a->1	r->1	
rst m	o->1	å->3	
rst n	o->1	ä->1	å->1	
rst o	c->22	m->1	
rst p	r->1	
rst r	e->1	i->1	ä->1	
rst s	e->1	k->6	l->1	t->3	v->1	ä->1	
rst t	a->3	
rst u	t->1	
rst v	a->1	i->12	ä->1	
rst.M	e->1	i->1	
rsta 	a->8	b->19	c->1	d->14	e->3	f->12	g->29	h->26	i->5	k->6	l->2	m->14	n->3	o->3	p->10	r->19	s->15	t->12	u->5	v->11	ä->10	å->1	ö->1	
rsta,	 ->10	
rsta:	 ->5	
rsta;	 ->2	
rstab	e->1	
rstad	 ->1	
rstag	a->1	
rstai	n->22	
rstak	l->1	
rstat	.->1	e->1	l->3	
rste 	a->1	
rstid	e->2	
rstig	e->1	l->4	
rstil	l->1	
rstkl	a->1	
rstod	 ->3	
rstol	e->1	
rstre	c->1	
rstry	k->27	
rsträ	v->12	
rströ	k->2	
rstäd	e->2	
rstäl	l->41	
rstär	k->29	
rstå 	a->8	d->2	f->2	h->2	n->1	o->1	v->4	
rstå,	 ->1	
rstå.	F->1	J->1	
rståd	d->2	
rståe	l->13	n->1	
rstån	d->9	
rstår	 ->40	,->1	.->1	
rstås	 ->4	
rståt	t->10	
rstöd	 ->2	e->2	j->5	
rstör	 ->3	a->5	d->3	e->5	i->2	s->1	t->2	
rsumb	a->1	
rsumm	a->2	e->6	
rsund	i->3	
rsvag	a->20	n->1	
rsvar	,->1	.->2	a->25	e->4	s->9	
rsvin	n->15	
rsvun	n->4	
rsväm	m->3	n->4	
rsvår	a->2	
rsydd	a->1	
rsyn 	a->1	
rsynt	,->1	
rsäkr	a->20	i->24	
rsäkt	 ->7	.->1	a->4	e->3	
rsälj	a->2	n->3	
rsämr	a->10	
rsänd	r->1	
rsänk	t->1	
rsätt	a->10	e->3	l->1	n->20	s->1	
rsågs	 ->1	
rsåte	 ->1	
rsök 	a->4	s->1	
rsök,	 ->2	
rsöka	 ->36	,->1	s->4	
rsöke	n->1	r->16	t->3	
rsökn	i->23	
rsökt	 ->13	e->5	
rsörj	n->4	
rsöve	r->1	
rt - 	d->1	m->1	n->1	o->2	ä->1	
rt Ca	m->1	
rt Du	i->1	
rt EG	-->1	
rt Eu	r->4	
rt FP	Ö->1	
rt Go	e->1	
rt ag	e->2	
rt al	l->1	
rt an	s->8	t->7	v->1	
rt ar	b->9	v->1	
rt at	t->89	
rt av	 ->28	g->1	s->3	t->1	
rt ba	r->1	
rt be	k->2	s->2	t->8	
rt bi	d->2	s->1	
rt bl	i->1	
rt bo	r->1	
rt br	e->1	
rt bu	d->1	
rt bä	t->2	
rt bö	r->2	
rt de	b->1	n->5	s->1	t->16	
rt dj	u->1	
rt dr	a->2	
rt dy	r->1	
rt dä	r->1	
rt eg	e->5	
rt ek	o->4	
rt el	l->1	
rt em	o->2	
rt en	 ->12	g->1	
rt er	 ->2	k->1	
rt et	t->10	
rt eu	r->3	
rt ex	a->1	
rt fa	l->1	s->4	t->1	
rt fi	n->3	
rt fr	a->3	å->8	
rt få	 ->1	r->1	
rt fö	l->2	r->48	
rt ge	 ->1	m->2	n->5	
rt go	d->1	
rt gr	e->1	ä->2	
rt gå	 ->2	
rt ha	n->3	r->2	
rt he	l->1	
rt hi	t->1	
rt ho	p->1	r->1	s->1	
rt hu	r->3	
rt hä	r->1	
rt hå	l->1	
rt i 	B->1	D->1	d->3	e->2	f->4	p->1	s->1	
rt if	r->1	
rt in	c->1	f->1	i->1	l->1	n->1	o->1	r->1	s->1	t->14	v->1	
rt ka	n->2	
rt kl	a->2	
rt kn	y->1	
rt ko	m->8	n->1	
rt kr	a->1	i->1	o->1	ä->1	
rt ku	l->2	n->1	
rt kä	r->1	
rt la	n->3	
rt li	k->1	
rt lo	b->1	
rt ly	c->1	
rt lä	g->1	m->1	r->1	
rt lö	f->1	p->1	
rt ma	n->1	r->1	t->2	
rt me	d->20	
rt mo	t->2	
rt my	c->2	
rt må	l->4	n->2	s->1	t->1	
rt mö	t->1	
rt ne	d->1	
rt nu	v->1	
rt ny	a->1	s->1	
rt nä	m->1	r->1	
rt nå	g->8	
rt oc	h->40	k->1	
rt ol	i->1	
rt om	 ->13	.->1	r->1	
rt or	d->6	
rt os	s->2	
rt pa	k->1	r->13	
rt pe	r->2	
rt po	l->2	s->2	
rt pr	i->1	o->5	
rt på	 ->8	m->1	
rt re	d->1	f->1	g->1	k->1	l->1	s->1	
rt ri	k->1	
rt rä	t->1	
rt sa	g->4	m->8	
rt se	r->1	t->4	
rt si	g->4	k->5	t->2	
rt sk	a->4	u->3	
rt sl	å->1	
rt so	m->24	
rt sp	e->1	r->1	
rt st	e->2	o->2	ä->2	ö->8	
rt sv	a->6	å->2	
rt sy	s->3	
rt sä	g->3	t->7	
rt så	 ->4	
rt ta	 ->1	c->6	l->2	s->1	
rt te	c->1	k->1	
rt ti	d->2	l->2	
rt to	l->1	p->1	
rt tr	ä->1	
rt ty	s->1	
rt un	d->5	
rt up	p->2	
rt ut	b->1	f->2	g->1	m->1	r->1	s->11	t->4	
rt va	d->1	l->1	
rt ve	r->1	t->2	
rt vi	 ->1	d->1	k->1	l->3	n->1	s->1	
rt vä	l->1	n->1	
rt vå	r->1	
rt yt	t->2	
rt Ös	t->1	
rt äm	b->1	
rt än	d->2	
rt är	 ->6	
rt åt	a->1	
rt ög	o->1	
rt öv	e->2	
rt!He	r->1	
rt!Ja	g->1	
rt) t	ä->1	
rt, a	t->1	
rt, b	ö->2	
rt, c	i->1	
rt, d	e->1	å->1	
rt, e	f->3	n->1	
rt, g	å->2	
rt, h	a->2	e->3	å->1	
rt, i	 ->1	
rt, k	a->1	u->1	
rt, l	ä->1	
rt, m	e->6	å->1	
rt, n	ä->1	
rt, o	c->6	
rt, p	å->1	
rt, s	o->2	å->1	
rt, t	a->1	o->1	r->1	
rt, v	i->4	
rt, ä	n->1	r->1	
rt- o	c->1	
rt-st	a->2	
rt. 7	)->1	
rt. I	n->1	
rt.Ar	t->1	
rt.De	n->4	s->1	t->2	
rt.Di	r->1	
rt.Då	 ->1	
rt.En	 ->1	
rt.Fr	u->1	
rt.Fö	r->1	
rt.Hä	r->1	
rt.I 	d->1	s->1	
rt.Ja	g->6	
rt.Ju	s->1	
rt.Ko	m->2	n->1	
rt.Lå	t->1	
rt.Me	n->2	
rt.Ni	 ->1	
rt.Oc	h->1	
rt.Ri	k->1	
rt.Sa	m->1	
rt.Sl	u->1	
rt.St	ö->1	
rt.Ut	b->1	
rt.Va	d->1	
rt.Vi	 ->5	l->1	
rt.Äv	e->1	
rt: E	f->1	
rt: e	t->1	
rt?Ja	g->1	
rtNäs	t->1	
rta a	l->1	
rta d	e->1	
rta e	g->1	
rta f	r->4	
rta k	l->1	
rta m	e->1	
rta o	c->1	m->1	r->1	
rta p	å->1	
rta r	ö->1	
rta s	o->1	
rta t	a->1	
rta u	t->1	
rta ä	r->1	
rtabl	a->1	
rtad 	f->1	s->1	
rtade	 ->2	s->1	
rtag,	 ->1	
rtaga	n->8	
rtagn	a->1	
rtal 	b->1	f->1	t->1	
rtala	 ->1	
rtale	t->4	
rtame	-->1	
rtand	e->1	
rtank	e->3	
rtann	a->3	
rtans	 ->2	
rtar 	a->1	o->1	
rtar,	 ->1	
rtar.	J->1	V->1	
rtas 	i->1	m->1	u->1	
rtast	e->1	
rtat 	-->1	a->2	d->1	g->1	o->1	p->1	s->2	t->1	
rtat,	 ->1	
rtat.	 ->1	D->1	
rtat:	 ->1	
rtats	 ->2	
rtbes	t->2	
rtbil	d->1	
rtdir	e->1	
rteck	e->4	n->20	
rtell	-->3	a->1	b->2	e->1	f->3	m->1	r->4	
rteme	n->9	
rten 	1->1	a->8	b->1	f->4	g->1	h->1	i->4	k->2	l->1	o->14	s->2	u->1	v->2	å->1	
rten,	 ->3	
rten.	D->1	E->1	I->1	O->1	S->1	
rten:	 ->1	
rtend	a->1	
rtens	 ->3	
rter 	(->1	-->1	a->5	d->1	e->1	f->3	i->2	k->2	m->1	o->4	p->4	r->1	s->6	t->4	u->1	
rter,	 ->7	
rter.	D->4	E->1	I->1	M->2	P->1	S->1	V->2	
rtera	 ->3	d->6	r->2	s->8	t->3	
rteri	n->1	
rtern	a->30	
rtet 	f->13	i->1	s->1	
rtet.	J->1	
rtets	 ->3	
rtext	 ->3	
rtfal	l->6	
rtfar	a->89	
rtfat	t->2	
rtfed	e->1	
rtfrå	g->1	
rtför	b->1	
rtgru	p->4	
rtgå.	D->1	N->1	
rtgåe	n->3	
rthet	s->1	
rthu 	o->1	
rthy 	o->1	
rti a	n->1	
rti d	e->1	
rti f	r->1	ö->1	
rti h	a->1	e->1	
rti i	 ->2	n->2	
rti k	o->1	
rti m	e->1	
rti p	å->1	
rti s	n->1	o->6	
rti t	i->2	
rti å	t->1	
rti, 	M->1	d->1	k->1	l->1	p->1	s->1	ä->1	
rti..	.->1	
rti.D	e->1	
rti.H	a->1	
rti.K	a->1	
rtid 	E->1	a->14	b->2	d->3	e->6	f->3	h->1	i->10	j->1	k->1	l->1	m->5	n->1	o->4	s->5	t->2	u->1	v->1	ä->3	å->1	
rtid,	 ->3	
rtids	p->6	
rtiel	l->2	
rtier	 ->5	,->1	n->4	
rtiet	 ->6	)->4	,->4	s->16	
rtifi	c->2	e->2	k->4	
rtigh	e->1	
rtiin	t->1	
rtika	l->3	
rtike	l->95	
rtikl	a->15	
rtikr	a->1	
rtile	d->1	
rtill	 ->2	v->1	
rtine	z->1	
rtino	t->1	
rtio 	g->1	å->2	
rtion	 ->3	a->1	d->1	e->5	
rtios	j->1	
rtipr	o->2	
rtis 	r->1	u->1	
rtis,	 ->1	
rtis.	D->1	
rtisk	 ->1	t->2	
rtisp	l->1	
rtjus	t->1	
rtjän	a->13	s->4	t->3	
rtkom	m->17	
rtkos	t->2	
rtlev	n->1	
rtlig	t->7	
rtläg	g->1	
rtmar	k->1	
rtmon	n->1	
rtner	 ->7	.->1	?->1	n->1	s->18	
rtnin	g->2	
rtnät	 ->1	
rtog 	m->1	
rtom 	a->6	b->1	f->2	h->1	i->2	s->2	t->1	
rtom!	T->1	
rtom,	 ->3	
rtom.	V->1	
rtomr	å->3	
rton 	a->1	m->6	s->1	
rtond	e->1	
rtone	r->1	
rtonh	u->1	
rtpla	t->1	
rtpri	o->1	
rtpro	b->1	
rtrak	t->1	
rtram	p->1	
rtran	s->1	
rtrap	p->1	
rtrar	 ->1	
rtreg	e->1	
rtroe	n->56	
rtrog	e->1	
rtros	 ->2	
rtrot	t->1	
rtryc	k->2	
rträd	d->1	e->5	
rträf	f->3	
rträn	g->1	
rtröt	t->1	
rts "	B->1	
rts a	n->2	v->11	
rts c	o->1	
rts d	i->3	
rts e	l->1	n->1	
rts f	a->1	r->2	ö->3	
rts h	i->1	ä->3	
rts i	 ->6	
rts m	e->2	
rts n	å->1	
rts o	c->4	m->2	
rts p	å->2	
rts s	e->1	
rts t	i->1	
rts u	t->1	
rts v	a->1	e->1	
rts, 	b->2	s->1	u->1	v->1	å->1	
rts.D	e->1	
rts.J	a->2	
rts.S	l->1	
rts.T	a->1	
rts.V	i->1	
rtsam	m->1	
rtsat	t->12	
rtse 	f->4	
rtser	 ->1	
rtset	t->1	
rtsif	f->1	
rtsik	t->4	
rtsin	s->1	
rtskr	i->1	
rtsme	d->1	
rtsmy	n->1	
rtsor	g->2	
rtsse	k->3	
rtsäk	e->7	
rtsät	t->82	
rtuga	l->26	
rtugi	s->70	
rtugu	e->1	
rtuni	s->2	
rtuse	n->3	
rtuts	k->2	
rtvin	 ->1	
rtviv	l->1	
rtydl	i->3	
rtyg 	d->1	f->2	i->4	m->3	o->1	s->14	u->3	
rtyg)	,->1	
rtyg,	 ->3	
rtyg.	E->1	F->1	V->2	
rtyg;	 ->1	
rtyga	 ->7	d->21	n->5	r->1	
rtyge	l->4	n->13	t->7	
rtygs	b->1	i->1	s->8	t->1	ä->1	
rtyre	n->1	
rtz o	c->1	
rtz s	o->1	
rtz, 	p->1	
rtäck	t->1	
rtänk	s->1	t->1	
ru Ah	e->2	
ru An	g->1	
ru Be	r->1	
ru Fr	a->1	
ru Ly	n->1	
ru Mc	N->1	
ru Pe	i->1	
ru Pl	o->1	
ru Re	d->3	
ru Sc	h->3	
ru Su	d->1	
ru Th	e->1	
ru Wa	l->1	
ru ko	m->46	
ru le	d->2	
ru ta	l->83	
ru, s	i->1	
ruari	 ->7	!->1	,->7	.->1	
rubba	 ->1	r->1	s->1	
rubri	k->2	
rucki	t->1	
ruckn	e->1	
ruera	 ->3	d->1	t->1	
ruhe 	o->1	
ruhe,	 ->1	
ruine	r->1	
ruk a	v->1	
ruk m	e->1	
ruk o	c->5	
ruk p	å->1	
ruk s	o->1	
ruk!A	n->1	
ruk, 	d->3	e->1	i->1	m->1	t->2	v->1	
rukad	e->2	
rukar	:->1	e->8	n->5	
rukas	 ->1	
ruken	.->1	
ruket	 ->13	,->2	.->1	;->2	s->1	
rukit	s->1	
rukni	n->1	
rukse	k->1	
ruksf	o->1	r->1	
ruksl	o->1	
rukso	m->2	
ruksp	o->6	r->3	
ruksr	e->2	
rukss	e->5	y->1	
rukt 	a->1	
rukt.	H->1	
rukta	n->7	r->3	t->1	
ruktb	a->2	
rukte	n->1	
rukti	o->18	v->12	
ruktu	r->153	
ruktö	r->3	
rulla	r->3	
rulls	t->3	
rum e	n->1	
rum f	i->1	ö->6	
rum h	a->1	ä->1	
rum i	 ->16	n->2	
rum m	e->1	
rum o	c->1	m->3	
rum p	å->3	
rum u	n->1	t->1	
rum y	t->1	
rum å	t->1	
rum!M	e->1	
rum, 	d->2	o->1	u->1	v->1	
rum. 	D->1	
rum.D	e->1	
rum.M	e->1	
rum.O	M->1	
rumen	t->52	
rumet	 ->3	
rumpe	r->2	
runa 	p->1	
rund 	a->81	f->16	i->3	o->1	s->1	t->1	u->1	v->1	ä->2	
rund,	 ->1	
rund.	P->1	
rund?	 ->1	
runda	 ->5	.->1	d->8	n->3	r->2	s->6	t->5	
rundb	u->1	
runde	n->32	r->6	
rundf	ö->4	
rundk	u->1	
rundl	i->16	ä->74	
rundo	r->1	
rundp	e->1	r->1	
rundr	e->2	
runds	a->1	t->1	
rundt	e->1	
rundv	a->25	
rung 	o->2	
rung.	I->1	O->1	
runge	t->2	
rungl	i->12	
rungs	l->1	
runkn	a->3	
runo 	L->1	
runt 	o->3	t->1	
runt.	D->1	
runta	 ->2	r->1	
runto	m->1	
runtp	r->1	
rupp 	(->2	a->9	b->2	e->1	f->3	h->4	i->2	k->4	l->2	m->1	n->1	o->2	p->3	r->2	s->6	t->3	u->3	v->4	ä->2	
rupp,	 ->9	
rupp.	F->1	M->1	
rupp?	H->1	
ruppb	y->12	
ruppe	n->63	r->57	
ruppk	o->1	
ruppl	i->1	
ruppo	r->1	
ruppr	e->1	ä->6	
rupps	 ->4	t->3	
ruppt	a->8	i->1	o->2	ä->1	
ruppu	n->1	
ruppv	i->1	
rupti	o->7	
rusa 	v->1	
rusal	e->2	
rusar	 ->2	
rusta	 ->1	d->2	
rustb	e->1	
ruste	n->1	r->3	
rustn	i->5	
rustr	a->1	e->1	
rut a	t->1	
rut o	c->1	
rut.D	e->1	
rutal	.->1	a->1	
rutbe	s->1	
rutbi	l->2	
rutea	u->3	
ruten	 ->1	
rutet	 ->1	
rutgi	f->1	
rutin	e->7	m->1	
rutit	 ->1	s->1	
rutom	 ->15	
rutsa	t->1	
rutse	 ->4	.->1	s->1	t->2	
rutsk	o->1	
rutsä	g->2	t->52	
rutte	n->1	
ruttn	a->2	
rutto	n->1	
rutva	r->2	
rutve	c->2	
rutöv	e->1	
ruva 	i->1	
ruvid	a->15	
rv få	r->1	
rv oc	h->2	
rv, a	t->1	
rv, e	n->1	
rv, s	o->1	
rv."D	e->1	
rv.Ba	r->1	
rv.En	 ->1	
rva d	e->1	
rva f	ö->1	
rva n	å->1	
rva o	c->1	
rva p	å->1	
rva r	e->1	
rvade	 ->1	
rvaka	 ->7	.->1	r->3	s->2	t->1	
rvakn	i->11	
rval 	a->2	e->1	
rvale	t->1	
rvals	k->1	
rvalt	a->2	n->47	
rvand	l->4	
rvans	k->2	
rvara	 ->3	n->39	
rvare	 ->1	
rvarn	i->1	
rvaro	 ->2	n->2	
rvarr	 ->1	
rvat 	d->1	
rvati	o->2	v->7	
rvats	 ->1	
rvatt	e->9	n->8	
rvatö	r->1	
rvbri	n->1	
rveck	a->1	
rven 	f->1	s->1	v->1	
rven.	D->1	T->2	
rvene	r->2	
rvent	i->5	
rver 	f->1	i->2	
rvera	d->1	t->1	
rverk	a->1	l->22	
rvet 	a->1	h->1	i->1	
rvet,	 ->1	
rvete	n->1	
rvhet	 ->1	
rvice	.->4	k->2	n->1	
rvid 	a->1	d->1	k->1	m->2	o->1	p->1	s->1	
rvidl	a->1	
rvinn	a->21	e->4	i->47	s->2	
rvirr	a->4	i->8	
rvis 	f->1	
rvisa	 ->1	d->1	
rviss	a->2	o->6	
rvju 	m->1	s->1	
rvjua	d->1	
rvlig	.->1	h->1	
rvrid	n->1	
rvrän	g->1	
rvsar	b->3	
rvsin	d->1	
rvsst	ö->2	
rvt p	r->2	
rvtru	p->1	
rvunn	a->1	e->1	i->1	
rväg 	a->2	f->1	h->1	i->1	
rväg,	 ->4	
rväg.	O->1	V->1	
rväga	 ->16	,->1	n->8	
rvägd	a->1	
rväge	r->7	
rvägr	a->3	
rvägt	 ->2	
rväld	i->3	
rvänd	a->2	e->1	
rvänt	a->22	n->7	
rvärd	e->5	
rvärl	d->2	
rvärr	a->4	
rvärt	.->1	
rvärv	a->4	s->3	
rvåna	 ->1	d->3	n->1	s->1	
rwell	s->1	
ry Fo	r->1	
ry oc	h->1	
ry, H	a->1	
ry.De	 ->1	
ryck 	a->7	e->1	f->10	i->2	k->1	m->1	p->1	s->1	
ryck,	 ->2	
ryck.	D->1	
rycka	 ->22	n->1	
ryckb	ä->1	
rycke	r->7	t->12	
ryckl	i->13	
ryckn	i->5	
rycks	 ->3	
ryckt	 ->4	e->9	s->1	
ryfta	 ->1	
rygga	 ->4	d->1	n->1	
rygge	n->3	
ryggh	e->6	
ryggr	a->1	
rygt 	4->1	e->1	t->1	
ryk.H	e->1	
ryka 	-->1	P->1	a->11	d->5	e->1	f->1	m->1	s->1	v->1	
ryka,	 ->2	
rykas	 ->4	
ryker	 ->2	
ryks 	o->1	v->1	
rykta	d->1	
ryktb	a->1	
rykte	 ->4	,->1	.->1	n->1	
rymd 	t->1	
rymde	n->1	
rymma	 ->1	
rymme	 ->10	,->1	
ryms 	i->1	
rymt 	a->1	
ryost	a->1	
ryphå	l->3	
ryps.	M->1	
rypto	g->2	
ryr e	r->1	
ryr j	a->1	
rys o	r->1	
rysa 	s->1	v->1	
rysk 	e->1	
ryska	 ->1	
rysni	n->1	
ryssa	 ->1	r->1	
rysse	l->19	
ryta 	d->2	k->1	m->3	
rytan	d->1	
rytas	 ->1	
rytel	s->2	
ryter	 ->6	i->1	
rytni	n->2	
rytte	r->2	
rzwal	d->1	
rä ut	g->1	
rä öv	e->1	
räck 	s->1	
räcka	 ->10	,->1	n->2	
räcke	n->1	r->21	
räckh	e->1	
räckl	i->77	
räckn	i->31	
räcks	 ->1	c->1	
räckt	 ->2	e->1	
räckv	i->3	
räd b	e->1	
räd f	ä->1	
räd h	a->2	
räd u	p->1	
räd, 	o->1	
räd.D	e->1	
räda 	E->1	e->1	i->6	s->1	u->1	
räda,	 ->1	
rädan	d->10	
rädar	e->47	n->10	
rädd 	a->2	f->3	
rädd,	 ->1	
rädda	 ->9	d->3	r->1	t->1	
rädde	 ->7	
räddn	i->4	
räde 	-->1	a->1	e->1	f->1	h->1	i->1	k->1	m->1	o->3	t->4	
räde.	H->1	J->2	
rädeH	e->1	
rädeP	r->1	
rädel	s->5	
räden	 ->3	a->1	
räder	 ->14	,->1	i->1	
rädes	p->7	v->2	
rädet	 ->10	,->1	.->1	
räds 	a->1	i->1	
rädsl	a->9	
räffa	 ->5	,->2	.->1	d->6	n->41	r->49	s->2	t->9	
räffl	i->2	
räfta	 ->11	,->1	d->3	r->3	s->5	t->6	
räfte	l->1	
rägar	n->1	
räger	i->36	
rägla	d->4	s->1	
rägli	g->1	
räken	s->9	
räkna	 ->8	d->1	r->21	s->4	t->5	
räkne	e->1	l->1	
räkni	n->14	
räkta	 ->1	
räkts	 ->1	
räl g	ä->1	
räl i	n->1	
räl, 	m->1	
rämbe	t->1	
rämd 	h->1	
rämel	s->1	
rämja	 ->36	.->1	n->17	r->6	s->1	t->1	
rämli	g->1	n->34	
rämma	n->3	
rämme	r->2	
rämst	 ->35	.->1	a->12	
rän m	a->1	y->1	
rän n	a->1	
rän s	t->1	
rän å	r->2	
räna 	r->1	s->2	
rända	 ->2	
rände	r->4	
rändr	a->27	i->46	
räng 	k->2	o->1	å->1	
ränga	 ->11	,->1	n->1	r->3	s->2	
rängd	 ->1	e->1	
ränge	r->5	
rängn	i->35	
rängt	 ->5	
ränin	g->1	
ränit	e->12	
ränka	 ->2	
ränkb	a->1	
ränke	r->5	
ränkn	i->13	
ränks	 ->3	
ränkt	a->5	s->2	
ränna	 ->2	s->1	
ränni	n->2	
räns 	v->2	
ränsa	 ->12	,->1	d->27	n->3	r->5	s->5	t->9	
ränse	n->4	r->30	
ränsf	r->2	
ränsk	o->7	
ränsl	e->7	
ränsn	i->12	
ränso	m->1	
ränsp	r->1	
ränsv	ä->1	
ränsö	v->12	
ränta	 ->1	
räpni	n->1	
räpro	d->1	
rär o	c->1	
rärt 	F->1	
räsch	 ->1	e->1	
räsk.	H->1	
rätas	 ->1	
rätor	 ->1	
rätt 	(->2	-->1	a->21	e->2	f->6	h->3	i->12	k->3	m->3	n->4	o->12	p->2	r->6	s->10	t->18	u->1	v->4	ä->1	ö->1	
rätt,	 ->10	
rätt.	 ->1	F->1	H->1	J->1	M->2	V->1	
rätt?	O->1	S->1	
rätta	 ->60	,->2	.->1	d->7	n->19	r->5	s->11	t->9	
rätte	g->1	l->4	n->84	r->1	
rättf	r->1	ä->7	
rätth	å->9	
rätti	g->122	
rättm	ä->1	
rättn	i->2	
rätts	a->4	f->1	h->2	i->2	k->9	l->118	o->6	p->2	r->1	s->52	t->3	v->4	
rättv	i->72	
rättä	n->1	
räva 	4->1	a->7	d->3	e->9	f->3	i->1	j->1	k->1	m->2	t->2	å->2	ö->1	
rävad	e->4	
rävan	 ->8	.->1	d->7	s->1	
rävar	 ->4	
rävas	 ->7	,->1	.->1	
rävat	 ->1	
rävde	 ->1	,->1	s->2	
räver	 ->43	.->2	
rävig	t->1	
rävs 	a->2	b->1	d->11	e->12	f->8	h->1	i->2	k->1	m->2	o->1	p->1	r->1	s->4	u->1	v->3	ä->1	
rävs,	 ->3	
rävt 	e->1	
rävts	 ->1	
rå so	m->1	
rå va	r->1	
rå är	 ->1	
råd (	a->1	
råd -	 ->1	
råd a	n->1	
råd b	e->1	
råd f	r->2	ö->1	
råd i	 ->1	
råd n	ä->1	
råd o	c->2	m->3	
råd s	o->3	
råd, 	b->1	m->1	o->2	
råd.D	e->1	
råd.J	a->1	
råd.K	a->1	
råd.L	å->1	
råd.M	e->1	
råd?Ä	r->1	
råda 	b->2	e->4	m->2	n->1	
rådan	d->4	
rådar	 ->1	.->1	n->1	
rådde	 ->1	
råde 	-->1	a->4	d->4	e->2	f->7	h->2	i->3	k->3	m->9	n->1	o->7	s->6	v->2	ä->5	å->1	
råde,	 ->14	
råde.	 ->1	D->4	F->4	I->2	J->3	M->4	O->2	P->1	T->1	V->1	
råde:	 ->1	
råde;	 ->1	
råde?	D->1	
råden	 ->61	)->1	,->10	.->20	:->2	;->1	?->2	a->36	s->1	
råder	 ->24	
rådet	 ->198	)->1	,->45	.->52	:->1	?->4	s->95	
rådfr	å->6	
rådgi	v->26	
rådgö	r->1	
rådsb	e->1	
rådsk	a->20	
rådsl	a->3	
rådsm	e->1	i->1	ö->1	
rådso	r->19	
rådsr	ä->1	
rådst	o->1	
råer,	 ->1	
rået.	D->1	
råga 	-->1	a->7	b->2	e->2	f->7	g->4	h->9	i->6	j->1	k->7	m->7	n->27	o->82	p->3	r->4	s->45	t->4	v->5	ä->9	
råga!	F->1	
råga,	 ->24	
råga.	 ->1	-->1	A->1	D->8	E->2	F->2	H->3	I->2	J->8	M->2	N->1	S->1	T->1	U->1	V->5	Ä->1	
råga:	 ->7	
råga?	.->1	
rågad	e->8	
rågan	 ->168	,->11	.->16	:->5	;->1	?->1	d->1	
rågar	 ->19	.->1	
rågas	a->1	ä->19	
rågat	 ->3	a->1	s->2	
rågav	a->1	
rågek	o->1	
råges	t->10	
råget	e->2	
rågni	n->8	
rågor	 ->176	)->1	,->37	.->28	:->4	;->1	n->28	
råk f	ö->1	
råk p	å->3	
råk t	i->1	
råk. 	D->1	
råka 	e->1	
råkar	 ->5	e->3	n->1	
råket	 ->2	.->2	
råkig	t->3	
råkli	g->3	
råkom	r->2	
råkra	t->30	
råkta	g->1	
råldr	a->3	
rålka	s->1	
rålni	n->3	
rålsk	y->1	
rån (	H->21	
rån -	 ->1	
rån 1	0->1	5->1	9->5	
rån 2	8->1	
rån 3	,->1	
rån 5	 ->2	0->1	
rån 8	9->1	
rån 9	5->1	
rån A	f->1	l->2	m->4	t->2	u->1	
rån B	S->1	a->1	o->1	r->2	
rån C	E->2	a->1	
rån D	a->1	e->1	
rån E	G->2	U->1	r->2	u->24	
rån F	M->1	l->3	r->1	ö->1	
rån G	U->1	a->1	o->1	ö->1	
rån H	e->2	
rån I	R->1	n->3	s->1	
rån J	a->1	
rån K	o->1	y->2	ö->2	
rån L	a->1	i->1	o->1	
rån M	a->1	
rån N	a->3	
rån O	S->1	
rån P	P->2	S->1	a->1	o->3	
rån R	o->1	
rån S	a->3	h->1	y->2	
rån T	a->4	e->1	y->1	
rån U	N->1	S->1	
rån V	e->1	
rån W	i->1	u->1	
rån a	l->4	n->3	t->26	v->2	
rån b	e->1	i->3	o->2	u->2	ö->5	
rån d	a->3	e->86	i->4	o->1	
rån e	n->19	r->3	t->17	u->1	x->3	
rån f	a->2	l->2	r->2	ö->27	
rån g	e->4	
rån h	a->3	e->1	ö->2	
rån i	 ->1	
rån j	u->4	
rån k	a->3	o->34	
rån l	a->1	e->3	ä->4	
rån m	a->4	e->6	i->8	o->1	å->2	
rån n	a->1	y->2	å->3	
rån o	b->1	c->11	f->1	l->4	p->1	r->2	s->2	
rån p	a->13	e->1	r->4	
rån r	a->1	e->3	å->13	
rån s	a->2	e->1	i->8	k->3	o->2	t->4	y->1	ä->3	ö->1	
rån t	.->1	i->5	o->2	r->16	u->1	
rån u	n->2	t->20	
rån v	a->2	e->1	i->5	ä->1	å->10	
rån Ö	s->1	
rån ä	r->1	
rån å	r->1	
rån ö	v->4	
rån, 	d->1	n->1	o->1	
rån.D	ä->1	
rån.Ä	n->1	
rång 	i->1	
rång,	 ->2	
rånge	l->1	
rångl	i->1	
rångm	å->1	
rångå	r->1	
rånko	m->3	
rånta	r->1	s->1	
rånto	g->1	
rånva	r->8	
rånvä	n->1	
råolj	a->1	
råpsl	a->1	
rårig	a->6	t->6	
rås f	ö->2	
råt k	o->1	
råtgä	r->1	
råtto	r->1	
råzon	 ->1	
rébet	o->1	
référ	e->1	
rêts 	(->1	
rínci	p->1	
rón C	r->2	
rón i	 ->1	
rón t	i->1	
rón v	i->1	
röd.-	 ->1	
röd.D	e->1	ä->1	
röda 	t->2	
rödan	d->3	
rödel	s->2	
röder	 ->1	
rödgr	ö->1	
rödor	.->1	
röghe	t->1	
röja 	d->3	k->1	t->1	
röja.	V->1	
röjar	e->1	
röjas	.->1	
röjde	 ->1	
röjer	 ->3	
röjor	.->1	
röjsm	å->2	
röjts	,->1	
rök b	e->1	
rök, 	d->1	
röks,	 ->1	
röm a	v->2	
röm b	e->1	
röm i	n->1	
röm, 	s->1	
röm: 	N->1	
römma	 ->1	r->3	
römme	n->4	
römni	n->6	
römt 	W->1	
römvä	r->1	
rön v	ä->2	
röna 	e->1	f->1	g->2	h->1	i->1	m->1	n->1	o->1	p->1	s->2	
röna/	E->1	
rönar	e->1	
rönas	 ->2	
rönbo	k->1	
rönit	z->1	
rönt 	l->1	
rör E	u->1	
rör P	o->1	
rör a	l->1	n->1	s->1	
rör b	e->1	
rör d	e->6	
rör f	l->1	r->2	ö->3	
rör i	 ->1	
rör j	u->1	
rör k	ä->1	
rör o	c->2	s->1	
rör p	a->1	r->1	å->1	
rör s	a->1	i->13	o->1	t->2	
rör t	.->1	i->1	
rör u	n->1	p->1	r->1	
rör v	i->1	
röra 	s->2	v->1	
röran	d->24	
röras	 ->2	
rörd 	a->1	o->1	
rörda	 ->17	,->1	.->1	
rörde	 ->1	s->1	
rördh	e->1	
rörel	s->9	
rörig	t->2	
rörli	g->24	
rörs 	a->7	k->1	
rört 	d->2	e->1	
rörts	 ->2	
rös o	c->1	
rös p	o->1	
rös r	a->1	
rösa 	m->1	r->1	v->1	
röske	l->3	
röst 	-->2	f->1	h->3	i->2	m->1	o->1	s->1	t->2	
röst,	 ->2	
röst.	J->1	Ä->1	
rösta	 ->43	.->2	d->15	r->15	t->15	
röste	n->1	r->4	
röstf	ö->7	
röstn	i->57	
röstr	ä->3	
röstt	o->1	
röstv	i->3	
röt h	a->1	
röt t	a->4	
röts 	k->2	
rött 	k->1	
rött.	D->1	
rötta	 ->1	t->1	
rötte	r->4	
röva 	E->1	d->1	h->1	v->1	
rövad	e->1	
rövar	 ->2	e->2	
rövas	 ->2	.->2	
rövat	s->1	
röver	s->1	
rövni	n->5	
rövoå	r->1	
rövra	d->1	n->1	
rövst	a->1	
s "Bi	g->1	
s "ge	m->1	
s (PP	E->1	
s (fi	s->1	
s (un	g->1	
s - a	l->1	t->1	
s - b	i->1	
s - e	n->1	
s - f	ö->1	
s - h	a->1	
s - i	 ->1	n->1	
s - j	a->1	
s - m	e->1	
s - n	å->1	
s - o	c->6	m->1	
s - s	e->1	
s - t	v->1	
s -, 	s->1	
s 195	7->1	
s 196	7->1	
s 199	6->2	8->1	
s 2 4	0->1	
s 20 	º->1	
s 200	0->1	
s 24 	n->1	
s 28:	e->1	
s 3,8	 ->1	
s 400	 ->1	
s 80 	p->1	
s Ado	l->1	
s Alg	e->1	
s BNI	 ->2	
s BNP	 ->1	
s Bal	k->1	
s Bar	c->1	n->1	
s Blo	k->1	
s CEN	:->1	
s Dam	a->1	
s Del	o->3	
s EG-	d->2	
s EU-	f->1	m->1	
s Eur	o->13	
s FPÖ	 ->1	
s Gen	e->1	
s Gil	-->1	
s Gol	f->1	
s Hel	i->1	
s Isr	a->1	
s Lei	n->1	
s Mit	t->1	
s Oz,	 ->1	
s Pac	k->1	
s REP	 ->1	
s Rui	z->1	
s SOL	A->1	
s Sjö	s->2	
s Spa	n->3	
s VD 	b->1	
s Vic	h->1	
s Wie	b->1	
s Wur	t->1	
s XXV	I->1	
s abs	o->3	
s adm	i->1	
s age	r->3	
s akt	i->1	
s alb	a->1	
s ald	r->1	
s alk	o->1	
s all	 ->1	a->14	d->2	e->3	m->5	s->1	t->18	
s alt	a->1	
s amb	i->3	
s an 	d->1	f->2	
s ana	l->3	
s and	e->4	l->1	r->6	
s anf	ö->2	
s ang	e->2	å->3	
s anh	ä->1	
s ani	n->1	
s anl	e->2	
s anm	ä->4	
s ann	o->1	
s anp	a->1	
s ans	e->2	i->1	l->3	t->9	v->42	
s ant	a->3	i->2	
s anv	ä->3	
s arb	e->36	
s arg	u->2	
s ark	i->1	
s art	i->2	
s att	 ->172	,->1	a->1	
s auk	t->3	
s aut	o->1	
s av 	-->2	B->2	D->2	E->15	F->5	G->1	O->1	P->1	R->1	S->1	T->1	U->1	W->1	a->9	b->8	d->49	e->28	f->18	g->8	h->4	i->3	j->1	k->26	l->6	m->8	n->5	o->6	p->13	r->10	s->17	t->4	u->5	v->5	y->2	ä->1	å->1	ö->1	
s avd	e->1	
s avg	å->2	ö->4	
s avs	i->1	k->1	l->4	p->1	
s avt	a->1	
s avv	i->1	
s axl	a->1	
s bac	i->1	
s bak	o->1	
s bar	a->1	k->1	n->2	
s bas	a->1	e->1	
s bef	a->1	o->11	
s beg	r->6	ä->6	
s beh	a->1	o->5	ö->8	
s bek	l->2	
s bel	ä->1	
s ben	h->1	
s ber	o->2	ä->1	
s bes	k->1	l->28	t->6	ö->1	
s bet	e->1	o->1	y->8	ä->49	
s bev	a->1	i->2	
s bid	r->4	
s bil	d->1	i->1	p->1	t->1	
s bis	t->1	
s bl.	a->2	
s bla	n->4	
s bli	 ->3	c->1	n->1	r->2	
s blo	c->1	t->1	
s bor	t->8	
s bra	 ->1	n->1	
s bri	s->4	
s bru	k->1	
s bry	r->1	
s brå	d->1	
s bud	g->14	s->1	
s byg	g->1	
s byr	å->3	
s bär	a->1	
s bäs	t->3	
s bät	t->3	
s båd	a->2	e->2	
s bör	 ->1	
s cen	t->7	
s cir	k->1	
s cos	t->1	
s da 	C->5	
s dag	 ->2	,->1	a->1	l->1	o->11	
s dat	o->1	
s de 	a->2	d->1	e->2	f->1	g->3	h->1	k->1	l->3	m->1	n->3	p->1	s->2	t->2	å->1	
s deb	a->7	
s def	i->3	
s del	 ->1	,->1	a->1	e->6	s->2	t->11	v->2	
s dem	 ->3	a->2	o->8	
s den	 ->24	n->3	
s der	a->2	
s des	s->3	
s det	 ->87	,->2	t->12	
s dim	e->2	
s dip	l->2	
s dir	e->18	
s dis	k->2	t->1	
s dit	 ->1	
s dju	r->1	
s doc	k->2	
s dog	m->1	
s dok	u->4	
s dom	a->1	i->1	s->4	
s dra	g->1	s->1	
s du 	c->1	
s dub	b->1	
s där	 ->8	,->3	.->2	?->1	e->4	f->12	v->1	
s då 	f->1	t->2	
s död	 ->3	.->2	
s eff	e->6	
s eft	e->18	
s ege	n->10	t->2	
s egn	a->6	
s eko	l->1	n->29	
s ell	e->23	
s emb	l->1	
s eme	l->5	
s emo	t->2	
s en 	a->5	b->5	d->9	e->6	f->5	h->4	i->2	k->5	l->2	m->7	n->1	o->3	p->4	r->4	s->16	t->5	u->3	v->5	ä->1	ö->2	
s end	a->9	
s ene	r->2	
s enh	e->4	ä->5	
s enl	i->6	
s eno	r->1	
s ens	 ->1	k->1	
s env	i->1	
s erf	a->2	
s ers	ä->1	
s et 	o->1	
s ett	 ->42	
s eur	o->3	
s eve	n->1	
s exa	m->1	
s exe	m->3	
s exi	s->3	
s exk	l->1	
s exp	e->2	
s ext	e->2	
s fab	r->1	
s fak	t->4	
s fal	l->5	
s fam	i->3	
s fan	t->1	
s far	l->1	t->2	v->3	
s fas	o->1	t->3	
s fav	o->1	
s fel	,->1	a->1	
s fem	 ->1	t->1	
s fil	o->1	
s fin	a->3	n->3	
s fis	k->4	
s fjo	r->1	
s fla	g->5	
s fle	r->6	x->3	
s flo	r->1	
s fly	g->1	
s fol	k->6	
s fon	d->2	
s for	d->1	m->3	s->1	t->11	ê->1	
s fot	s->2	
s fra	m->55	
s fre	d->1	k->1	
s fri	a->4	h->2	k->1	v->2	
s frä	m->5	
s frå	g->14	n->28	
s ful	l->13	
s fun	d->1	g->1	k->6	
s fyl	l->1	
s fyr	a->1	t->1	
s fys	i->1	
s få 	b->2	e->1	g->1	m->1	p->1	s->2	
s får	 ->2	
s föl	j->4	
s för	 ->134	.->1	b->3	d->7	e->33	f->5	h->1	l->3	m->4	n->1	o->5	r->4	s->72	t->17	u->1	v->5	ä->2	
s gal	n->1	
s gan	s->1	
s gar	a->3	
s gas	k->1	
s ge 	o->1	
s gem	e->26	
s gen	e->5	o->29	t->2	
s geo	g->1	
s ger	 ->1	
s gil	t->4	
s giv	a->1	
s gjo	r->1	
s god	a->3	k->4	t->1	
s gra	n->4	
s gru	n->8	p->13	
s grä	m->1	n->4	
s grö	n->1	
s guv	e->1	
s gäl	l->1	
s gär	n->2	
s gå 	t->1	
s gån	g->2	
s går	 ->1	
s gör	 ->1	a->3	
s ha 	e->2	v->1	
s had	e->4	
s haf	t->1	
s ham	n->4	
s han	d->8	t->1	
s har	 ->31	,->1	m->1	
s hav	,->1	e->4	
s hek	t->1	
s hel	a->2	t->2	
s het	t->1	
s hin	d->1	
s his	t->7	
s hit	t->4	
s hjä	l->3	r->2	
s hop	p->2	
s hos	 ->3	
s hot	a->1	
s hur	 ->3	
s huv	u->4	
s hyc	k->1	
s häl	s->8	
s hän	d->5	v->1	
s här	 ->13	,->7	
s hål	l->2	
s hår	d->3	t->2	
s hög	a->1	t->1	
s höj	a->1	
s i 2	0->1	
s i A	d->1	m->3	
s i B	e->1	i->1	
s i D	a->1	
s i E	u->12	
s i F	ö->3	
s i G	e->1	o->1	
s i I	n->1	
s i J	o->1	
s i K	o->5	
s i L	a->1	o->1	
s i M	a->1	c->1	o->1	
s i P	P->1	
s i S	a->1	c->1	h->2	r->1	t->1	v->1	y->1	
s i T	a->3	
s i U	S->1	
s i a	b->1	l->1	r->4	t->1	v->1	
s i b	e->4	i->3	r->1	ö->1	
s i d	a->13	e->41	i->1	o->1	
s i e	f->1	n->10	t->8	
s i f	e->1	o->1	r->9	ö->16	
s i g	e->3	å->3	
s i h	a->5	e->3	å->1	
s i j	u->1	
s i k	a->4	o->4	r->1	
s i l	a->1	j->1	
s i m	a->3	e->1	i->2	å->1	
s i n	a->1	o->1	y->1	ä->2	
s i o	c->1	l->2	m->1	n->1	r->1	
s i p	a->2	o->4	r->6	
s i r	a->2	e->7	i->1	å->8	
s i s	a->6	e->2	i->3	k->1	l->2	m->1	o->1	p->1	t->5	y->1	å->1	
s i t	a->1	i->3	o->1	
s i u	t->2	
s i v	i->6	ä->2	å->8	
s i Ö	s->1	
s i ä	n->3	
s i å	r->1	
s i ö	v->3	
s ide	n->1	o->1	
s idé	e->1	n->1	
s ige	n->4	
s iho	p->1	
s ikr	a->2	
s ill	e->2	
s imm	u->1	
s in 	d->1	i->4	p->2	u->1	
s in,	 ->3	
s inb	l->2	
s ind	i->2	u->1	
s inf	ö->5	
s ing	a->5	e->20	r->2	å->2	
s ini	t->6	
s ink	o->4	
s inl	e->1	ä->3	
s inn	a->6	e->9	
s ino	m->15	
s inr	e->4	i->7	ä->1	
s ins	a->5	p->1	t->22	
s int	a->1	e->69	r->17	ä->1	
s inv	ä->3	
s irr	g->1	
s jag	 ->9	,->1	.->1	
s jor	d->2	
s ju 	a->1	s->1	
s jud	e->1	
s jur	i->11	
s jus	t->5	
s juv	e->1	
s jäm	s->1	
s kab	i->1	
s kal	l->3	
s kan	 ->9	s->1	
s kap	a->3	
s kat	a->1	
s kem	i->1	
s kl.	 ->6	
s kla	r->4	s->1	u->1	
s kli	m->1	
s kol	l->4	
s kom	 ->1	m->40	p->1	
s kon	c->1	k->25	s->11	t->4	
s kop	p->1	
s kor	r->4	t->1	
s kra	f->3	v->5	
s kre	t->1	
s kri	n->1	t->2	
s krä	v->1	
s kul	t->4	
s kum	u->2	
s kun	n->2	s->1	
s kus	t->5	
s kva	l->3	n->1	r->6	
s kvi	n->1	
s kvo	t->1	
s käl	l->1	
s kän	s->2	
s kär	n->2	
s köp	a->1	
s lag	 ->1	,->2	a->2	e->1	s->12	
s lan	d->6	s->1	
s le 	b->1	
s led	a->12	n->2	s->1	
s leg	a->5	i->2	
s let	t->1	
s lev	n->3	
s lib	e->2	
s lig	a->1	
s lik	a->9	n->1	s->2	
s lil	l->1	
s lin	j->1	
s lit	t->1	
s liv	.->2	s->8	
s lju	s->1	
s lob	b->1	
s log	i->2	
s lop	p->2	
s lov	o->1	
s luc	k->1	
s lug	n->1	
s läg	e->1	s->1	
s läm	p->2	
s län	d->5	g->1	
s lär	o->1	
s läs	e->1	
s lån	g->1	
s löf	t->2	
s löp	a->1	
s mak	t->5	
s man	 ->4	d->2	
s mar	k->2	
s mas	s->1	
s mat	c->1	
s med	 ->118	,->3	.->3	a->2	b->16	d->3	f->1	l->19	v->3	
s mel	l->15	
s men	 ->4	
s mer	 ->6	.->1	
s mes	t->3	
s met	o->3	
s mig	 ->1	
s mil	d->1	i->1	j->10	
s min	 ->1	a->1	d->2	i->1	o->1	s->2	u->2	
s mis	s->1	
s mon	o->2	
s mor	a->1	
s mot	 ->14	i->1	o->1	s->2	
s myc	k->17	
s män	 ->1	n->3	
s mär	k->2	
s mål	 ->5	,->3	.->2	:->1	i->1	
s mån	 ->4	a->1	g->15	
s mås	t->9	
s möj	l->15	
s mör	d->1	
s möt	e->3	
s nac	k->2	
s nam	n->6	
s nat	i->9	u->7	
s ned	 ->3	.->2	
s neg	a->4	
s ni 	i->1	s->1	
s nio	 ->1	
s niv	å->4	
s nog	a->1	
s nor	r->1	
s nu 	a->1	e->1	f->2	l->1	o->1	v->1	
s nuv	a->9	
s nya	 ->6	
s nyf	ö->1	
s nyl	i->4	
s nys	s->1	
s näm	l->2	n->2	
s när	 ->12	a->3	m->1	v->1	
s näs	t->1	
s någ	o->24	r->9	
s nöd	v->3	
s oac	c->1	
s oan	s->1	v->1	
s obe	r->3	
s obl	i->3	
s och	 ->188	,->1	
s ock	s->39	
s odi	s->1	
s odj	u->1	
s oen	i->1	
s off	e->4	i->1	
s oft	a->2	
s ofö	r->3	
s ohj	ä->1	
s ohö	v->1	
s oin	s->2	t->3	
s oku	n->1	
s ola	g->1	
s oli	k->6	
s olj	e->1	
s oly	c->1	
s olä	m->1	
s om 	3->2	H->1	L->1	a->19	b->2	d->13	e->4	f->1	h->5	i->6	m->4	n->2	o->3	r->1	t->1	v->3	y->1	ä->1	
s om)	;->1	
s om,	 ->1	
s om.	 ->1	D->1	J->2	M->1	V->1	
s omb	o->1	
s omf	a->5	
s omr	å->7	
s oms	o->1	
s omv	ä->1	
s ord	 ->3	:->1	e->2	f->34	
s org	a->5	
s ori	g->1	
s oro	 ->7	,->1	.->1	a->1	
s ors	a->1	
s oss	 ->2	.->1	
s osä	k->2	
s oti	l->3	
s otr	o->1	
s otv	i->1	
s ova	n->1	
s pap	p->1	
s par	l->3	t->19	
s pas	 ->1	
s pat	i->1	
s pel	a->1	
s pen	g->2	n->1	
s per	i->1	s->5	
s pha	r->1	
s pla	c->1	n->1	t->3	
s ple	n->1	
s pol	i->24	
s pop	u->1	
s por	t->3	
s pos	i->4	
s pot	e->1	
s poä	n->1	
s pra	x->1	
s pre	c->2	l->1	m->2	s->2	
s pri	n->7	o->3	s->1	v->2	
s pro	b->5	c->1	d->2	g->6	j->2	k->1	p->1	t->2	
s pub	l->1	
s pun	k->1	
s på 	9->1	E->3	a->9	b->5	c->1	d->16	e->38	f->7	g->8	h->1	i->4	j->3	k->3	l->4	m->8	n->4	o->4	p->2	r->6	s->10	t->2	v->16	Ö->1	å->1	
s på,	 ->1	
s på.	D->1	
s påp	e->3	
s påt	r->1	
s quo	 ->1	,->1	
s rad	i->1	
s ram	 ->2	v->1	
s ran	d->1	
s rap	p->15	
s ras	i->3	
s rat	i->1	
s rea	k->2	
s red	a->7	
s ref	e->1	o->4	
s reg	e->18	i->16	l->6	
s rek	o->3	
s rel	a->1	
s rep	u->1	
s res	e->2	o->10	p->1	t->1	u->9	
s ret	r->1	
s rig	o->1	
s rik	a->1	e->1	t->6	
s ris	k->4	
s ro,	 ->1	
s roc	k->1	
s rol	l->10	
s rot	s->1	
s run	t->3	
s rut	i->1	
s ryk	t->2	
s räd	d->1	
s räk	n->10	
s rät	t->40	
s råd	.->1	e->3	
s rör	a->1	e->1	l->1	
s rös	t->2	
s röt	t->1	
s sad	e->3	
s sak	 ->3	.->1	e->1	k->1	n->1	
s sam	a->2	b->1	h->1	l->2	m->17	o->1	s->2	t->9	
s sat	t->1	
s sci	e->1	
s se 	t->2	ö->1	
s sed	a->4	
s seg	e->1	
s sek	e->1	r->1	t->1	
s sem	e->1	
s sen	a->2	
s ser	b->1	
s ses	s->2	
s sex	,->1	
s sid	a->26	
s sif	f->1	
s sik	t->1	
s sin	 ->2	a->1	n->1	
s sis	t->1	
s sit	t->2	u->5	
s sjä	l->14	t->1	
s ska	d->1	l->14	p->3	t->3	
s ske	p->1	
s ski	c->2	l->1	
s sko	g->4	l->1	
s skr	i->2	
s sku	l->24	
s sky	d->1	l->2	
s skä	l->3	
s skö	r->2	t->1	
s sla	p->3	v->1	
s slo	t->1	v->1	
s slu	t->13	
s små	 ->2	
s sna	b->3	r->3	
s soc	i->12	
s sol	i->2	s->1	
s som	 ->107	
s spe	c->9	
s spå	r->1	
s spö	k->1	
s sta	b->1	d->1	r->1	t->7	
s ste	l->1	n->1	
s sto	d->1	r->3	
s str	a->11	i->1	u->16	y->1	ä->1	
s stu	d->1	n->1	
s sty	r->2	
s stä	l->6	n->1	r->1	v->1	
s stå	l->1	n->12	r->1	
s stö	d->15	r->1	t->1	
s sub	s->1	v->1	
s suv	e->6	
s sva	g->1	r->4	
s svå	r->5	
s syf	t->2	
s syn	 ->2	d->1	p->3	v->2	
s säg	a->2	
s säk	e->10	
s säl	j->1	
s sän	d->1	
s sär	a->1	s->7	
s sät	t->4	
s så 	a->5	d->1	e->1	h->1	k->2	m->1	s->6	
s såd	a->1	
s sål	e->4	
s sår	b->1	
s såv	ä->1	
s sön	d->2	
s ta 	h->2	u->1	
s tac	k->1	
s tak	t->2	
s tal	.->1	a->2	m->3	
s tan	k->2	
s tap	p->1	
s tek	n->2	
s ten	d->2	
s ter	r->5	
s tex	t->4	
s tid	 ->4	,->1	.->2	e->1	i->4	s->1	
s til	l->142	
s tio	 ->2	
s tjo	c->1	
s tju	g->1	
s tjä	n->11	
s tog	 ->1	
s tot	a->2	
s tra	d->1	n->1	
s tre	 ->3	,->1	
s tro	 ->1	d->1	r->2	t->2	v->7	
s tul	l->1	
s tur	 ->1	.->1	i->1	
s tvi	n->1	s->1	v->3	
s tvä	r->2	
s två	 ->4	n->1	
s tyd	l->6	
s typ	 ->3	
s tyv	ä->1	
s und	a->3	e->39	v->1	
s uni	l->1	
s upp	 ->28	,->4	.->8	d->3	e->1	f->7	g->9	l->1	m->3	n->5	r->1	s->1	
s ur 	e->1	m->1	
s urs	p->6	
s ut 	a->1	f->2	g->1	m->1	o->1	p->4	s->1	u->1	
s ut,	 ->4	
s ut.	D->1	F->2	G->1	K->1	
s uta	n->10	
s utb	i->2	r->1	
s utf	o->7	
s utg	j->1	å->2	ö->1	
s uti	f->3	
s utm	ä->7	
s utn	y->1	
s utr	e->2	i->2	y->1	
s uts	e->1	k->4	t->2	
s utt	a->23	r->2	
s utv	e->17	i->5	ä->1	
s utö	v->1	
s vac	k->1	
s vad	 ->5	
s val	 ->1	f->1	k->1	
s van	 ->1	
s vap	e->2	
s var	 ->3	a->16	d->1	e->1	f->1	i->4	j->3	t->1	
s vat	t->3	
s vec	k->1	
s ver	k->29	
s vet	e->2	
s vi 	a->2	e->1	f->1	j->1	k->1	m->1	s->1	u->1	
s via	 ->1	
s vic	e->1	
s vid	 ->19	a->4	
s vik	t->9	
s vil	j->4	k->1	l->12	
s vin	s->1	
s vis	a->2	s->4	
s vit	b->5	
s vol	u->1	
s vot	u->1	
s vux	n->1	
s väc	k->2	
s väg	a->1	e->1	n->15	r->5	
s väk	t->1	
s väl	d->2	j->1	s->1	
s vän	s->1	t->2	
s väp	n->1	
s vär	d->5	l->2	
s väs	e->1	
s vån	i->1	
s vår	 ->1	a->1	t->1	
s yrk	e->2	
s yta	.->1	
s ytt	e->10	r->8	
s äga	n->1	r->5	
s ägg	"->1	
s än 	e->1	p->1	
s änd	a->1	r->9	å->2	
s änn	u->7	
s är 	a->7	d->14	e->7	f->4	h->2	j->3	m->1	n->2	o->1	p->2	r->1	s->3	t->1	v->2	
s äve	n->7	
s åld	e->5	
s år 	-->1	2->1	
s år.	T->1	
s årh	u->1	
s årl	i->4	
s åsi	k->8	
s åst	a->3	
s åt 	a->2	d->5	g->1	h->1	n->1	r->1	s->2	t->1	ä->3	
s åt,	 ->1	
s åt.	N->1	
s åta	g->2	
s åte	r->5	
s åtg	ä->10	
s åtm	i->2	
s öde	 ->1	,->4	
s ögo	n->2	
s öka	d->3	t->2	
s öms	e->1	
s ömt	å->1	
s öns	k->2	
s öpp	e->2	
s öre	g->2	
s öro	n->1	
s öve	r->37	
s övr	i->1	
s! Ja	g->1	
s! Va	d->1	
s!Det	 ->1	
s!Eur	o->1	
s!För	 ->1	
s!Gen	o->1	
s!Her	r->1	
s!Vi 	b->1	
s".De	n->1	
s".Ja	g->1	
s".Ka	n->1	
s) fö	r->1	
s) oc	h->1	
s, 12	 ->1	
s, Ev	a->1	
s, Lu	x->1	
s, Mi	s->1	
s, St	o->1	
s, To	m->1	
s, Wu	l->1	
s, al	l->2	
s, an	d->2	s->1	
s, at	t->12	
s, av	 ->1	
s, be	l->1	s->1	t->1	
s, bl	.->1	
s, bä	r->1	
s, bö	r->1	
s, de	 ->1	n->1	s->1	t->4	
s, di	a->1	
s, dv	s->1	
s, dä	r->4	
s, då	 ->3	
s, ef	t->8	
s, el	l->2	
s, en	 ->5	l->1	
s, et	t->3	
s, eu	r->1	
s, fo	r->1	
s, fr	a->1	e->1	ä->4	å->1	
s, fö	r->15	
s, ge	n->2	
s, gi	v->1	
s, gö	r->1	
s, ha	r->3	
s, he	l->1	r->1	
s, hu	r->2	
s, hä	l->1	
s, i 	d->1	s->5	
s, in	k->1	n->1	o->1	t->5	
s, ja	g->3	
s, jo	r->1	
s, ka	n->1	
s, ko	m->6	
s, le	g->1	
s, me	d->5	n->20	
s, mi	n->1	s->1	
s, mo	t->1	
s, my	c->1	
s, mä	n->2	
s, må	s->1	
s, nä	m->3	r->4	
s, nå	g->2	
s, oc	h->44	
s, om	 ->8	
s, pa	r->1	
s, på	 ->6	
s, re	g->1	
s, sa	m->1	
s, sk	e->1	r->1	
s, so	m->10	
s, sp	e->2	
s, sä	l->1	r->1	
s, så	 ->10	s->3	v->2	
s, t.	e->1	
s, ti	l->1	
s, tr	a->1	o->2	
s, ty	c->1	
s, un	d->1	
s, up	p->1	
s, ur	 ->1	
s, ut	a->7	t->1	
s, va	d->1	r->3	
s, vi	l->8	s->1	
s, vä	d->1	
s, vå	l->1	
s, är	 ->4	
s, äv	e->2	
s, åt	e->2	m->2	
s- fö	r->1	
s- oc	h->42	
s-, u	t->1	
s-Car	p->1	
s-Jør	g->2	
s-bel	o->1	
s-bes	t->1	
s-bil	e->1	
s-de-	L->1	
s-för	k->1	
s-int	ä->2	
s-not	i->1	
s-nyt	t->1	
s-pro	g->1	
s-sit	u->1	
s. 11	 ->1	,->1	
s. De	s->1	t->2	
s. Eq	u->1	
s. Eu	r->1	
s. Me	n->2	
s. Pa	r->1	
s. Wa	l->1	
s. ar	b->1	
s. at	t->10	
s. de	n->2	s->1	t->1	
s. en	h->1	
s. er	t->1	
s. et	t->1	
s. fo	r->1	
s. fö	r->2	
s. gr	a->1	
s. ho	s->1	
s. hu	r->1	
s. i 	d->1	
s. id	é->1	
s. in	f->1	n->1	t->1	
s. ja	g->1	
s. ma	n->2	
s. me	d->1	
s. mi	n->1	
s. nä	r->1	
s. om	 ->2	
s. på	 ->1	
s. sp	e->1	
s. va	r->1	
s. vi	 ->1	
s.(EN	)->1	
s.)Åt	e->1	
s.- (	P->1	
s..(F	R->1	
s.All	a->1	m->1	t->1	
s.Anh	å->1	
s.Ant	a->1	
s.Att	 ->1	
s.Bet	r->2	ä->1	
s.Bev	i->1	
s.Bla	n->2	
s.Cen	t->1	
s.Dag	l->1	
s.De 	h->1	m->1	s->2	
s.Den	 ->11	n->4	
s.Des	s->2	
s.Det	 ->46	a->1	t->15	
s.Dir	e->1	
s.Där	 ->1	e->1	f->9	m->1	
s.Då 	f->1	g->1	m->1	ö->1	
s.Eft	e->2	
s.Eko	n->1	
s.En 	b->1	d->2	k->1	v->1	
s.End	a->1	
s.Enl	i->2	
s.Ert	 ->1	
s.Ett	 ->5	
s.Eur	o->3	
s.Fac	k->1	
s.Flo	r->2	
s.Fru	 ->4	t->1	
s.Frå	g->2	
s.För	 ->8	
s.Gen	e->1	o->3	
s.Gre	k->1	
s.Han	 ->1	
s.Hel	t->1	
s.Her	r->10	
s.His	t->1	
s.Hit	 ->1	
s.Hop	p->1	
s.Hur	 ->1	
s.Huv	u->1	
s.Här	 ->1	
s.I a	l->1	n->1	
s.I d	a->2	e->1	
s.I e	g->1	
s.I k	o->1	
s.I l	i->1	
s.I r	a->1	
s.I s	l->1	t->1	
s.I ö	v->1	
s.Ing	e->1	
s.Ino	m->1	
s.Int	e->1	
s.Jag	 ->28	
s.Jon	c->1	
s.Jus	t->1	
s.Jäm	s->1	
s.Kom	m->6	
s.Kon	k->1	
s.Kos	o->1	
s.Lan	d->1	
s.Led	a->1	
s.Låt	 ->2	
s.Man	 ->3	
s.Med	l->3	
s.Mel	l->1	
s.Men	 ->9	
s.Min	 ->2	
s.Myn	d->1	
s.Män	n->1	
s.Mån	g->1	
s.Ni 	f->1	
s.Nu 	h->1	ä->1	
s.När	 ->4	
s.Någ	r->1	
s.OLA	F->1	
s.Oav	s->1	
s.Om 	p->1	v->1	
s.Onö	d->1	
s.Par	l->3	
s.Per	s->1	
s.Pre	s->1	
s.Pro	c->1	
s.På 	l->1	u->1	
s.Rap	p->1	
s.Rea	k->1	
s.Red	a->1	
s.Res	t->1	u->1	
s.Råd	e->1	
s.Sam	t->2	
s.San	n->1	
s.Sed	a->1	
s.Slu	t->5	
s.Sna	r->1	
s.Som	 ->2	
s.Så 	k->1	
s.Tac	k->1	
s.Tal	a->1	
s.Tan	k->1	
s.Til	l->1	
s.Tyv	ä->1	
s.Und	e->4	
s.Utf	o->1	
s.Utm	a->1	
s.Vad	 ->4	
s.Var	 ->1	f->1	
s.Vi 	a->1	b->3	f->3	g->1	h->5	i->1	k->2	m->6	s->1	t->1	v->2	ä->3	
s.Vid	a->1	
s.Vil	l->1	
s.Vår	 ->1	t->2	
s.Ytt	e->2	
s.k. 	a->1	i->1	s->2	
s.Änd	r->2	
s.Änn	u->1	
s.Äve	n->2	
s.Åta	g->1	
s.Åtg	ä->1	
s/den	 ->1	
s/int	ä->1	
s: an	t->1	
s: at	t->1	
s: en	 ->1	
s: fö	r->1	
s: hö	g->1	
s: ko	m->1	
s: va	d->1	
s; at	t->1	
s; b)	 ->1	
s; de	t->1	
s; en	 ->1	
s; oc	h->1	
s; vi	 ->1	
s?. (	F->1	
s?.He	r->1	
s?Den	 ->1	
s?Ett	 ->1	
s?Frå	g->1	
s?Har	 ->1	
s?I s	å->1	
s?Ja,	 ->1	
s?Jo,	 ->1	
s?Kom	m->1	
s?Och	 ->1	
s?Sku	l->1	
s?Til	l->1	
s?Vil	k->2	
s?Är 	d->1	
sNäst	a->1	
sa (a	r->1	
sa - 	a->1	
sa 10	0->1	
sa 25	 ->3	
sa 35	 ->1	
sa PP	E->1	
sa Ry	s->1	
sa al	l->2	t->2	
sa am	b->1	
sa an	a->1	d->3	f->1	s->6	t->1	v->2	
sa ar	b->5	
sa as	p->2	
sa at	t->7	
sa av	 ->18	s->3	t->2	
sa be	b->1	f->3	s->7	t->3	
sa bi	l->5	
sa bl	i->2	
sa br	a->1	i->2	
sa bå	d->4	
sa bö	r->1	
sa ce	r->1	
sa da	g->1	
sa de	 ->5	l->3	m->1	n->5	s->1	t->8	
sa di	s->1	
sa do	k->2	
sa dr	a->1	
sa ef	f->1	t->1	
sa eg	n->1	
sa el	e->1	
sa en	 ->2	o->1	
sa er	 ->2	
sa fa	l->8	n->1	r->1	t->1	
sa fe	m->1	
sa fi	n->1	s->1	
sa fo	n->6	
sa fr	a->1	ä->1	å->21	
sa fu	l->1	
sa fö	r->22	
sa ga	r->1	
sa ge	m->5	n->1	
sa go	d->2	
sa gr	e->1	u->2	ä->3	
sa ha	d->2	m->1	r->1	
sa he	r->1	
sa hi	n->3	s->4	
sa ho	t->1	
sa hu	r->2	
sa hä	n->2	
sa hö	g->1	
sa i 	E->3	f->1	h->1	l->1	s->1	u->2	v->2	
sa in	 ->1	b->1	c->1	d->2	i->1	l->1	n->2	o->1	s->2	t->7	v->1	
sa ka	n->4	t->3	
sa kl	y->1	
sa ko	l->3	m->4	n->9	
sa kr	a->3	i->1	
sa ku	s->1	
sa kv	i->3	
sa la	g->2	n->1	
sa li	t->1	
sa lä	k->1	m->1	n->10	t->1	
sa lö	f->1	s->1	
sa ma	k->1	t->3	
sa me	d->12	n->2	r->3	
sa mi	g->1	n->5	s->2	
sa mo	n->1	r->1	t->1	
sa mä	n->1	
sa må	l->10	n->1	s->2	
sa mö	j->2	
sa ni	o->2	
sa no	r->1	
sa ny	a->1	
sa nå	g->1	
sa ob	l->1	
sa oc	h->18	
sa ok	l->1	
sa ol	y->1	
sa om	 ->6	r->8	s->6	v->1	
sa or	d->2	g->2	
sa os	s->1	
sa pa	r->5	
sa pe	n->8	r->2	
sa pi	r->1	
sa pl	a->3	
sa po	l->1	
sa pr	a->1	i->2	o->19	
sa pu	n->5	
sa på	 ->13	s->1	
sa re	d->2	g->13	k->2	s->5	
sa ri	k->7	s->2	
sa ru	t->1	
sa rä	t->1	
sa s.	k->1	
sa sa	k->3	m->5	
sa se	s->1	x->1	
sa si	f->2	g->6	n->4	t->1	
sa sj	ö->1	
sa sk	i->2	o->2	u->1	ä->3	
sa sl	a->1	u->1	
sa sm	å->2	
sa so	c->1	l->1	m->2	
sa sp	e->3	ä->2	
sa st	a->2	i->1	o->1	r->4	ä->1	å->2	ö->2	
sa sv	å->1	
sa sy	n->1	
sa sä	g->2	r->1	
sa så	 ->1	
sa ta	l->1	n->1	
sa te	r->1	x->1	
sa ti	d->2	l->13	
sa to	l->1	n->1	
sa tr	a->3	e->5	
sa tv	i->1	å->3	
sa ty	c->1	
sa un	d->5	
sa up	p->11	
sa ur	 ->1	
sa ut	a->1	n->2	s->1	v->1	
sa va	d->2	l->1	p->2	r->2	
sa ve	r->2	
sa vi	d->1	k->2	n->1	s->2	
sa vä	l->1	r->7	
sa vå	r->2	
sa äm	n->2	
sa än	d->25	n->1	
sa är	 ->7	
sa äv	e->1	
sa år	t->1	
sa åt	a->2	g->6	
sa öv	e->3	
sa!Lå	t->1	
sa, 5	0->1	
sa, b	l->1	
sa, d	j->2	v->1	
sa, e	n->1	
sa, f	u->1	ö->4	
sa, g	e->1	
sa, h	ö->1	
sa, l	å->1	
sa, m	e->2	
sa, o	c->1	
sa, s	a->1	o->1	
sa, u	t->1	
sa, v	i->1	
sa, å	t->1	
sa...	(->1	
sa.An	n->1	
sa.Ba	k->1	
sa.Bl	a->1	
sa.De	t->4	
sa.Dä	r->2	
sa.Eu	r->1	
sa.Fr	a->1	
sa.Fö	r->1	
sa.He	r->1	
sa.I 	d->1	f->1	
sa.Ja	g->3	
sa.Kä	r->1	
sa.Ma	n->1	
sa.Me	n->2	
sa.Mi	n->1	
sa.Rå	d->1	
sa.Sa	m->1	
sa.Up	p->1	
sa.År	 ->1	
sa?Pr	o->1	
sabel	 ->2	
sabet	h->1	
sabla	n->1	
sabon	 ->4	,->1	.->1	m->2	
saca 	s->1	
sace 	o->1	
sace.	D->1	J->1	
sad a	v->1	
sad d	a->2	
sad e	l->1	u->1	
sad g	i->1	
sad h	a->1	
sad o	c->1	m->2	
sad s	e->1	o->1	
sad t	i->6	
sad, 	f->1	v->1	
sad.D	e->1	
sad.J	a->1	
sad.V	i->1	
sade 	"->2	-->2	E->1	a->14	d->4	f->5	h->3	i->7	j->2	k->1	m->3	n->4	o->11	r->1	s->5	t->11	u->1	v->5	ä->2	
sade,	 ->14	
sade.	D->2	H->1	J->1	S->2	
sade:	 ->1	
sades	 ->2	,->1	
sadör	 ->1	
safet	y->1	
saffä	r->2	
safto	n->1	
sag i	 ->1	
sager	a->1	
sagt 	-->1	a->12	b->2	d->2	f->2	i->3	j->1	m->2	o->1	s->1	ä->1	
sagt,	 ->8	
sagt.	 ->1	
sagts	 ->10	,->2	
saill	e->1	
sak a	t->4	
sak b	e->2	
sak g	ä->3	
sak h	a->1	o->1	ä->1	
sak j	a->1	
sak k	o->1	
sak m	e->2	o->1	å->1	
sak n	ä->1	
sak s	j->1	o->8	
sak t	i->3	
sak u	t->1	
sak v	a->1	i->4	
sak ä	r->2	
sak, 	h->1	m->1	
sak.A	t->1	
sak.D	e->1	
sak.E	t->1	
sak.N	i->1	
sak.T	y->1	
sak: 	g->1	
saka 	e->2	o->1	p->1	r->1	
sakad	e->3	
sakar	 ->4	
sakas	 ->2	
sakat	 ->2	.->2	s->2	
saken	 ->7	,->2	.->1	:->1	?->1	s->3	
saker	 ->25	,->3	.->5	:->1	n->11	
sakfö	r->1	
sakku	n->2	
sakli	g->11	
sakna	d->5	r->12	s->20	t->2	
sakom	r->2	
sakpr	o->1	
sakre	r->1	
sakt 	o->1	v->1	
sakt.	B->1	
sakte	n->1	r->2	
sakti	o->1	v->1	
saktö	r->1	
sala 	v->1	
salem	 ->2	
salin	a->1	
salme	d->1	
salte	r->1	
saluf	ö->1	
sam a	c->1	r->1	s->2	
sam b	e->2	u->1	
sam c	o->1	
sam d	a->1	e->2	i->2	
sam e	r->1	u->2	
sam f	o->1	r->1	ö->2	
sam g	r->1	
sam h	e->1	å->1	
sam i	n->2	
sam l	a->1	ö->1	
sam m	a->2	e->3	i->1	
sam n	ä->1	
sam o	c->1	m->2	
sam p	o->1	å->4	
sam r	a->1	e->4	ä->1	
sam s	a->2	t->5	ä->3	
sam t	i->2	r->1	
sam u	t->2	
sam v	a->1	e->2	
sam å	k->1	t->1	
sam ö	k->1	v->1	
sam, 	n->1	o->1	
sam.I	 ->1	
samar	b->83	
samba	n->47	
samex	i->2	
samfi	n->1	
samfu	n->5	
samfö	r->7	
samhe	t->97	
samhä	l->47	
samka	r->1	t->2	
samla	 ->10	d->1	r->3	s->1	t->5	
samle	v->1	
samli	n->25	
samma	 ->250	,->4	.->2	d->1	n->228	r->5	s->2	
samme	 ->1	
samor	d->37	
samrä	t->1	
samrå	d->9	
samst	ä->4	
samsy	n->3	
samt 	G->1	H->1	a->12	b->4	d->2	e->7	f->11	h->1	i->3	j->1	k->5	l->3	m->5	n->1	o->9	p->2	r->6	s->7	t->4	u->7	v->1	y->1	ä->3	å->1	ö->1	
samt,	 ->2	
samt.	P->1	U->1	Å->1	
samta	l->16	
samti	d->53	
samtl	i->25	
samty	c->6	
samve	r->3	t->2	
san h	o->1	
san i	 ->2	
san o	c->2	
san t	i->1	
san ä	r->1	
san, 	k->1	ä->1	
san.M	e->1	
san.S	å->1	
san.V	a->1	
sanal	f->1	y->5	
sanda	 ->1	,->2	.->1	
sande	 ->11	.->1	l->3	t->1	
sanfö	r->1	
sankt	i->8	
sanlä	g->9	
sanmä	l->1	
sann 	e->1	
sanna	 ->1	
sanne	r->4	
sanni	n->3	
sanno	l->8	
sans 	n->1	
sansa	t->2	
sansp	r->1	
sanst	r->1	
sansv	a->1	
sant 	-->2	a->10	d->3	f->2	i->1	n->1	p->1	s->2	t->1	ä->1	
sant!	"->1	
sant,	 ->3	
sant.	D->1	V->1	
sant:	 ->1	
santa	 ->5	
sar a	n->1	t->9	
sar d	e->6	
sar e	l->1	m->1	n->3	r->1	
sar f	ö->3	
sar h	u->2	
sar i	 ->2	n->2	v->1	
sar j	a->1	u->1	
sar k	a->1	o->2	
sar m	a->1	e->1	i->1	
sar n	e->1	u->1	
sar o	c->4	m->1	s->1	
sar p	r->1	å->8	
sar r	e->2	
sar s	i->3	k->1	t->1	
sar t	i->6	r->1	y->2	
sar u	p->1	t->1	
sar v	a->4	e->1	i->2	å->1	
sar ä	n->1	v->2	
sar å	s->1	
sar!D	e->1	
sar, 	a->1	i->1	l->1	m->1	
sar.D	ä->1	
sar.S	å->1	
sarbe	t->27	
sare 	E->1	d->1	h->1	o->1	
sare.	V->1	
sargu	m->1	
sarna	 ->1	
sarti	k->3	
sas a	v->1	
sas b	e->1	o->1	
sas d	e->1	i->1	
sas e	f->1	
sas i	 ->2	n->1	
sas k	o->1	
sas m	e->1	å->1	
sas o	c->1	m->3	
sas p	å->1	
sas s	o->2	ö->1	
sas t	i->10	
sas v	i->1	
sas, 	i->1	
sas.D	e->1	
saspe	k->3	
sat a	l->1	n->1	t->8	
sat b	e->1	
sat d	e->2	
sat e	n->2	t->3	
sat f	i->1	
sat h	u->1	
sat i	 ->2	
sat m	e->1	o->1	
sat n	e->1	
sat o	c->1	s->1	
sat p	r->3	å->1	
sat s	i->8	ä->1	
sat t	i->1	
sat v	i->1	
sat, 	h->1	
sat.D	e->2	
sat.F	ö->1	
sat.H	e->1	
sat.N	i->1	
satel	l->1	
satio	n->46	
sator	 ->1	,->1	i->1	
sats 	a->2	f->2	i->1	o->2	p->1	s->1	t->13	u->1	ä->1	
sats,	 ->5	
sats.	D->1	H->1	J->1	
satsa	 ->7	r->3	s->2	t->1	
satse	n->20	r->65	
satsf	ö->1	
satsn	i->4	
satso	s->3	
satss	t->3	
satt 	b->1	d->3	e->1	f->2	i->1	l->1	o->2	r->1	s->4	t->1	u->1	v->2	ö->1	
satt,	 ->3	
satt.	D->1	N->1	
satta	 ->25	.->2	
satte	 ->3	s->6	
satts	 ->2	.->1	
sauro	,->1	
savbr	o->1	
savgi	f->1	
savgr	ä->1	
savgå	n->1	
savgö	r->5	
savi 	I->1	
savta	l->15	
savve	r->1	
sbank	e->2	
sbar 	h->1	
sbara	 ->1	
sbart	 ->3	
sbas.	D->1	
sbase	r->1	
sbedr	ä->2	
sbedö	m->2	
sbefo	g->1	l->2	
sbefr	i->6	
sbegr	e->1	ä->3	
sbeha	n->3	
sbeho	v->1	
sbekä	m->3	
sbela	g->4	
sbelo	p->2	
sbelä	g->1	
sberä	t->2	
sbesk	r->1	y->1	
sbesl	u->7	
sbest	ä->14	å->9	
sbesä	t->1	
sbeta	l->2	
sbeto	n->1	
sbetä	n->2	
sbeva	r->1	
sbevi	s->6	
sbidr	a->2	
sbild	n->7	
sbist	å->2	
sbola	g->3	
sbord	 ->1	e->2	
sbour	g->5	
sbris	t->2	
sbrot	t->2	
sbruk	 ->2	!->1	,->5	a->1	e->6	s->1	
sbudg	e->3	
sburn	a->1	
sbuss	a->1	
sbuti	k->1	
sbygd	 ->1	.->1	e->31	s->10	
sbygg	n->1	
sbåda	n->1	
sbörd	a->12	
scaya	b->2	g->4	
scen 	m->1	
scena	r->5	
scene	n->1	
scens	a->1	
scent	r->7	
scert	i->1	
sch f	ö->1	
sch i	 ->1	
sch o	c->1	
sch s	o->1	
sch! 	U->1	
sch.E	f->1	
sch?F	r->1	
schab	l->1	
sche 	B->1	
schef	e->12	
schem	a->1	
schen	 ->4	;->1	
scher	 ->1	a->1	n->2	
schho	f->1	
schle	r->4	
schwi	t->1	
scien	t->1	
scipl	i->14	
scism	,->1	e->2	
scist	 ->1	e->3	i->5	
score	b->1	
scyke	l->3	
sdag 	a->1	f->1	h->1	i->1	k->1	o->2	s->1	
sdag.	A->1	D->1	J->1	L->1	
sdag:	D->1	
sdage	n->1	
sdags	,->1	
sdeba	t->3	
sdel 	i->2	s->1	u->1	
sdel.	V->1	
sdela	r->8	
sdele	n->1	
sdepa	r->1	
sdigr	a->2	
sdikt	i->5	
sdime	n->1	
sdire	k->7	
sdoku	m->6	
sdom 	ä->1	
sdomi	n->1	
sdoms	t->2	
sdrab	b->4	
sdrän	g->1	
sdugl	i->5	
sduka	r->1	
sdömd	,->1	
sdömt	 ->1	
se (a	r->1	
se - 	a->2	e->1	
se Gr	o->1	
se an	s->1	
se ar	t->1	
se at	t->38	
se av	 ->14	
se ba	r->1	
se be	r->1	
se de	 ->2	m->1	n->6	r->1	s->1	t->5	
se do	m->1	
se el	l->1	
se en	 ->3	
se et	t->3	
se fo	r->1	
se fr	a->5	å->5	
se fö	r->22	
se ge	n->1	r->1	
se gi	v->1	
se ha	n->1	r->2	
se ho	n->1	s->1	
se hu	r->4	
se hä	r->1	
se i 	B->1	I->1	a->1	d->2	f->1	o->1	t->1	u->1	
se in	t->2	
se ja	g->2	
se ju	s->1	
se ka	n->2	
se ko	l->1	m->4	
se ly	s->1	
se me	d->16	l->2	r->2	
se mo	t->1	
se my	n->1	
se no	t->2	
se nä	r->3	
se oc	h->14	k->1	
se ol	i->1	
se om	 ->12	.->1	
se pe	s->1	
se på	 ->11	
se re	s->2	
se ri	k->1	
se sa	d->1	m->1	
se si	n->1	
se sk	a->1	u->1	
se sn	a->2	
se so	m->17	
se sp	å->1	
se st	a->1	
se sä	k->1	
se så	 ->1	
se ta	g->1	
se ti	l->70	
se un	d->1	
se up	p->2	
se ut	 ->1	,->2	
se va	d->3	r->1	
se ve	m->1	
se vi	l->10	
se än	d->1	
se är	 ->3	
se öv	e->14	
se", 	i->1	
se, d	e->3	
se, e	f->2	x->1	
se, i	 ->1	n->2	
se, j	a->1	
se, k	a->1	
se, l	i->1	
se, m	e->3	
se, s	k->1	
se, t	y->1	
se, u	r->1	
se, v	i->1	
se- o	c->1	
se-No	r->1	
se.Be	t->1	
se.De	n->2	t->4	
se.Ef	t->1	
se.En	l->2	
se.Et	t->1	
se.Fö	r->1	
se.Ja	g->3	
se.Ko	m->1	
se.Lå	t->1	
se.Ma	n->1	
se.Me	n->1	
se.Mi	n->2	
se.Ni	 ->1	
se.Om	 ->1	
se.Sa	m->1	
se.Sk	a->1	
se.Va	r->1	
se.Vi	 ->1	n->1	
se; j	a->1	
se?En	l->1	
seakt	 ->1	
sebal	l->1	
sebyg	d->1	
sed s	o->1	
sedan	 ->83	,->9	.->10	?->2	
sedd 	f->2	
sedda	 ->2	.->1	
seder	 ->1	
seend	e->60	
seffe	k->7	
seful	l->11	
seg t	e->1	
segdr	a->1	
seger	 ->2	.->1	n->1	
segla	 ->5	d->2	r->6	
segra	d->2	t->1	
sehin	d->1	
seill	e->1	
seism	i->2	
sekel	 ->2	,->1	s->1	
sekle	r->1	t->1	
sekon	f->2	o->24	
sekre	t->16	
sekti	o->2	
sekto	r->89	
sekun	d->3	
sekve	n->61	
sel f	a->1	ö->1	
sel i	n->1	
sel k	a->2	
sel m	e->1	
sel n	u->1	
sel o	c->5	
sel v	e->1	
sel ä	r->1	
sel å	t->1	
sel! 	J->1	
sel!T	i->1	
sel, 	A->1	d->1	n->1	v->1	ä->1	
sel- 	o->1	
sel-I	)->1	I->1	
sel.D	e->1	
sel.F	r->1	
sel.S	c->1	
selby	r->1	
seled	a->2	
selek	t->1	
selfe	d->1	
sell 	n->1	t->1	
sella	 ->1	
selod	l->1	
selsa	t->1	
selsä	t->102	
selös	 ->1	t->2	
semel	l->3	
semes	t->4	
semin	a->1	
semit	i->3	
semön	s->1	
sen "	E->1	
sen (	1->2	
sen -	 ->6	
sen 1	9->2	
sen 2	0->1	
sen E	U->1	u->1	
sen M	i->1	
sen a	l->2	n->1	t->22	v->24	
sen b	e->3	l->4	ä->1	ö->2	
sen d	e->2	o->2	u->1	ä->1	
sen e	l->1	n->1	
sen f	r->5	ö->11	
sen g	a->1	e->2	
sen h	a->7	e->1	o->1	ä->1	
sen i	 ->33	n->6	
sen k	a->1	o->5	u->1	
sen l	i->1	y->1	å->1	
sen m	a->1	e->14	i->3	y->1	å->4	
sen n	e->1	y->1	ä->1	
sen o	c->19	m->6	r->1	
sen p	å->5	
sen r	e->1	
sen s	a->2	e->1	k->13	o->13	t->2	å->1	
sen t	a->2	i->7	r->2	
sen u	n->1	p->1	t->4	
sen v	a->1	e->1	i->5	
sen ä	r->10	
sen ö	k->1	
sen!N	ä->1	
sen, 	B->1	P->1	d->4	e->3	f->3	h->1	i->2	k->1	l->1	m->1	n->1	o->6	p->1	s->7	t->3	u->4	v->1	ä->2	ö->1	
sen. 	D->1	J->1	M->1	
sen.A	n->2	t->1	v->1	
sen.D	e->17	
sen.E	m->1	
sen.F	r->2	ö->2	
sen.G	å->1	
sen.H	a->1	e->5	u->1	
sen.I	 ->2	n->1	
sen.J	a->8	u->1	
sen.K	o->1	
sen.L	å->1	
sen.M	e->2	i->1	
sen.N	i->1	ä->1	
sen.O	c->1	m->1	r->2	
sen.P	a->1	
sen.R	e->1	å->1	
sen.S	a->2	o->2	å->1	
sen.T	i->1	
sen.V	a->2	i->11	å->1	
sen.Ä	n->1	
sen; 	s->1	
sen?F	o->1	r->1	
senNä	s->2	
sena 	i->3	u->2	ö->1	
sena,	 ->1	
senad	 ->5	,->1	?->1	e->3	
senar	 ->1	e->29	
senas	 ->1	t->67	
senat	e->1	
senbe	r->3	
sende	 ->2	n->1	s->1	t->5	
senfä	r->1	
senhe	t->4	
senin	g->13	
senli	g->3	
senrö	t->1	
sens 	a->3	b->2	d->9	e->2	i->2	m->2	n->1	o->1	p->1	r->1	u->2	v->2	ö->1	
sens,	 ->1	
sensi	b->1	
sent 	i->1	s->1	t->1	
sent,	 ->1	
sent.	D->2	F->1	J->1	
senta	b->1	l->10	n->10	t->12	
sente	r->24	
sentl	i->26	
seomr	å->1	
separ	a->1	
septe	m->15	
ser -	 ->4	
ser 4	0->1	
ser A	r->1	
ser E	U->1	
ser a	l->3	n->4	r->1	t->121	v->3	
ser b	e->2	l->2	ö->3	
ser d	e->28	o->2	ä->1	å->3	
ser e	j->1	l->4	m->3	n->1	r->1	t->1	x->1	
ser f	o->2	r->20	ö->37	
ser g	ä->1	å->2	
ser h	a->5	o->1	u->1	ä->2	
ser i	 ->10	n->20	
ser j	a->38	
ser k	a->2	o->8	r->1	
ser l	e->1	
ser m	a->2	e->8	y->3	
ser n	a->1	i->2	u->1	ä->1	
ser o	c->36	l->2	m->8	
ser p	a->1	å->9	
ser r	e->1	i->1	å->3	
ser s	a->1	i->2	k->4	l->1	o->41	t->1	å->3	
ser t	i->16	
ser u	n->2	p->2	r->1	t->7	
ser v	a->9	e->2	i->19	å->1	
ser ä	r->5	
ser å	t->1	
ser ö	v->4	
ser!D	e->1	
ser, 	a->2	d->6	f->1	h->1	i->3	j->1	m->3	n->1	o->8	s->6	t->1	u->3	v->3	ä->1	
ser. 	H->1	M->1	
ser.(	A->1	
ser.-	 ->1	
ser..	(->1	
ser.9	0->1	
ser.A	l->1	
ser.B	e->1	
ser.D	e->10	ä->1	
ser.E	n->1	
ser.F	ö->1	
ser.H	e->2	
ser.I	 ->1	n->2	t->1	
ser.J	a->3	
ser.K	a->1	i->1	o->3	
ser.O	m->1	
ser.S	t->1	
ser.T	i->1	
ser.V	a->2	i->3	
ser: 	e->1	
ser?E	u->1	
ser?M	e->1	
ser?V	i->1	
sera 	a->4	b->2	d->14	e->9	f->2	g->1	h->3	i->2	k->4	l->1	n->1	o->6	p->2	s->4	u->2	ä->1	ö->1	
sera.	 ->1	
serad	 ->13	e->30	
seran	d->3	
serar	 ->22	,->1	
seras	 ->15	,->2	.->2	
serat	 ->6	,->1	.->3	s->5	
serb,	 ->1	
serbe	r->7	
serbi	s->6	
serbj	u->1	
seri 	m->1	n->1	
seri.	M->1	
serie	r->1	
serik	a->1	
serin	g->90	
seriö	s->7	
serli	g->13	
serna	 ->100	!->1	,->12	.->23	;->1	H->1	s->2	
sers 	f->1	
serva	t->11	
serve	r->4	
servi	c->7	
servt	r->1	
ses d	e->2	
ses f	ö->1	
ses g	e->1	
ses i	n->1	
ses m	e->1	o->1	ö->1	
ses p	h->1	
ses s	o->4	
ses t	i->1	
ses u	t->1	
ses v	a->2	
ses ö	v->5	
ses.A	n->1	
sesid	i->5	
sessi	o->6	
set -	 ->2	
set a	v->6	
set b	e->2	
set e	l->1	t->1	
set f	a->1	ö->5	
set h	i->1	
set i	 ->3	n->1	
set k	a->1	o->1	
set m	i->2	
set o	c->1	
set p	å->3	
set u	p->1	
set, 	o->1	
set.D	e->1	
set.F	r->1	
set.J	a->1	
setap	p->1	
setik	 ->1	
sets 	e->1	
sett 	a->10	b->1	d->3	e->3	f->3	h->2	i->3	k->1	l->1	m->5	n->2	o->6	p->2	s->3	u->2	v->4	ä->6	ö->1	
sett,	 ->3	
sett.	D->2	H->1	J->1	M->1	
sett:	 ->1	
setts	 ->2	
setêt	e->2	
seuro	p->1	
seutv	e->1	
sevis	 ->2	
sevär	d->8	t->6	
sewie	s->1	
sex a	l->1	v->1	
sex e	u->1	
sex m	i->1	å->10	
sex p	l->1	
sex t	i->1	
sex ö	v->1	
sex, 	s->1	
sexis	m->1	
sexmå	n->1	
sexpo	r->1	
sexto	n->1	
sexue	l->3	
sexvä	r->1	
sfakt	o->1	
sfall	 ->3	,->1	e->1	s->1	
sfara	 ->1	.->1	
sfas,	 ->1	
sfase	n->4	
sfast	i->1	
sfatt	a->11	
sfel,	 ->1	
sfele	n->1	
sfien	t->31	
sfina	n->1	
sfisk	e->3	
sflag	g->15	
sflot	t->2	
sflyg	n->1	
sfond	 ->1	e->21	
sford	o->1	
sform	e->3	u->1	
sfors	k->1	
sforu	m->2	
sfost	e->1	
sfri 	f->1	i->2	
sfria	 ->2	
sfrih	e->45	
sfris	t->10	
sfräm	j->4	
sfråg	a->14	o->30	
sfrån	v->1	
sfull	 ->2	.->1	a->2	h->1	t->10	
sfunk	t->2	
sfäre	n->1	
sfäst	 ->1	
sfång	a->1	
sförb	e->1	
sförd	e->10	r->3	
sföre	t->5	
sförf	a->16	
sförh	a->14	å->6	
sförk	l->5	
sförl	u->2	
sförm	å->8	
sföro	r->3	
sförs	l->214	t->2	ä->2	ö->1	
sgara	n->3	
sgase	r->4	
sgeme	n->1	
sgill	a->1	
sgiva	r->15	
sgivn	i->1	
sgrad	 ->3	e->2	
sgren	a->2	
sgrun	d->1	
sgrup	p->10	
sgrän	s->3	
sgynn	a->7	
sgå K	i->1	
sgå d	e->1	
sgås:	 ->1	
sgör 	d->1	
sh Pe	t->1	
sh Po	r->1	
sh, a	t->1	
shall	"->1	
shand	e->8	l->5	
shant	e->2	
shate	t->1	
shaus	s->1	
shave	n->1	
shem 	ä->1	
sherr	a->1	
shet 	i->1	k->1	m->1	o->8	p->1	s->2	v->1	
shet,	 ->4	
shet.	 ->1	B->1	D->1	L->1	
shete	n->25	
shets	p->1	s->2	
shind	e->11	
shing	t->3	
ship 	m->1	
shjäl	p->2	
shop,	 ->1	
shota	d->1	
shus.	E->1	
shush	å->1	
shämm	a->2	
shäns	y->1	
shåll	n->1	
siasm	 ->3	
siati	s->2	
sibil	i->1	
sida 	f->2	g->1	i->4	o->2	s->2	v->2	
sida,	 ->9	
sida.	D->1	F->1	H->1	I->1	J->1	O->1	V->1	Ä->1	
sida?	I->1	
sidan	 ->43	,->2	.->1	
sidar	i->1	
siden	t->9	
sides	 ->2	
sidia	r->21	
sidig	 ->5	a->1	h->1	t->6	
sidiä	r->1	
sidka	r->1	
sidoe	f->1	
sidor	 ->3	.->1	n->2	
sidue	r->1	
siell	 ->6	,->1	a->19	t->11	
sien 	h->1	i->1	o->2	
sien,	 ->1	
sien.	S->1	
siens	 ->1	
siera	 ->3	d->3	r->1	s->6	t->3	
sieri	n->34	
siffr	a->7	o->15	
sific	e->9	
sifie	r->5	
siful	l->1	
sig E	u->1	
sig O	L->1	
sig a	l->2	n->7	r->1	t->26	v->8	
sig b	a->4	e->3	l->1	o->1	r->1	ä->2	
sig d	e->9	i->1	j->1	o->1	ö->2	
sig e	f->1	l->1	m->3	n->9	t->4	
sig f	r->9	ö->27	
sig g	i->2	ä->1	ö->1	
sig h	e->1	u->3	
sig i	 ->24	h->1	n->13	v->1	
sig j	u->1	
sig k	a->1	v->1	ä->1	
sig l	ä->2	
sig m	a->4	e->11	i->1	o->4	y->4	å->2	ö->1	
sig n	a->1	e->1	o->1	ä->3	ö->1	
sig o	c->9	e->1	m->23	n->1	
sig p	e->1	o->1	r->1	å->24	
sig r	e->2	
sig s	a->1	i->3	j->11	k->1	o->3	t->3	ä->1	å->2	
sig t	.->1	i->23	v->1	y->1	
sig u	n->1	t->8	
sig v	a->9	i->1	ä->1	
sig ä	n->1	r->3	v->1	
sig å	s->1	t->12	
sig ö	v->4	
sig, 	a->1	d->2	e->1	f->1	g->1	h->1	n->1	
sig.A	v->1	
sig.B	r->1	
sig.D	e->2	
sig.E	m->1	n->1	
sig.H	e->2	
sig.J	a->2	
sig.K	o->1	
sig.M	a->1	
sig.S	a->1	
sig.T	a->1	
sig.V	a->1	i->2	
sig.Ä	r->1	
sig; 	d->1	
siga 	a->1	f->1	h->1	i->1	k->3	m->1	o->1	p->1	r->2	s->2	
siga,	 ->2	
signa	l->14	
signe	l->1	r->1	
sigt 	a->4	b->1	h->1	i->1	m->1	o->2	s->2	t->1	
sigt.	G->1	
sik i	 ->1	
sik m	å->1	
sike.	F->1	
siken	 ->1	
siker	,->1	
sikt 	-->2	F->1	a->21	b->2	e->1	f->2	g->1	h->1	i->2	k->5	m->2	o->9	p->1	s->8	v->2	ä->8	ö->1	
sikt,	 ->9	
sikt.	D->2	J->1	K->1	O->1	V->1	
sikta	d->1	r->1	
sikte	,->2	.->1	n->22	r->23	
sikti	g->76	
siktl	i->4	
siktn	i->2	
sikts	f->2	p->1	
sil e	n->1	
sila 	b->2	
silie	n->1	
silve	r->3	
simis	t->2	
simma	 ->1	
simul	a->2	
sin a	k->1	n->2	r->2	
sin b	e->4	i->3	r->1	u->2	
sin d	a->2	e->3	o->1	
sin e	g->7	k->3	n->2	x->2	
sin f	a->1	r->4	u->1	ö->6	
sin g	e->1	o->1	
sin h	a->3	e->12	u->1	ä->1	ö->2	
sin i	 ->1	n->3	
sin k	a->1	o->2	
sin l	i->3	
sin m	a->3	e->1	o->1	å->1	
sin n	a->4	u->2	y->1	ä->1	
sin o	b->1	c->1	r->5	
sin p	e->2	l->2	o->3	r->1	å->1	
sin r	a->1	e->2	i->2	o->6	ä->5	ö->1	
sin s	e->1	i->1	j->1	k->1	l->2	o->5	p->1	t->4	u->1	ä->2	
sin t	i->3	u->3	
sin u	n->1	p->5	t->3	
sin v	a->2	i->2	ä->1	
sin w	e->1	
sin ä	r->1	
sin å	s->2	
sin ö	n->1	
sin.B	e->1	
sina 	a->6	b->6	d->2	e->16	f->12	g->3	h->7	i->6	j->1	k->6	l->5	m->8	n->3	o->3	p->1	r->15	s->13	t->5	u->8	v->7	y->1	å->3	ö->1	
sindu	s->8	
sine 	d->1	q->2	
sinfo	r->2	
sinfr	a->1	
singf	o->20	
sinit	i->9	
sinna	t->1	
sinne	,->1	h->1	l->1	n->2	s->1	
sinni	g->1	
sinom	 ->1	
sinri	k->4	
sinsa	m->1	t->3	
sinse	m->3	
sinsp	e->2	
sinst	a->3	i->3	r->6	ä->1	
sinte	n->2	r->1	
sintr	e->1	
sion 	H->1	P->2	a->2	b->2	e->1	f->4	h->2	i->2	k->3	m->2	o->10	s->15	t->1	u->1	ä->1	å->2	
sion)	 ->2	
sion,	 ->4	
sion.	 ->1	D->2	F->1	I->1	J->1	K->1	S->1	V->2	
sion?	D->1	K->1	Ä->1	
sione	l->1	n->895	r->41	
sions	-->1	d->2	f->4	h->1	k->3	l->11	o->1	p->1	r->13	s->2	t->1	u->3	ä->1	
sionä	r->248	
sis a	v->2	
sis n	ä->1	
sis o	c->1	
sis, 	k->1	
sisk 	f->3	p->2	t->1	
sisk,	 ->1	
siska	 ->83	
siske	 ->2	
siskt	 ->6	
sism 	-->1	e->1	o->3	s->1	
sism,	 ->2	
sism.	D->1	O->1	V->2	
sisme	n->3	
sist 	a->3	f->1	k->2	v->1	ä->1	
sist,	 ->4	
sist.	G->1	
sista	 ->43	n->1	
siste	n->1	r->6	
sisti	s->11	
sistn	ä->2	
sitet	 ->1	
sitio	n->15	
sitiv	 ->18	,->1	a->23	l->2	t->31	
sitla	n->2	
sitlä	n->1	
sitru	t->1	
sitt 	a->20	b->11	d->1	e->7	f->8	g->1	h->1	i->1	j->1	k->1	l->5	m->9	o->1	p->3	r->4	s->8	t->1	u->3	v->1	y->4	ä->1	ö->2	
sitt,	 ->1	
sitta	n->1	
sitte	r->8	
sittn	i->2	
sittr	a->1	
situa	t->126	
siv a	v->1	
siv b	l->1	
siv k	v->1	
siv m	i->1	
siv r	o->1	
siv s	t->2	
siv t	a->1	
siv..	 ->1	
siva 	a->1	e->1	l->1	s->1	t->1	u->2	
sivar	e->1	
sive 	a->1	b->2	d->3	e->3	k->2	l->1	r->3	s->1	t->1	
sivt 	a->2	d->1	f->2	i->3	o->2	u->1	
siära	 ->1	
siäre	r->1	
sjovi	s->17	
sju g	å->1	
sju i	n->1	
sju m	o->1	
sju p	u->1	
sju r	e->1	
sju, 	å->1	
sjuk.	J->1	
sjuka	,->1	
sjukd	o->1	
sjukf	ö->1	
sjukh	u->6	
sjukv	å->3	
sjund	e->4	
sjunk	a->4	e->2	i->2	n->1	
sjuri	s->2	
sjutt	o->2	
själ,	 ->1	
själ.	F->2	
själe	n->2	
själv	 ->38	,->5	.->4	a->69	b->5	f->3	h->1	k->20	p->1	s->16	t->5	ä->1	
sjätt	e->19	
sjöfa	r->8	
sjömä	n->2	
sjön.	F->1	
sjönk	 ->3	.->1	
sjöss	 ->3	)->1	
sjötr	a->1	
sjövä	r->1	
sk - 	n->1	
sk TV	 ->1	
sk a 	p->1	
sk ag	i->1	
sk al	l->7	
sk an	a->1	d->1	g->2	t->1	
sk ar	t->3	
sk as	p->1	
sk at	t->2	
sk ba	l->2	s->2	
sk be	l->1	r->1	s->2	t->3	
sk bi	l->4	
sk bl	o->1	
sk bo	j->1	
sk br	o->1	
sk by	r->2	
sk bö	j->1	
sk ci	v->2	
sk da	g->1	
sk de	b->4	m->2	t->1	
sk di	a->2	m->1	s->4	
sk ek	o->1	
sk en	e->1	
sk er	s->1	
sk fe	d->1	
sk fi	e->1	l->1	
sk fl	a->2	
sk fo	n->1	r->2	
sk fr	a->2	å->2	
sk fy	s->1	
sk fö	r->6	
sk ge	m->1	n->2	s->1	
sk gl	u->1	
sk gr	u->1	ö->2	
sk ha	m->1	n->4	
sk hj	ä->2	
sk hä	n->1	
sk i 	s->1	
sk id	e->1	
sk im	m->1	
sk in	r->3	s->5	t->2	
sk jo	r->1	
sk ju	r->1	s->1	
sk jä	m->1	t->1	
sk ka	m->1	n->4	r->1	t->3	
sk kl	o->1	
sk ko	m->1	n->21	s->1	
sk ku	l->3	
sk kv	i->1	
sk la	g->5	
sk le	d->2	g->3	
sk li	v->5	
sk lä	k->1	
sk lö	s->1	
sk ma	k->3	r->2	t->1	
sk me	d->2	n->1	
sk mi	l->2	n->1	
sk mo	d->1	
sk my	n->2	
sk na	t->3	
sk ni	v->14	
sk nj	u->1	
sk nä	r->1	
sk oc	h->21	
sk of	f->3	
sk oj	ä->1	
sk om	s->1	
sk op	e->1	
sk pa	r->2	
sk pe	r->2	
sk pl	a->2	
sk po	l->15	ä->1	
sk pr	o->5	
sk pu	n->1	
sk ra	m->1	s->1	
sk re	f->3	g->3	n->2	t->1	
sk ri	s->1	
sk ro	l->5	
sk rä	t->1	
sk rå	d->1	
sk rö	r->1	
sk si	g->2	t->3	
sk sk	a->1	
sk sm	i->1	
sk so	l->2	m->3	
sk st	a->7	r->5	
sk sy	n->6	
sk te	r->1	
sk ti	g->1	l->5	
sk tr	a->2	
sk ty	p->1	
sk un	d->2	i->5	
sk up	p->3	
sk ur	s->1	
sk ut	b->2	m->2	v->8	
sk ve	r->1	
sk vi	l->1	
sk vä	g->2	
sk än	 ->1	
sk åk	l->13	
sk öv	e->2	n->1	
sk, e	f->2	
sk, f	ö->1	
sk, k	o->1	
sk, m	e->2	
sk, s	k->1	
sk-br	i->1	
sk-fr	a->1	
sk-is	r->1	
sk-sk	a->1	
sk. J	a->1	
sk.De	t->1	
sk.He	r->4	
sk.I 	b->1	g->1	
sk.In	f->1	
sk.Ja	g->1	
sk.Me	n->1	
sk.Om	 ->1	
sk.Vi	 ->1	
ska "	s->1	
ska E	u->3	
ska F	P->1	
ska K	u->1	
ska P	a->1	
ska T	V->1	
ska a	b->1	k->3	l->3	m->1	n->12	r->12	s->2	t->8	u->1	v->2	
ska b	a->4	e->34	i->12	l->1	u->5	y->3	å->1	ö->2	
ska c	e->3	
ska d	a->1	e->27	i->5	j->1	o->3	y->1	
ska e	f->2	k->8	l->2	n->3	r->3	t->3	x->5	
ska f	a->7	i->4	l->3	o->31	r->17	u->2	å->1	ö->45	
ska g	a->1	e->16	i->1	r->29	
ska h	a->10	e->1	i->2	o->1	u->1	ä->5	å->4	ö->1	
ska i	 ->6	d->1	m->1	n->76	s->1	
ska j	o->2	ä->1	
ska k	a->9	i->1	l->2	o->104	r->18	u->11	v->1	y->1	ä->3	
ska l	a->3	e->10	i->14	ä->10	ö->1	
ska m	a->9	e->33	i->9	o->5	y->15	å->16	ö->1	
ska n	a->3	e->1	i->2	o->1	u->1	ä->3	ö->2	
ska o	c->49	e->1	f->3	i->1	k->1	m->17	p->2	r->75	
ska p	a->17	e->7	l->5	o->14	r->29	u->5	å->2	
ska r	a->19	e->57	i->8	u->1	ä->6	å->18	ö->1	
ska s	a->10	c->2	e->4	i->13	j->2	k->14	l->2	o->29	p->3	t->40	v->3	y->10	ä->2	å->2	
ska t	a->3	e->8	i->10	j->1	r->4	v->1	y->1	
ska u	m->1	n->242	p->3	t->27	
ska v	a->9	e->10	i->7	o->2	ä->10	
ska ä	m->1	n->1	
ska å	k->4	t->14	
ska ö	a->1	g->1	s->1	v->2	
ska, 	b->1	e->1	f->2	h->2	k->1	m->3	n->1	o->1	r->1	s->3	ä->1	ö->1	
ska.D	e->1	
ska.E	f->1	m->1	n->1	
ska.F	ö->1	
ska.H	u->1	
ska.J	a->2	
ska.P	å->1	
ska.V	i->3	
ska: 	"->1	a->1	
skabe	l->1	
skad 	a->1	k->1	m->1	s->2	t->1	
skada	 ->9	!->1	,->1	.->1	d->2	n->1	r->6	t->4	
skade	 ->8	.->1	e->2	f->1	m->1	s->3	
skadl	i->10	
skado	r->25	
skaff	a->25	e->1	
skaka	d->1	t->1	
skal:	 ->1	
skala	.->1	n->2	
skald	j->1	
skali	g->3	
skall	 ->670	
skalv	 ->1	
skam 	f->1	o->1	
skam!	D->1	
skaml	i->2	
skamm	a->1	e->1	
skamp	 ->1	a->1	å->1	
skan 	-->1	I->1	a->4	f->2	o->4	s->1	v->1	ä->2	
skan,	 ->1	
skan.	V->1	
skana	l->3	
skand	a->9	e->20	i->2	
skans	 ->1	l->1	
skap 	-->1	a->22	b->2	d->3	e->1	f->3	g->1	h->1	i->7	k->1	m->2	n->1	o->15	s->11	t->1	u->2	v->1	
skap"	 ->1	!->1	,->1	
skap,	 ->16	
skap.	 ->1	D->7	E->1	I->2	J->2	S->1	T->1	V->2	
skap:	 ->1	
skapa	 ->100	d->4	n->24	r->29	s->13	t->10	
skape	n->125	r->22	t->97	
skapi	t->2	
skapl	i->37	
skaps	 ->1	-->1	a->2	b->3	d->1	f->1	i->14	k->3	l->3	m->20	n->11	o->1	p->7	r->18	s->4	å->2	
skar 	a->6	b->1	d->1	e->4	f->3	g->1	i->1	j->1	l->1	m->1	o->2	p->1	r->1	s->4	v->3	
skar,	 ->2	
skar.	M->1	O->1	V->1	
skara	n->1	
skare	 ->5	,->1	
skarn	a->2	
skarp	t->2	
skarr	i->1	
skart	e->1	
skas 	e->1	f->1	i->3	m->8	o->1	
skas,	 ->1	
skas.	F->1	
skast	e->1	
skat 	a->1	d->2	f->1	m->1	p->1	r->1	s->1	
skat,	 ->1	
skat.	D->1	H->1	
skats	 ->1	,->1	.->1	
skatt	 ->3	,->2	.->2	a->17	e->32	n->10	
skbed	ö->4	
skbes	t->4	
ske -	 ->1	
ske I	t->1	
ske a	n->1	t->1	
ske b	a->1	e->1	l->1	
ske d	e->4	
ske e	n->3	
ske f	i->2	ö->2	
ske g	e->2	ö->1	
ske h	a->2	
ske i	 ->5	n->8	
ske k	a->1	o->4	u->1	ä->1	
ske l	e->1	i->1	ä->2	å->1	
ske m	e->3	
ske n	i->3	
ske o	c->4	m->4	
ske p	r->3	å->5	
ske r	e->2	
ske s	k->1	n->1	o->1	ä->1	
ske t	a->1	i->1	y->1	
ske u	n->1	t->5	
ske v	a->1	i->2	o->2	
ske ä	r->5	v->1	
ske!Ä	v->1	
ske) 	f->1	o->1	
ske, 	d->1	m->1	o->2	u->1	å->1	
ske.-	 ->1	
ske.D	e->1	
sked 	l->1	o->1	t->1	
sked.	D->1	
skeda	 ->2	n->1	t->1	
skede	 ->3	.->1	t->3	
skekv	o->1	
skeln	 ->3	
skemå	l->3	
skemö	j->4	
sken 	a->7	f->6	g->1	h->1	i->2	
sken,	 ->1	
skeom	r->2	
skepp	 ->2	s->6	
skeps	i->1	
skept	i->8	
sker 	-->1	a->1	b->3	d->2	e->3	f->3	i->10	k->1	m->3	n->1	o->3	p->1	r->1	s->5	t->1	v->1	ä->1	
sker,	 ->1	
sker.	D->1	G->1	H->1	N->1	V->2	
skera	d->2	r->14	s->1	t->1	
skere	s->1	
skeri	k->1	p->1	s->2	u->1	
skern	a->6	
skerä	t->1	
skese	k->1	
sket 	(->1	i->2	
sket,	 ->1	
sketr	y->3	
skets	 ->1	
skett	 ->13	,->1	.->1	
skeva	t->2	
skfak	t->1	
skfri	t->1	
skfyl	l->1	
skför	e->1	
skhan	t->6	
skhet	.->1	
skick	 ->3	.->1	a->12	l->1	
skien	 ->1	,->1	
skift	e->6	
skild	 ->17	.->1	a->37	e->4	r->3	
skilj	a->10	e->10	t->1	
skill	i->2	n->45	
skilt	 ->129	
skin 	o->1	s->2	
skine	n->2	r->1	
sking	r->3	
skinl	i->1	
skipa	 ->2	n->1	
skipn	i->9	
skisk	 ->1	a->3	
skiss	 ->1	e->3	
skjut	a->13	e->7	i->5	s->5	v->1	
skkap	i->1	
skkom	m->2	
sklan	d->22	
sklar	a->1	
sklau	s->2	
sklig	 ->2	a->39	h->1	t->1	
sklim	a->2	
sknin	g->77	
skniv	å->1	
skoal	i->2	
skoef	f->1	
skofö	r->2	
skog 	e->1	f->1	i->1	
skoga	r->10	
skoge	n->5	
skogr	i->1	
skogs	a->2	b->6	f->1	k->1	o->1	p->1	s->4	u->1	ä->2	
skoha	n->3	
skola	 ->2	n->4	
skoli	v->3	
skoll	e->1	
skolo	r->3	
skomm	e->15	i->26	u->2	
skomn	a->3	
skona	d->1	r->1	
skonc	e->3	
skonf	e->144	
skonk	u->1	
skons	t->1	u->1	
skont	r->18	
skop,	 ->3	
skor 	d->2	f->4	h->2	i->7	l->2	m->1	o->2	p->1	s->15	t->1	u->1	v->1	ä->1	
skor,	 ->3	
skor.	D->1	
skorn	a->24	
skors	 ->14	
skort	 ->1	,->1	
skosl	ä->1	
skost	n->10	
skott	 ->20	,->2	.->4	e->135	s->5	
skour	i->1	
skov 	o->1	
skove	t->1	
skraf	t->48	
skrar	 ->1	
skrat	t->2	
skrav	 ->1	.->1	e->8	
skret	 ->1	
skrev	 ->6	s->2	
skrid	a->12	e->7	s->2	
skrif	t->22	
skrig	e->6	
skrik	.->1	
skrim	i->20	
skris	 ->3	e->1	
skrit	e->5	
skriv	a->11	b->1	e->25	i->8	n->8	s->8	
skrot	.->1	a->10	f->1	n->15	
skrov	 ->6	"->1	,->1	.->2	e->3	k->1	s->1	
skräc	k->9	
skräd	d->1	
skräm	d->1	l->1	m->3	
skrän	k->11	
skräp	n->1	
skt E	U->2	u->1	
skt K	o->1	
skt M	ü->1	
skt a	l->1	n->5	r->1	t->4	v->1	
skt b	e->6	i->10	l->1	r->1	u->1	y->1	
skt c	i->1	
skt d	e->3	
skt e	g->2	n->3	r->1	t->1	x->1	
skt f	a->3	e->2	i->2	l->1	r->1	u->1	ä->1	å->3	ö->10	
skt g	e->2	r->3	ö->1	
skt h	a->4	e->1	ä->1	å->2	
skt i	 ->1	n->11	s->2	
skt j	u->1	
skt k	a->1	l->1	o->6	u->2	v->1	ä->1	
skt l	a->3	e->1	
skt m	a->2	e->5	i->3	o->1	å->1	ö->1	
skt n	y->1	ö->2	
skt o	c->17	m->3	p->1	r->1	
skt p	a->4	e->3	å->3	
skt r	a->1	ä->2	ö->1	
skt s	a->2	e->10	i->1	k->4	o->1	p->1	t->8	v->2	y->2	ä->10	
skt t	a->6	e->1	i->1	o->1	v->1	
skt u	n->1	p->3	r->3	t->5	
skt v	a->8	e->1	i->3	ä->3	
skt ä	n->1	r->4	
skt å	t->1	
skt ö	g->1	l->1	
skt!N	ä->1	
skt, 	m->4	o->1	r->1	ä->1	
skt.(	P->1	
skt.A	l->1	
skt.B	e->1	
skt.D	e->4	
skt.G	e->1	
skt.J	a->2	
skt.S	l->1	
skt.Å	 ->1	
sktal	a->1	
skugg	a->2	b->1	
skuld	a->1	b->1	e->1	
skull	 ->13	,->2	.->3	e->478	
skult	u->9	
skunn	i->1	
skupp	g->1	
skur 	f->1	
skura	r->1	
skurs	 ->1	,->1	e->4	
skus 	s->1	
skuss	i->61	
skuta	 ->1	b->3	n->2	
skute	r->78	
skva,	 ->1	
skval	i->7	
skvot	e->3	
skvär	d->6	t->7	
sky f	ö->1	
skydd	 ->34	)->1	,->3	.->6	a->31	e->17	s->16	
skyfa	l->1	
skyhö	g->1	
skyld	i->29	
skyll	a->3	e->1	s->1	
skymt	s->1	
skynd	a->11	s->4	
skyvä	r->1	
skäl 	-->2	6->1	a->2	b->1	d->1	e->1	f->4	h->3	i->4	n->1	o->2	s->6	t->5	ä->2	
skäl,	 ->1	
skäl.	A->1	D->1	F->1	J->1	
skäle	n->3	t->8	
skäli	g->1	
skämd	a->1	
skämm	a->2	
skämt	s->1	
skänk	a->2	
skänn	a->1	
skäns	l->2	
skär 	n->1	p->1	
skärn	i->3	
skärp	a->8	n->1	t->2	
skärs	 ->1	
skåda	d->2	r->1	
skådl	i->6	
skådn	i->1	
skåle	n->1	
skår,	 ->1	
skönh	e->1	
sköpa	r->1	
skör.	K->1	
sköra	 ->2	
skörd	 ->1	a->1	e->1	
skört	 ->1	
sköt 	9->1	l->1	
sköta	 ->6	s->1	
sköte	r->1	
sköts	 ->2	.->1	e->5	
skött	 ->2	e->2	s->1	
skövl	a->1	
sla -	 ->1	
sla a	v->7	
sla f	ö->1	
sla g	å->1	
sla h	o->1	
sla m	e->4	å->1	
sla o	c->1	p->1	
sla".	B->1	
sla, 	c->1	r->1	
sla.B	i->1	
slade	 ->1	
slag 	-->2	1->18	2->7	3->5	4->8	5->2	6->2	a->14	b->9	d->3	e->4	f->33	g->7	h->15	i->22	j->1	k->7	l->1	m->3	n->3	o->31	p->2	r->3	s->60	t->58	u->2	v->4	ä->3	å->1	ö->1	
slag,	 ->33	
slag.	 ->1	)->3	.->1	D->7	F->4	H->4	I->2	J->5	K->1	L->1	M->2	P->1	S->1	T->1	U->1	V->4	
slag;	 ->1	
slag?	D->1	F->2	
slaga	r->1	
slage	n->69	r->1	t->68	
slagi	t->16	
slagn	a->16	i->17	
slagr	e->1	
slags	 ->15	d->1	f->1	k->1	t->9	
slakt	a->1	
slam 	l->1	
slan 	d->1	f->2	o->1	
sland	 ->8	,->1	.->2	e->5	s->1	
slapp	h->3	
slar 	m->5	
slat 	i->1	
slava	r->1	
slavi	e->1	
sleda	m->39	
slen,	 ->1	
slen.	K->1	
sler 	S->1	
slesk	a->1	
slesn	å->4	
slibe	r->1	
slier	n->1	
slig 	b->1	d->2	f->7	g->5	h->2	i->1	k->2	m->2	o->3	r->2	s->2	
sliga	 ->82	.->1	r->1	
sligh	e->13	
sligt	 ->29	,->2	.->1	
sling	a->2	
slinj	e->2	
slins	b->1	
slipp	e->2	
slira	r->1	
slist	a->48	
slita	 ->1	
slive	t->14	
slo o	c->1	
slo, 	W->1	s->1	
slobb	y->1	
slog 	a->1	b->2	e->3	f->1	i->3	m->1	t->1	v->1	å->1	
slogi	k->2	
slogs	 ->4	
slola	d->1	
slomä	s->1	
slopp	 ->1	,->1	
slor 	h->1	m->1	o->1	t->1	
slor.	J->1	
slott	s->1	
slove	n->1	
sluka	r->2	s->1	
slump	 ->3	.->1	
slumr	a->1	
slunt	o->1	
sluss	a->2	
slut 	-->1	8->2	9->1	a->6	b->1	e->1	f->7	g->1	h->4	i->8	k->3	l->3	m->1	n->1	o->26	p->11	s->14	u->4	v->3	ä->3	å->1	
slut,	 ->14	
slut.	 ->1	D->3	F->1	I->1	N->2	O->1	S->1	T->1	V->1	
slut;	 ->1	
sluta	 ->39	,->4	d->30	n->27	r->9	s->8	t->14	
slute	n->15	r->8	t->54	
slutf	ö->9	
slutg	i->8	
sluth	a->1	
sluti	t->4	
slutk	o->1	
slutl	i->38	
slutn	a->2	i->40	
slutp	e->1	
slutr	e->2	
sluts	 ->1	a->52	c->1	f->12	p->4	r->1	t->1	
slutv	e->1	
slutä	n->5	
slyck	a->18	
släck	a->2	e->1	
släge	 ->1	.->1	t->6	
slägr	e->1	
släka	r->1	
släkt	a->1	e->1	i->1	
slämn	a->2	
sländ	e->34	
släng	d->1	
släpa	d->1	
släpp	 ->2	,->1	.->1	a->6	e->5	h->1	s->1	t->3	
slå E	u->1	
slå a	t->6	
slå e	l->1	n->3	
slå f	a->6	
slå i	h->1	
slå k	o->4	
slå m	e->2	
slå n	å->1	
slå p	r->1	
slå r	å->1	
slå s	a->1	i->1	
slå v	a->2	e->1	i->1	
slåda	 ->1	
slåen	d->1	
slång	a->1	
slår 	B->1	a->7	d->3	e->6	f->1	i->4	j->4	k->2	m->2	n->1	r->1	s->2	t->1	v->6	ä->2	
slår"	.->1	
slår.	 ->1	M->1	
slår?	S->1	
slås 	a->3	b->2	d->2	e->1	g->2	i->11	m->1	p->1	t->2	
slås.	D->1	
slåss	 ->1	
slöja	d->1	n->1	r->3	s->1	
slös 	d->1	s->1	
slösa	 ->4	,->2	.->1	r->1	s->1	
slöse	r->3	
slösh	e->39	
slösn	i->2	
slöst	 ->3	
slöt 	a->1	d->1	v->1	
sm - 	m->1	
sm el	l->2	
sm et	c->1	
sm fö	r->1	
sm hä	n->1	
sm in	t->1	
sm må	s->1	
sm oc	h->12	
sm om	 ->6	
sm på	 ->1	.->1	
sm sa	m->1	
sm so	m->5	
sm un	d->1	
sm än	 ->1	
sm är	 ->1	
sm öv	e->1	
sm, a	l->1	
sm, f	r->1	
sm, i	d->1	
sm, m	e->1	
sm, n	a->1	å->1	
sm, o	c->2	
sm, s	p->1	
sm, v	i->1	
sm, ä	r->1	
sm.De	s->1	t->5	
sm.Dä	r->1	
sm.Fr	u->1	
sm.He	r->1	
sm.I 	n->1	r->1	
sm.Ja	g->1	
sm.Me	d->1	
sm.Nä	r->1	
sm.Oc	h->2	
sm.Va	d->1	
sm.Vi	 ->2	l->1	
sm?Vi	l->1	
smajo	r->1	
smakt	 ->2	.->1	e->1	
smakä	m->1	
sman 	t->1	
sman.	S->1	
smann	 ->1	a->1	e->12	
smark	n->15	
smask	i->2	
smatt	a->1	
smedb	o->9	
smedd	e->2	
smede	l->95	
smedi	a->3	
smedl	e->5	
smedv	e->2	
smeka	n->2	
smen 	-->2	i->2	o->5	p->1	s->1	ä->1	
smen,	 ->3	
smen.	O->1	
smen;	 ->1	
smen?	V->1	
smens	 ->4	
smer 	f->2	o->1	s->1	
smer.	V->2	
smern	a->3	
smeto	d->6	
smidi	g->3	
smilj	ö->5	
smini	s->16	
smisk	 ->1	a->1	
smita	 ->1	
smitn	i->1	
smitt	a->1	
smode	l->2	
smoln	 ->1	
smome	n->5	
smono	p->1	
smoto	r->1	
smugg	l->1	
smula	 ->1	
smuss	l->1	
smuts	a->2	i->1	
smynd	i->31	
smäde	l->1	
smält	n->1	
smän 	a->1	e->1	f->1	i->2	n->1	o->1	p->1	s->6	t->2	
smäng	d->2	
smänn	e->15	
smärk	e->1	
smärr	e->1	
smärt	a->1	s->1	
smäss	i->12	
små E	u->1	
små a	n->1	
små b	l->1	
små e	k->1	
små f	a->1	r->1	ö->2	
små l	ä->2	
små m	e->2	ä->1	ö->1	
små o	c->32	
små p	l->1	
små s	p->1	t->4	
små å	t->1	
små, 	m->1	s->1	
små.D	e->1	
småfö	r->5	
smågr	ä->1	
smål 	(->1	g->1	h->1	i->1	o->1	s->2	
smål.	B->1	Ä->1	
småle	n->1	t->1	
småls	s->1	
småni	n->4	
småsk	a->1	
smöjl	i->4	
smöns	t->1	
smöte	 ->1	t->1	
sna d	e->2	
sna m	ö->1	
sna n	o->1	
sna o	r->1	
sna p	å->4	
sna t	i->4	
sna, 	f->1	m->1	
snabb	 ->3	a->24	t->43	v->1	
snack	d->2	
snade	 ->4	
snar 	f->1	t->3	u->1	
snar.	D->1	H->1	
snara	r->23	s->13	
snark	o->1	
snarl	i->1	
snart	 ->26	.->1	
snat 	m->1	p->2	t->6	
snedl	ä->1	
snedv	r->12	
snier	 ->1	,->1	
sning	 ->44	,->2	.->10	a->31	e->14	s->7	
snitt	 ->7	,->1	e->5	l->1	s->1	
snivå	 ->15	,->4	.->5	?->1	e->5	n->3	
snorm	e->7	
snyck	e->1	
snyhe	t->1	
snäll	a->1	
snät 	o->1	
snäte	n->1	t->1	
snäva	r->1	
snåla	 ->2	,->1	r->2	
snåri	g->1	
snöjd	 ->1	a->1	
snöje	 ->1	
snövi	t->1	
so et	t->1	
so fa	r->1	
so i 	a->1	
so oc	k->1	
so är	 ->1	
so äv	e->1	
so, d	e->1	
so- o	c->1	
sochi	s->1	
socia	l->202	
socie	r->1	t->1	
socio	e->3	
sodli	n->1	
soeff	e->1	
soffe	r->2	
sofi 	o->1	s->1	
sofi,	 ->1	
sofin	 ->1	
sofis	k->1	
soft 	l->1	
sola 	s->1	
solda	t->2	
soler	a->6	i->1	
solid	a->30	e->3	
sollm	ä->1	
solsk	e->1	
solut	 ->38	a->3	i->99	
solyc	k->1	
som "	E->2	n->1	v->1	
som -	 ->3	
som 1	9->1	
som 2	0->1	
som 3	-->1	
som 4	0->1	5->1	
som A	g->1	h->1	l->1	m->1	p->1	
som B	S->1	a->1	e->5	l->1	o->1	r->1	
som C	e->1	o->2	
som D	a->4	e->1	
som E	G->2	U->6	h->1	l->1	u->31	
som F	B->1	P->1	r->2	ö->2	
som G	a->1	o->1	r->1	
som H	a->2	e->1	
som I	n->1	t->1	
som J	o->2	ö->1	
som L	a->3	l->1	
som M	a->1	c->1	
som N	e->1	
som O	f->1	
som P	a->3	r->1	
som R	a->1	i->1	o->1	
som S	e->2	k->1	
som T	h->1	o->2	u->1	
som W	a->2	
som a	 ->1	b->2	d->2	g->2	l->29	m->2	n->46	p->1	r->10	s->1	t->13	v->22	
som b	)->1	a->4	e->93	i->8	l->8	o->13	r->6	u->1	y->2	ä->5	å->2	ö->11	
som c	)->1	a->1	e->1	h->2	
som d	a->2	e->212	i->8	j->1	o->4	r->13	u->1	y->1	ä->7	å->3	ö->2	
som e	f->5	g->3	j->1	k->2	m->1	n->82	r->4	t->45	u->5	x->10	
som f	a->29	e->1	i->36	j->1	l->8	o->18	r->35	u->3	y->1	ä->2	å->9	ö->137	
som g	a->5	e->26	i->3	j->10	l->1	o->6	r->10	ä->21	å->11	ö->33	
som h	a->170	e->52	i->13	j->3	o->8	u->1	y->1	ä->28	å->6	ö->7	
som i	 ->81	f->1	n->134	
som j	a->102	o->1	u->12	
som k	a->56	l->1	o->97	r->20	u->1	v->1	ä->5	ö->2	
som l	a->14	e->35	i->22	y->5	ä->19	å->2	
som m	a->49	e->32	i->14	o->8	u->1	y->5	ä->2	å->25	ö->48	
som n	a->7	e->2	i->37	o->1	u->24	y->4	ä->8	å->10	ö->1	
som o	b->2	c->17	f->7	l->1	m->25	n->1	r->13	t->1	
som p	a->17	e->5	l->4	r->8	u->1	å->31	
som r	a->3	e->50	i->5	u->2	y->1	ä->6	å->19	ö->17	
som s	a->26	c->1	e->12	i->5	j->1	k->115	l->4	m->2	n->3	o->1	p->7	t->47	u->1	y->16	ä->11	å->13	ö->3	
som t	.->2	a->18	i->42	j->1	o->7	r->13	u->1	v->2	y->9	ä->4	
som u	n->20	p->26	r->3	t->39	
som v	a->35	e->17	i->241	o->3	r->1	u->1	ä->11	å->8	
som y	t->1	
som Ö	s->1	
som ä	g->4	n->13	r->168	t->1	v->12	
som å	k->1	l->2	s->5	t->10	
som ö	k->2	n->1	p->3	s->2	v->6	
som, 	d->2	e->4	g->1	i->4	j->2	o->1	p->1	s->1	u->2	v->1	ä->3	
somgi	v->1	
somli	g->3	
somma	r->3	
sområ	d->40	
somrö	s->1	
somsp	ä->1	
son a	n->1	
son f	ö->1	
son h	a->3	
son i	 ->2	n->1	
son k	a->1	
son o	c->1	
son s	o->2	
son v	a->1	
son, 	m->1	
son.N	i->1	
sonal	 ->8	,->2	.->3	e->1	f->1	p->3	r->3	s->1	u->1	
sonan	d->1	s->1	
sonel	l->2	
sonem	a->3	
sonen	 ->1	
soner	 ->29	,->4	.->2	;->1	n->3	s->1	
songs	b->1	
soni 	o->1	
sonin	g->4	
sonli	g->34	
sons 	t->1	
sonta	l->2	
sonte	l->1	
sopa 	a->1	
sor M	o->2	
sor T	e->1	s->2	
sor e	n->1	
sor m	e->1	
sor o	c->1	
sor, 	m->1	o->1	t->1	u->1	
sor.F	ö->1	
sor.J	a->1	
sorbe	r->1	
sordf	ö->21	
sordn	i->15	
sorel	a->1	
sorg 	a->1	o->7	s->1	
sorga	n->11	
sorgl	i->3	
sorgs	f->1	
sorie	n->1	
soris	k->3	
sorna	 ->1	
sorte	n->1	
sorts	 ->7	
sos o	c->2	
sos, 	k->1	
sosky	d->1	
sosäk	e->2	
sot s	o->1	
sovje	t->1	
sovo 	(->2	T->1	a->1	b->1	f->3	h->1	i->1	k->2	m->1	o->6	t->1	u->1	v->1	ä->3	
sovo,	 ->11	
sovo.	-->1	A->1	D->2	E->1	F->1	H->1	K->1	L->1	M->1	O->1	V->1	
sovo?	 ->1	H->1	
sovoN	ä->1	
sovok	o->1	r->1	
sovos	 ->7	
sovåd	l->1	
sovår	d->2	
sp", 	a->1	
sp. s	ä->1	
sp. t	r->1	
spake	t->4	
spakt	 ->1	e->3	
spane	l->1	
spanj	o->1	
spans	k->10	
spara	 ->4	r->3	
spari	n->3	
spark	 ->2	a->3	
sparl	a->1	
spars	a->1	
spart	e->1	n->3	
spati	e->2	
speci	a->14	e->42	f->29	
spegl	a->11	i->1	
spekt	 ->27	:->1	a->6	e->68	i->38	r->2	ö->6	
speku	l->4	
spel 	f->1	i->1	m->1	t->1	u->1	
spel,	 ->2	
spel.	D->1	I->1	
spel;	 ->1	
spela	 ->14	?->1	d->1	r->15	s->1	t->5	
spele	n->1	t->1	
speln	i->1	
spelp	l->1	
spelr	e->4	u->1	
spend	e->5	
spens	e->1	i->7	
speri	o->18	
spers	p->1	
spets	.->1	f->1	
spice	 ->1	
spill	o->1	
spin 	h->1	
spire	r->3	
spisk	a->1	
splac	e->3	
splan	 ->10	.->2	N->1	e->18	
splat	s->9	
splik	t->7	
split	t->4	
spo, 	s->1	
spoli	c->1	t->127	
spond	e->1	
spons	 ->1	r->1	
spont	a->4	
sport	 ->42	,->2	-->1	.->1	a->1	b->2	d->1	e->41	f->2	g->1	k->2	m->1	n->1	o->3	p->1	s->7	u->1	
spos 	b->1	
sposi	t->3	
spost	e->1	
spots	 ->1	
sprax	i->1	
sprid	a->4	e->5	i->1	n->8	s->2	
sprin	c->78	i->1	
sprio	r->1	
spris	e->3	
sprob	l->10	
sproc	e->53	
sprod	u->6	
sprog	r->32	
sproj	e->3	
sprot	o->1	
sprun	g->19	
språk	 ->5	.->1	a->9	e->3	l->3	o->2	t->1	
språn	g->2	
spunk	t->18	
spänn	a->4	i->7	
spärr	 ->1	a->2	
spåfö	l->1	
spår 	a->1	h->1	i->1	t->1	
spår,	 ->2	
spåra	 ->2	n->1	s->1	
spåre	n->1	
spårn	i->2	
spöke	 ->1	.->1	n->1	
spöks	t->1	
sque,	 ->1	
squin	s->1	
srad 	s->1	
srael	 ->22	,->4	-->1	.->3	?->1	e->5	i->15	k->1	s->6	
sram 	f->1	
sram,	 ->1	
srama	r->4	
srame	n->2	
srapp	o->6	
sreak	t->1	
sreda	r->2	
srefo	r->2	
srege	l->3	r->8	
sregi	o->4	s->3	
sregl	e->21	
sreko	m->5	
srela	t->1	
srepr	e->2	
srepu	b->4	
sresa	 ->2	
sreso	l->7	
sresu	l->1	
srik 	i->3	n->1	p->1	
srik,	 ->1	
srika	 ->4	,->1	
srikt	 ->5	.->1	
srila	n->1	
srisk	e->3	
sroll	e->1	
srubr	i->1	
sruhe	 ->1	,->1	
srum 	i->1	
srund	a->2	
sruti	n->1	
sryck	t->1	
srymd	 ->1	e->1	
sräds	l->1	
srätt	 ->3	,->1	.->1	e->50	i->2	s->4	
sråd 	-->1	f->1	
sråd,	 ->1	
sråd.	D->1	K->1	
sråde	t->4	
srådg	i->14	
sröre	l->2	
ss - 	j->1	
ss al	l->7	
ss an	 ->3	l->1	m->1	s->1	
ss ar	b->1	
ss at	t->29	
ss av	 ->4	s->2	
ss ba	s->1	
ss be	f->2	g->2	t->2	
ss bi	l->1	
ss br	a->1	i->1	
ss bu	d->1	
ss da	g->2	
ss de	 ->2	f->1	l->1	m->1	n->4	s->2	
ss do	c->1	m->2	
ss dä	r->6	
ss då	 ->2	
ss eg	e->1	n->2	
ss ek	o->1	
ss el	l->2	
ss em	e->2	
ss en	 ->7	h->1	l->2	
ss et	t->4	
ss eu	r->1	
ss ex	p->1	
ss fl	e->1	
ss fo	l->2	r->2	t->1	
ss fr	a->3	å->2	
ss fu	l->1	n->2	
ss få	 ->1	
ss fö	r->19	
ss ge	 ->1	m->3	n->1	
ss gj	o->1	
ss gr	a->1	u->1	
ss gä	l->1	
ss ha	d->1	r->3	
ss he	t->1	
ss hi	s->1	
ss ho	p->1	
ss hu	r->1	
ss hä	r->1	
ss i 	E->1	P->1	a->1	b->1	d->2	e->4	f->4	k->2	m->1	n->1	s->2	t->1	u->1	v->3	
ss id	é->1	
ss in	 ->1	d->1	f->1	n->4	r->1	s->2	t->6	
ss ka	l->1	
ss kl	a->1	
ss ko	m->4	n->3	
ss kv	a->1	
ss la	g->1	
ss le	d->1	
ss li	k->2	
ss lu	g->1	
ss lå	n->1	
ss ma	k->2	
ss me	d->11	l->1	n->1	s->1	
ss mi	l->1	
ss mo	r->1	t->2	
ss my	c->3	
ss mä	r->1	
ss må	l->1	n->5	
ss na	t->2	
ss ne	g->2	
ss ny	a->2	
ss nä	m->2	r->2	
ss nå	g->1	
ss oa	n->1	
ss oc	h->10	k->4	
ss od	i->1	
ss oe	n->1	
ss of	f->1	
ss om	 ->16	,->1	.->1	f->1	
ss or	d->4	o->3	
ss os	ä->1	
ss pa	r->1	
ss pe	r->1	
ss po	s->2	
ss pr	i->1	o->1	
ss på	 ->16	
ss ra	s->1	
ss re	g->1	l->1	s->3	
ss ry	k->1	
ss rä	t->3	
ss rö	r->1	
ss sa	d->2	m->4	
ss se	 ->1	
ss si	n->1	t->1	
ss sj	ä->10	
ss sk	a->1	o->1	y->1	
ss sl	a->1	u->2	
ss so	c->3	m->17	
ss st	r->2	ö->2	
ss sv	å->1	
ss sy	f->1	
ss sä	g->1	
ss så	 ->2	l->1	
ss ta	p->1	
ss ti	d->2	l->15	
ss tj	o->1	
ss to	t->1	
ss tr	e->1	o->1	
ss tv	i->1	
ss ty	p->2	
ss un	d->4	
ss up	p->1	
ss ut	a->1	f->1	n->1	s->3	v->1	ö->1	
ss va	d->1	r->6	
ss ve	r->3	
ss vi	 ->1	k->1	l->3	
ss vä	g->1	n->2	
ss vå	n->1	
ss yt	t->1	
ss än	d->2	n->1	
ss är	 ->10	
ss ås	i->2	
ss åt	 ->8	,->1	.->1	e->1	g->3	
ss öd	e->1	
ss öm	t->1	
ss ör	e->1	
ss öv	e->3	
ss".D	e->1	
ss) o	c->1	
ss, T	o->1	
ss, a	t->1	v->1	
ss, d	ä->1	
ss, e	f->1	
ss, f	ö->2	
ss, g	i->1	
ss, h	u->1	
ss, i	n->2	
ss, m	e->3	
ss, o	c->3	
ss, s	k->1	å->2	
ss, v	i->2	
ss, ä	r->1	
ss, å	t->1	
ss.Al	l->1	
ss.De	n->1	t->5	
ss.Di	r->1	
ss.Dä	r->1	
ss.En	 ->2	
ss.Eu	r->1	
ss.Fr	u->2	
ss.He	r->2	
ss.Ja	g->4	
ss.Ma	n->1	
ss.Må	n->1	
ss.Nä	r->1	
ss.Nå	g->1	
ss.Sl	u->1	
ss.Va	r->1	
ss.Vi	 ->5	
ss.Vå	r->1	
ss.Äv	e->2	
ss: k	o->1	
ss?. 	(->1	
ss?Jo	,->1	
ss?Vi	l->1	
ssa -	 ->1	
ssa 1	0->1	
ssa 2	5->3	
ssa 3	5->1	
ssa P	P->1	
ssa a	l->2	m->1	n->12	r->3	s->2	t->1	v->23	
ssa b	e->12	i->5	l->2	r->3	å->4	
ssa c	e->1	
ssa d	a->1	e->6	i->1	o->2	
ssa e	f->1	g->1	l->1	n->1	
ssa f	a->10	e->1	i->2	o->6	r->21	u->1	ö->20	
ssa g	a->1	e->5	o->2	r->4	
ssa h	a->4	e->1	i->6	o->1	u->1	ä->2	
ssa i	 ->3	n->16	
ssa k	a->7	l->1	o->11	r->4	u->1	v->3	
ssa l	a->3	ä->13	ö->2	
ssa m	a->3	e->13	i->5	o->2	ä->1	å->9	ö->2	
ssa n	i->2	o->1	y->1	
ssa o	b->1	c->1	k->1	l->1	m->17	r->3	
ssa p	a->4	e->10	i->1	l->3	o->1	r->14	u->5	å->4	
ssa r	e->21	i->9	u->1	ä->1	
ssa s	.->1	a->8	e->2	i->3	j->1	k->6	l->2	m->2	o->3	p->5	t->8	v->1	y->1	ä->2	å->1	
ssa t	a->2	e->2	i->3	o->1	r->8	v->3	y->1	
ssa u	n->4	p->6	t->2	
ssa v	a->3	i->3	ä->8	
ssa ä	m->2	n->25	r->4	v->1	
ssa å	r->1	t->8	
ssa ö	v->2	
ssa!L	å->1	
ssa, 	f->2	s->1	u->1	
ssa.B	l->1	
ssa.D	e->1	ä->1	
ssa.I	 ->1	
ssa.J	a->1	
ssa.M	a->1	e->1	i->1	
ssabo	n->8	
ssad 	h->1	o->1	s->1	t->2	
ssad,	 ->1	
ssade	 ->2	
ssadö	r->1	
ssag 	i->1	
ssage	r->1	
ssakr	e->1	
ssala	 ->1	
ssama	r->3	
ssamh	ä->5	
ssamm	a->1	
ssamt	a->5	
ssand	e->3	
ssank	t->1	
ssant	 ->14	,->1	.->1	a->5	
ssar 	e->1	o->1	p->1	v->1	
ssar,	 ->1	
ssarb	e->3	
ssarn	a->1	
ssas 	d->1	e->1	i->1	s->1	t->3	
ssat 	e->1	
ssavg	å->1	
ssbel	a->4	ä->1	
ssbru	k->10	
ssche	m->1	
sse (	a->1	
sse a	n->1	t->2	v->3	
sse d	e->3	
sse f	ö->5	
sse l	y->1	
sse o	c->1	
sse p	å->1	
sse s	a->1	o->1	
sse t	a->1	
sse, 	d->2	e->1	s->1	v->1	
sse-N	o->1	
sse.F	ö->1	
sse.M	a->1	i->1	
sse?E	n->1	
ssed 	s->1	
ssekr	e->1	
ssekt	o->18	
ssel 	f->2	i->1	k->2	m->1	n->1	o->1	v->1	ä->1	å->1	
ssel!	T->1	
ssel,	 ->5	
ssel-	 ->1	I->2	
ssel.	F->1	S->1	
sselb	y->1	
sself	e->1	
sselo	d->1	
ssels	a->1	ä->102	
ssen 	-->1	1->1	a->2	b->1	d->1	e->1	f->3	h->3	i->11	k->2	l->2	m->5	n->1	o->10	s->10	u->1	ä->2	
ssen,	 ->21	
ssen.	A->1	D->5	F->3	H->4	I->2	J->5	M->2	S->4	V->6	
ssen?	F->1	
ssenN	ä->1	
ssena	 ->4	,->1	
ssens	 ->7	
ssent	e->1	
sser 	-->1	A->1	i->1	m->1	o->1	
sser,	 ->2	
ssera	 ->4	d->8	r->5	s->1	t->1	
sseri	e->1	
sserl	i->13	
ssern	a->8	
sserv	i->1	
sset 	-->1	a->1	e->1	m->1	
sset,	 ->1	
ssetê	t->2	
ssfal	l->1	
ssfor	m->1	
ssfos	t->1	
ssför	h->1	s->3	
ssgyn	n->7	
sshet	 ->4	
sshus	h->1	
sshän	s->1	
ssida	n->1	
ssiff	r->3	
ssifi	c->9	
ssig 	a->1	b->1	k->1	
ssiga	 ->13	,->2	
ssigt	 ->13	.->1	
ssil 	e->1	
ssila	 ->2	
ssimi	s->2	
ssin 	i->1	
ssion	 ->41	,->2	.->4	?->3	e->906	s->20	ä->247	
ssisk	 ->1	a->2	t->2	
ssist	a->1	e->1	
ssitu	a->4	
ssiv 	a->1	m->1	s->1	
ssiv.	.->1	
ssiva	 ->4	
ssivt	 ->4	
ssjöf	a->1	
sskad	l->1	o->2	
sskan	d->1	
sskap	a->1	
sskat	t->1	
ssked	e->3	
sskic	k->1	
sskif	t->2	
sskil	j->4	l->1	
sskip	a->1	n->2	
sskon	f->2	
sskri	v->1	
sskro	v->7	
sskyd	d->3	
sskyl	d->2	
sskäl	 ->3	
ssköt	s->5	t->1	
ssla 	m->1	
sslad	e->1	
sslan	 ->1	d->5	
sslar	 ->5	
sslat	 ->1	
sslyc	k->18	
sslös	e->1	n->1	
ssmed	d->1	i->3	
ssna 	n->1	p->4	t->4	
ssna,	 ->1	
ssnad	e->4	
ssnar	 ->3	.->2	
ssnat	 ->9	
ssnin	g->7	
ssnöj	d->2	e->1	
sso e	t->1	
sso i	 ->1	
sso o	c->1	
sso ä	r->1	v->1	
sso, 	d->1	
ssoci	e->1	
ssoni	 ->1	
ssor 	M->2	T->3	e->1	o->1	
ssor,	 ->2	
sspel	a->1	
sspri	d->1	
ssprå	n->1	
ssreg	l->1	
ssres	o->2	
ssrät	t->2	
sst b	e->1	
sst d	a->1	
sst f	o->1	
sst j	u->1	
sst k	a->1	o->1	
sst m	i->1	
sst n	ä->1	
ssta 	o->1	
sstad	g->1	i->2	
sstag	 ->2	,->1	.->3	e->2	
sstan	d->3	k->4	
sstar	 ->2	t->1	
sstat	 ->28	,->5	.->8	e->239	l->2	s->11	
sstav	 ->1	
sste 	a->2	d->1	v->1	
sstex	t->1	
sstil	 ->1	
sstol	k->1	
sstra	t->11	
sstro	e->2	t->1	
sstru	k->5	
ssträ	v->2	
sströ	m->4	
sstyr	k->6	n->1	
sstäl	l->24	
sstäm	d->1	m->19	n->1	
sstän	k->4	
sstål	s->1	
sstêt	e->1	
sstöd	 ->9	,->4	.->5	;->1	e->10	s->1	
sstör	n->1	
ssuel	l->1	
ssupp	f->2	
ssuse	n->1	
ssuto	m->61	
ssvär	r->4	
ssvår	i->1	
ssyne	n->1	
ssynp	u->1	
ssys 	f->1	
ssyss	e->1	
ssyst	e->55	
ssäke	r->65	
ssäkr	a->1	
ssäll	s->7	
ssänk	n->1	
ssätt	 ->8	.->2	
st - 	f->1	s->1	v->1	
st 1 	0->1	
st 10	 ->1	
st 12	 ->1	
st 25	 ->1	
st 3 	p->2	
st 40	0->1	
st 5,	5->1	
st 70	0->1	
st 9 	f->1	
st Da	l->1	
st Eu	r->3	
st In	t->1	
st Mi	d->1	
st Pe	t->1	
st ac	c->2	
st ak	t->1	
st al	b->1	l->3	
st an	g->1	m->1	s->4	t->3	
st ar	b->2	t->1	
st at	t->12	
st av	 ->11	l->2	s->2	t->1	
st be	f->1	h->2	k->1	r->3	s->2	t->2	
st bi	l->1	
st bl	i->1	
st ca	s->1	
st da	t->1	
st de	 ->7	f->1	m->1	n->2	s->1	t->13	
st dr	a->4	
st dy	n->1	
st dä	r->6	
st då	 ->2	l->1	
st ef	t->5	
st en	 ->8	
st er	i->1	
st et	t->8	
st ex	p->1	
st fa	n->1	s->3	
st fl	e->1	
st fo	g->1	
st fr	a->6	e->1	å->2	
st fu	l->1	
st få	 ->2	
st fö	r->28	
st ge	n->4	r->1	t->1	
st gj	o->3	
st gl	ä->2	
st gr	u->1	
st gä	l->1	
st gå	 ->1	
st gö	r->2	
st ha	 ->3	f->2	r->15	
st hä	r->3	
st hö	r->1	
st i 	E->1	I->1	N->1	a->1	b->3	d->5	e->2	f->2	m->1	n->1	o->1	s->4	v->3	
st il	s->1	
st in	n->2	o->4	r->1	s->1	t->7	v->1	
st ju	r->1	s->1	
st ka	n->7	
st ko	m->5	n->3	r->1	s->1	
st kr	a->1	i->2	ä->1	
st ku	n->4	
st la	n->2	
st le	d->1	
st li	k->1	
st lo	t->3	
st lä	m->1	s->1	x->1	
st lå	n->2	
st lö	n->1	s->1	
st me	d->7	l->1	n->2	r->1	
st mi	n->3	s->2	t->1	
st mo	d->1	t->4	
st må	n->1	s->8	
st mö	j->3	
st ne	g->1	
st ni	o->1	
st no	g->1	t->1	
st nu	 ->10	
st ny	a->1	
st nä	m->1	r->9	
st nå	g->1	r->1	
st nö	d->1	
st ob	s->1	
st oc	h->34	
st of	f->1	
st ol	y->1	
st om	 ->9	d->1	r->1	
st op	t->1	
st or	d->1	
st ov	ä->1	
st pe	k->1	n->1	r->3	
st pl	a->1	
st po	l->1	p->1	r->1	
st pr	e->1	i->2	o->3	
st på	 ->29	?->1	
st ra	t->1	
st re	k->1	n->1	p->2	s->1	
st ri	m->1	s->1	
st ru	b->1	
st rä	c->1	t->1	
st rö	r->2	s->1	
st sa	d->3	g->2	m->2	
st se	d->1	r->2	x->1	
st si	g->1	
st sk	a->6	e->1	i->1	u->6	ä->1	
st sl	u->1	
st so	m->7	
st st	r->2	ä->1	ö->4	
st sv	a->1	å->2	
st sy	f->1	m->1	
st sä	g->1	t->2	
st så	 ->2	
st ta	 ->1	c->5	
st ti	d->1	l->15	
st tr	a->1	e->2	o->1	
st tv	e->1	i->1	å->2	
st tä	n->1	
st un	d->1	
st up	p->3	
st ut	a->2	n->1	o->1	s->3	t->2	v->3	ö->1	
st va	d->2	g->1	k->1	r->3	
st ve	m->1	
st vi	 ->4	d->10	k->7	l->16	
st vä	l->2	x->1	
st är	 ->11	
st år	 ->1	
st åt	 ->1	e->1	f->1	g->1	
st ön	s->1	
st öv	e->3	
st!Dä	r->1	
st!Tv	ä->1	
st, P	V->1	
st, a	t->1	
st, d	e->3	ä->2	
st, e	f->3	n->1	
st, f	r->1	
st, h	e->2	
st, i	n->2	
st, k	o->1	
st, m	e->2	i->1	
st, o	c->1	m->1	
st, p	å->1	
st, s	o->1	å->1	
st, v	i->1	
st- o	c->1	
st-be	n->5	
st. A	v->1	
st.Ac	c->1	
st.De	 ->1	n->1	t->1	
st.Ef	t->1	
st.Fö	r->2	
st.Gi	v->1	
st.Ja	g->3	
st.Ko	m->1	
st.Kä	r->1	
st.Me	d->1	
st.Mi	n->1	
st.Nu	 ->1	
st.Nä	r->1	
st.Va	d->1	
st.Vi	 ->3	
st.Är	 ->1	
st: m	i->1	
st?Ne	j->1	
st?Vi	 ->1	
sta a	d->1	l->2	n->3	t->4	v->7	
sta b	e->17	i->1	r->1	u->2	ö->2	
sta c	h->1	
sta d	a->3	e->22	i->4	
sta e	f->1	m->5	n->1	r->5	
sta f	a->5	e->1	r->12	ö->34	
sta g	a->2	e->6	r->5	ä->6	å->21	
sta h	a->32	i->1	
sta i	 ->4	g->2	n->9	
sta k	l->2	o->9	u->1	v->1	ä->2	
sta l	a->1	i->2	ä->1	
sta m	a->3	e->9	o->2	å->7	ö->18	
sta n	a->1	o->1	y->2	ä->3	
sta o	c->4	f->1	l->2	m->7	r->2	s->1	
sta p	l->1	o->2	r->8	u->37	å->4	
sta r	a->15	e->13	i->3	u->1	ö->2	
sta s	a->9	i->2	k->6	l->2	m->2	o->5	t->9	v->2	y->1	ä->13	
sta t	a->6	e->3	i->5	j->1	o->3	r->1	y->1	
sta u	n->1	p->2	r->1	t->4	
sta v	a->3	e->1	i->11	ä->3	
sta ä	g->6	m->1	n->1	r->12	
sta å	r->2	
sta ö	k->1	v->3	
sta, 	a->3	d->2	e->1	f->1	i->1	o->5	s->2	u->1	
sta.)	F->1	
sta.-	 ->1	
sta..	 ->1	
sta.D	e->3	
sta.E	m->1	
sta.H	e->1	
sta.S	j->1	
sta.V	a->1	i->4	
sta: 	I->1	J->1	V->1	u->1	v->1	
sta; 	d->1	v->1	
sta?N	ä->1	
staNä	s->1	
staaf	f->1	
stab 	s->1	
stabe	h->1	
stabi	l->22	
stabu	l->1	
stack	a->1	
stad 	f->2	m->2	o->3	
stad,	 ->1	
stad.	"->1	D->1	H->1	
stade	 ->16	,->1	l->2	s->1	
stadg	a->27	o->1	
stadi	e->4	u->4	
stadk	o->24	
stads	b->1	c->1	o->1	p->1	
stadt	,->1	
stag 	p->1	s->1	
stag,	 ->1	
stag.	I->2	S->1	
staga	n->12	r->40	
stage	n->2	
stagn	a->1	e->1	
stain	s->22	
stak,	 ->1	
staka	 ->5	
stakl	a->1	
stali	n->2	
stall	e->1	k->2	
stalt	e->1	
stamp	 ->1	
stan 	1->3	a->1	b->1	d->1	e->2	f->4	h->1	i->3	k->2	m->1	o->10	p->1	t->2	u->2	v->1	ä->26	ö->3	
stan,	 ->5	
stan.	(->2	A->1	F->1	H->1	J->3	S->1	T->1	U->1	V->3	
stanb	u->1	
stand	a->25	e->16	
stank	a->4	r->1	
stann	a->7	
stans	 ->8	,->4	.->1	?->1	e->6	r->22	
stant	e->1	i->3	
star 	d->2	e->2	f->2	g->1	i->1	j->3	m->6	o->5	p->2	t->1	
stare	 ->2	
stari	n->1	
stark	 ->11	,->1	a->25	e->1	t->23	
start	a->11	e->4	p->1	
stas 	a->1	l->3	v->1	
stas,	 ->1	
stasi	e->1	
stast	r->1	
stat 	-->1	a->1	b->1	d->2	e->3	f->12	g->1	h->6	i->4	l->1	m->3	n->1	o->9	p->1	s->7	t->2	u->2	v->1	å->1	
stat,	 ->7	
stat.	B->1	D->4	G->1	H->1	I->1	J->2	K->1	L->1	O->1	
state	 ->2	n->26	r->335	
stati	o->15	s->8	
statl	i->98	
stats	 ->14	-->5	b->2	k->1	m->4	n->4	p->1	s->19	
statt	a->1	
statu	e->2	s->8	
staur	e->1	
stav 	o->1	
stavl	i->1	
stban	k->4	
stbes	t->1	
stbev	a->1	
stbil	d->1	
stblo	c->1	
stbri	n->1	
stdem	o->11	
ste -	 ->3	
ste E	M->1	k->1	u->6	
ste F	N->1	
ste I	s->1	
ste a	b->1	c->2	g->1	l->11	n->13	r->4	s->1	t->3	v->4	
ste b	e->25	i->1	l->15	y->1	ä->2	ö->5	
ste c	e->1	h->1	
ste d	a->5	e->37	i->1	o->5	r->1	ä->10	å->3	
ste e	k->1	l->1	m->1	n->3	p->1	r->7	u->2	v->1	x->1	
ste f	a->8	e->2	i->7	o->1	r->5	u->1	y->1	å->13	ö->20	
ste g	a->2	e->14	i->1	r->4	å->5	ö->15	
ste h	a->6	e->1	i->1	j->2	o->3	ä->1	å->2	
ste i	 ->9	a->2	f->1	n->23	
ste j	a->8	o->1	u->2	
ste k	a->2	l->1	n->1	o->17	r->6	u->4	ä->2	
ste l	a->1	e->2	i->1	y->1	ä->1	ö->4	
ste m	a->24	e->7	i->2	o->2	å->10	ö->1	
ste n	a->4	e->1	i->2	o->3	u->5	å->2	
ste o	c->28	f->1	l->1	m->1	r->1	
ste p	a->2	e->1	o->1	r->3	u->1	å->6	
ste r	a->1	e->17	i->1	ä->2	å->6	
ste s	a->6	e->15	j->3	k->12	l->1	n->2	o->1	t->15	y->6	ä->14	å->3	ö->4	
ste t	a->26	e->4	i->15	o->1	r->2	y->1	ä->2	
ste u	n->5	p->14	t->17	
ste v	a->31	e->10	i->70	ä->3	
ste ä	g->2	n->7	v->4	
ste å	r->16	t->6	
ste ö	k->2	p->1	v->5	
ste, 	k->1	n->1	v->1	ä->1	
ste.D	e->1	
ste.F	ö->1	
ste.V	i->1	
ste: 	V->1	
stedt	 ->2	,->2	
steen	h->5	
steer	i->1	
stefe	l->1	
stefr	å->1	
stefö	r->5	
steg 	a->1	b->1	f->11	g->1	h->2	i->13	j->1	l->2	m->4	n->2	o->2	p->3	s->7	t->3	u->1	v->1	
steg,	 ->3	
steg.	D->2	
stege	n->5	t->2	
stein	.->1	
stekn	i->1	o->1	
stela	 ->1	,->1	
stele	v->1	
stels	e->5	
stelt	.->1	
stem 	-->1	a->3	d->3	e->1	f->21	g->1	i->5	k->2	m->10	o->7	p->3	s->16	ä->1	ö->1	
stem,	 ->9	
stem.	 ->1	D->3	E->1	G->1	H->2	M->1	T->1	U->1	
stem:	 ->1	
stema	n->5	t->10	
steme	n->12	t->69	
stemä	n->37	
sten 	A->1	I->1	a->4	d->2	f->2	g->1	h->1	i->5	k->1	m->2	o->2	p->6	s->2	t->1	v->1	å->1	
sten"	 ->1	
sten,	 ->12	
sten.	D->2	E->1	H->1	J->1	K->1	O->1	S->1	V->1	
stenN	ä->1	
stena	r->3	
stend	e->1	ö->1	
stene	n->1	
stenk	o->1	
stens	 ->5	,->1	b->1	e->1	
stent	 ->1	
stepr	o->1	
ster 	-->2	B->2	C->1	E->1	F->1	G->6	J->1	S->1	T->1	a->6	b->2	d->3	e->4	f->3	h->2	i->8	k->6	l->2	m->6	o->14	p->4	s->24	t->3	u->2	v->3	ä->4	ö->7	
ster!	J->1	
ster"	 ->1	,->1	
ster,	 ->19	
ster.	.->1	D->5	E->4	F->1	H->2	J->4	K->1	M->1	N->2	O->2	P->1	S->2	T->2	V->2	Ä->1	Å->1	
stera	 ->7	,->1	.->1	d->4	n->3	r->16	s->1	
sterd	a->39	
sterf	a->1	i->2	
steri	l->1	n->16	
sterm	ö->2	
stern	 ->20	,->2	.->9	/->2	a->47	f->1	i->1	s->5	
sterp	o->2	r->1	
sterr	e->3	i->130	å->14	
sters	 ->1	
stes 	i->2	
stese	k->2	
stest	 ->1	
stet 	k->1	
stet.	)->3	
steur	o->9	
stext	e->3	
stfli	r->1	
stful	l->1	
stfäl	l->8	
stför	d->1	k->7	
stgru	p->3	
stgör	 ->1	a->2	
sthan	d->1	
sthom	 ->3	
sthäl	s->1	
sthål	l->1	
stian	 ->1	
stice	 ->4	
stick	 ->1	e->1	p->3	
stid 	k->1	o->1	
stid,	 ->1	
stide	n->5	r->1	
stidn	i->2	
stids	d->3	
stier	,->1	
stift	a->15	n->113	
stig 	s->1	
stiga	 ->2	n->1	s->1	
stige	r->2	
stigh	e->1	
stigi	t->2	
stigl	i->4	
stigm	a->1	
stigt	 ->4	
stik 	p->1	s->2	
stike	n->3	
stil 	-->1	m->1	
still	a->1	d->1	f->34	h->2	s->14	v->5	ä->2	
stimu	l->11	
stina	 ->6	-->1	f->2	s->1	
stind	u->2	
stini	e->4	
stink	t->3	
stinr	i->1	
stins	k->8	
stion	e->1	
stipe	n->1	
stisk	 ->9	.->5	a->57	t->22	
stiti	e->6	
stitu	e->1	t->158	
stjän	s->7	
stjär	n->2	
stkla	s->1	
stkom	p->1	
stkub	i->1	
stkus	t->1	
stkäl	l->1	
stlag	t->1	
stlan	d->2	
stlig	 ->1	
stlin	j->2	
stläg	g->2	
stlän	d->1	
stmak	t->1	
stmar	g->1	
stmyn	d->3	
stmän	g->2	
stnad	 ->10	.->1	;->1	e->74	s->22	
stnar	 ->1	
stnin	g->72	
stnäm	n->2	
sto h	å->1	
sto v	i->1	
stod 	a->3	d->2	e->2	f->1	i->1	j->1	m->1	n->1	p->2	s->1	
stodo	n->1	
stol 	b->1	d->1	i->1	o->1	s->2	v->1	
stol.	D->1	E->1	
stola	r->25	
stole	n->46	
stolk	a->1	
stolp	e->1	
stols	a->1	b->1	f->2	k->1	p->1	s->1	t->1	u->1	v->1	
stolt	 ->6	a->3	h->2	
stomr	å->2	
stone	 ->27	
stop-	s->1	
stopp	 ->8	a->10	m->1	
stor 	a->3	b->16	c->1	d->13	e->3	f->4	g->2	h->5	i->2	j->2	k->3	l->1	m->12	o->3	p->3	r->6	s->1	t->2	u->16	v->4	ö->1	
stor,	 ->1	
stor.	O->1	
stora	 ->151	,->2	.->3	?->1	
stord	r->2	
store	 ->1	r->3	
storf	ö->2	
storh	e->1	
stori	a->10	e->9	k->1	s->16	
stork	a->1	
storm	 ->1	,->1	a->18	e->6	f->1	
stors	k->2	l->2	
stort	 ->41	
stown	 ->2	,->1	
stpar	t->5	
stra 	A->1	E->1	F->1	J->1	T->1	c->1	m->1	o->1	
strad	i->1	
straf	f->40	
strak	t->1	
stram	 ->1	n->2	
stran	d->1	
strar	 ->6	,->3	.->1	:->1	n->5	s->1	
strat	e->63	i->28	
strax	 ->2	
strea	m->8	
strec	k->1	
streg	i->1	
strer	a->12	i->3	
stres	 ->2	
stret	 ->1	
stri 	b->1	d->1	i->1	o->2	s->6	
stri,	 ->3	
stri-	 ->1	
strib	u->1	
stric	h->6	
strid	 ->9	a->2	d->2	e->8	i->1	l->1	
strie	l->6	r->2	
strif	r->4	
strik	t->25	
stril	i->1	o->1	
strin	 ->39	!->1	,->15	.->14	:->1	?->1	g->3	s->9	
strip	o->2	
stris	 ->3	
stroe	n->2	
strof	 ->24	,->4	.->4	a->1	d->1	e->51	h->1	s->4	
stron	o->4	
strot	t->1	
strue	r->5	
struk	i->1	t->185	
strum	e->52	
strun	t->4	
stryk	.->1	a->29	e->2	s->2	
stryp	s->1	
sträc	k->32	
strän	d->2	g->63	
strät	t->3	
sträv	a->30	i->1	
stråe	t->1	
strål	k->1	n->3	s->1	
ströj	o->1	
strök	 ->1	,->1	s->1	
ström	 ->4	,->1	:->1	m->7	n->6	
sts p	u->1	
sts v	i->1	
sts.D	å->1	
sts.S	l->1	
stsam	 ->1	m->1	
stsek	t->2	
stsla	g->2	
stslo	g->2	
stslå	 ->5	r->4	s->8	
ststä	l->51	
stsva	g->1	
stton	e->1	
sttys	k->2	
stu m	e->1	
stude	n->2	r->3	
studi	e->9	
stugo	r->1	
stull	a->1	
stum 	o->1	
stund	 ->8	a->2	e->7	
sturi	e->1	s->1	
stutv	i->2	
stvak	t->1	
stver	k->1	
stvik	t->3	
stvis	t->1	
stvär	l->1	
styck	e->5	
stymp	a->1	n->2	
styr 	a->1	
styra	 ->6	n->4	s->1	
styre	 ->1	,->1	k->3	l->7	t->3	
styrk	a->13	e->2	o->2	
styrn	i->7	
styrs	 ->2	
städa	 ->1	t->1	
städe	r->17	s->2	
ställ	a->136	b->1	d->67	e->104	i->6	n->70	s->20	t->22	
stämd	 ->5	a->8	e->5	h->1	
stämm	a->24	e->158	i->4	
stämn	i->2	
stämp	e->1	l->1	
stäms	 ->1	
stämt	 ->13	,->3	
stän 	e->1	
ständ	i->107	l->1	
stäng	a->2	d->1	e->1	n->6	t->1	
stänk	a->2	e->1	s->1	t->2	
stärk	a->28	e->3	n->6	s->5	t->9	
stäth	e->1	
stäv 	m->1	
stävj	a->1	
stå a	l->1	t->11	v->4	
stå d	e->3	
stå e	n->1	
stå f	o->1	r->8	ö->12	
stå h	u->2	
stå i	 ->4	n->1	
stå k	l->3	v->1	
stå n	y->1	ä->1	
stå o	c->2	m->1	
stå s	o->1	
stå t	i->1	
stå u	t->2	
stå v	a->4	
stå, 	a->1	f->1	s->1	
stå.F	P->1	
stå.J	u->1	
stå: 	å->1	
stådd	 ->1	a->1	
ståel	i->6	s->8	
ståen	d->32	
stålf	ö->5	
stålg	e->1	
ståli	n->25	
ståls	e->4	t->1	
stålv	e->5	
stånd	 ->54	,->8	.->10	?->2	a->5	e->30	i->1	p->97	s->19	
står 	a->25	d->13	e->6	f->20	g->1	h->9	i->44	j->3	k->10	l->2	m->7	n->2	o->2	p->14	s->2	t->4	u->1	v->8	ä->1	å->1	ö->2	
står,	 ->3	
står.	D->2	H->1	
stås 	d->1	f->1	k->1	s->1	u->1	v->1	
stått	 ->27	,->1	.->1	s->1	
stête	 ->1	
stöd 	-->2	a->5	b->1	d->3	e->3	f->26	g->1	h->2	i->11	k->5	l->1	m->4	o->16	p->7	s->19	t->42	v->4	ä->2	å->2	ö->1	
stöd,	 ->14	
stöd.	"->1	.->1	A->1	D->10	E->1	F->2	H->5	I->2	J->2	M->1	N->1	O->1	R->1	S->1	T->1	U->1	V->2	Ä->2	Å->2	
stöd;	 ->1	
stöd?	-->1	
stödd	e->2	
stöde	n->31	r->56	t->32	
stödj	a->71	e->1	
stödm	e->1	o->1	
stödn	i->1	
stödp	o->1	
stödr	a->2	
stöds	 ->8	p->1	y->3	
stödå	t->5	
stöld	,->1	
stör 	b->1	k->1	m->1	s->1	
störa	 ->2	s->3	
störd	a->1	e->2	
störe	l->5	
störi	n->2	
störn	i->5	
störr	e->73	
störs	 ->1	,->1	t->35	
stört	n->1	s->2	
stöta	 ->1	n->1	r->1	
stöte	r->1	s->1	
stötf	å->1	
stött	 ->10	a->2	s->1	
suali	s->1	
subje	k->1	
subsi	d->23	
subst	a->4	
subve	n->10	
succe	s->5	
sudda	 ->1	
suell	 ->1	a->1	
sugar	e->1	
sul o	m->1	
sul s	o->1	
sul.V	i->1	
suler	 ->3	
sulta	t->111	
sultb	a->1	
sulte	r->9	
sum o	c->1	
sumba	r->1	
sumen	t->61	
summa	 ->2	d->1	n->2	t->1	
summe	l->6	
summo	r->8	
sumti	o->2	
sund 	v->1	
sunda	 ->2	,->1	r->1	
sunde	r->3	
sundi	 ->2	:->1	
suner	a->1	
suppe	h->1	
suppf	a->2	ö->1	
suppg	ö->1	
supps	k->1	
supra	n->1	
surd 	i->1	
sursb	r->1	
surse	n->1	r->45	
sursf	ö->1	
surss	l->1	
surst	i->1	
surt 	a->1	m->1	
sus k	a->1	r->1	
sus o	c->1	
susen	 ->1	
suspe	n->1	
sutan	 ->3	
sutbi	l->9	
sutby	t->6	
sutom	 ->59	,->2	
sutru	s->1	
sutry	m->4	
sutsa	t->1	
sutsk	o->2	
sutsl	a->1	
sutsä	t->2	
sutti	t->1	
suttr	y->1	
sutve	c->2	
sutvä	r->1	
sutöv	n->1	
suver	ä->17	
sv. M	e->1	
sv. V	a->1	
sv. m	e->1	
sv., 	ä->1	
sv.?A	n->1	
sv.Sv	e->1	
svag 	i->1	p->1	s->1	
svaga	 ->8	,->2	d->3	r->6	s->7	t->2	
svagh	e->12	
svagn	i->1	
sval,	 ->1	
svans	e->1	i->1	
svar 	-->1	a->6	b->2	d->2	f->26	g->4	h->4	i->7	k->2	m->2	n->2	o->4	p->17	r->1	s->9	t->2	v->2	ä->3	
svar,	 ->26	
svar.	 ->1	D->12	E->1	F->1	G->3	I->1	J->4	M->4	O->1	P->1	S->2	V->4	
svar?	I->1	
svara	 ->30	,->1	.->2	d->10	n->9	r->35	s->2	t->5	
svare	n->3	t->70	
svari	g->56	
svars	.->1	a->1	b->3	f->55	k->4	m->3	o->7	p->5	t->2	
svart	a->2	
svarv	,->1	e->1	
svatt	e->1	n->1	
svek 	h->1	o->1	
svens	k->2	
svent	i->1	
svep 	a->1	
sveps	k->1	
svept	e->1	
sverk	 ->1	a->1	e->1	s->4	
svike	l->4	n->2	t->1	
svikn	a->1	
svilj	a->2	
svill	k->20	
svinn	a->3	e->12	
svins	t->1	
svis 	-->2	e->1	f->1	g->1	h->3	i->1	k->2	o->1	s->6	v->7	
svis,	 ->6	
svis.	J->1	
svunn	i->4	
sväg,	 ->1	
svält	 ->1	s->1	
svämm	a->3	
svämn	i->4	
svänl	i->2	
svärd	 ->2	.->1	a->8	e->3	
sväre	t->1	
svärl	i->6	
svärr	e->4	
svärt	 ->3	,->1	
sväse	n->6	
sväts	k->1	
svävn	a->1	
svåg 	a->1	
svåge	r->1	
svång	r->1	
svår 	a->1	b->1	f->1	p->1	s->1	
svåra	 ->19	,->1	r->5	
svårb	e->2	
svård	s->1	
svåri	g->31	
svårl	ö->2	
svårt	 ->27	,->1	
svårö	v->1	
swage	n->1	
sydda	 ->1	
sydeu	r->1	
sydku	s->1	
sydvä	s->1	
sydös	t->1	
syfta	d->3	r->30	s->3	
syfte	 ->15	.->1	n->6	t->16	
sykol	o->1	
syl g	e->1	
syl o	c->3	
syl, 	f->1	r->1	
syl- 	o->1	
syl.D	e->1	
syl.J	a->1	
syl.V	i->1	
sylbe	s->1	
sylfö	r->2	
sylrä	t->2	
sylsö	k->6	
symbo	l->9	
sympa	t->8	
sympt	o->1	
syn -	 ->1	
syn a	t->1	v->1	
syn g	e->1	
syn i	 ->2	
syn o	c->5	
syn p	å->4	
syn t	i->65	
syn v	a->1	
syn ä	n->1	v->1	
syn, 	m->1	o->1	
syn.A	t->1	
syn.E	t->1	
syn.S	i->1	l->1	
syn; 	d->1	
syna 	h->1	
synas	 ->1	.->2	
synd 	a->1	f->1	g->1	ä->1	
synda	b->2	
synde	r->1	
syndr	o->1	
synen	 ->5	.->1	
syner	g->2	
synes	 ->1	
synli	g->8	
synne	r->52	
synon	y->1	
synpu	n->29	
syns 	s->1	
synst	a->2	
synsä	t->4	
synt 	n->1	v->1	
synt,	 ->1	
synte	s->1	
synvi	n->12	
syra 	a->1	d->1	i->1	
syrie	r->4	
syris	k->4	
sys f	l->1	
sysse	l->103	
syssl	a->6	
syste	m->190	r->1	
säg: 	D->1	
säga 	"->1	-->1	F->1	S->2	a->76	b->1	d->9	e->4	f->4	g->1	h->4	i->5	j->1	k->2	l->2	m->1	n->11	o->6	r->1	s->2	t->8	v->2	ä->2	å->1	
säga,	 ->15	
säga.	J->1	M->1	
säga:	 ->4	
sägan	d->2	
sägar	e->4	
sägas	 ->4	,->1	
sägel	s->8	
säger	 ->63	,->3	.->2	:->5	
sägne	r->1	
sägni	n->1	
sägs 	d->2	e->1	h->1	i->1	
säker	 ->20	,->1	.->1	h->232	l->15	s->24	t->28	
säkra	 ->31	r->4	s->5	
säkri	n->24	
säkt 	f->7	
säkt.	O->1	
säkta	 ->4	
säkte	n->2	r->1	
sälja	 ->2	r->2	s->1	
säljn	i->3	
sälla	n->2	
sälls	k->8	y->2	
sämne	n->2	
sämra	 ->2	d->4	n->1	r->1	s->2	
sämre	 ->5	
sämst	 ->4	a->1	
sända	 ->4	r->2	
sände	 ->2	b->9	
sändn	i->1	
sändr	i->4	
sänka	 ->3	s->2	
sänkn	i->2	
sänkt	s->1	
sär d	e->2	
sär s	o->1	
särar	t->1	
särbe	s->1	
sären	 ->1	d->3	
särki	l->1	
särsk	i->156	
säson	g->1	
säte.	O->1	
sätt 	-->1	H->1	a->31	b->9	e->5	f->11	g->7	h->5	i->6	k->19	l->2	m->2	o->11	p->7	s->36	t->2	u->7	v->7	ä->9	å->2	ö->1	
sätt,	 ->25	
sätt.	 ->1	A->1	B->1	D->13	E->3	F->1	H->5	I->1	J->6	K->1	L->1	M->3	N->2	S->4	V->3	Ä->1	
sätt:	 ->2	
sätt?	A->1	D->1	
sätta	 ->86	!->1	,->2	.->2	n->5	r->2	s->13	
sätte	n->1	r->64	t->23	
sättl	i->1	
sättn	i->211	
sätts	 ->11	,->2	.->1	
så "m	e->1	
så - 	d->1	i->1	
så 19	9->1	
så Eu	r->4	
så Fl	a->1	
så Mo	r->1	
så ab	s->1	
så ak	t->1	
så al	l->7	
så am	b->1	
så an	d->3	l->1	s->3	t->3	v->1	
så ar	b->1	
så at	t->179	
så av	 ->6	g->2	s->2	
så ba	l->1	r->3	
så be	 ->1	f->1	g->1	h->3	k->2	r->4	s->2	t->2	
så bi	d->1	l->1	
så bl	i->5	
så bo	r->3	
så br	a->3	e->2	
så by	g->2	
så bä	r->1	t->1	
så bö	r->4	
så de	 ->10	l->3	m->1	n->2	s->1	t->12	
så di	s->1	
så do	m->1	
så dr	a->1	u->1	
så dä	r->2	
så ef	f->2	t->1	
så ek	o->1	
så en	 ->24	k->1	l->1	
så er	k->1	
så et	t->10	
så fa	k->1	l->2	r->1	s->1	
så fi	n->7	
så fo	r->4	
så fr	a->3	e->1	å->6	
så fu	l->1	n->1	
så få	 ->3	r->4	t->2	
så fö	l->1	r->28	
så ga	r->1	
så ge	 ->2	m->1	n->1	r->1	
så gl	a->1	
så go	d->2	
så gr	a->2	u->1	
så gä	l->1	r->2	
så gå	 ->1	r->2	
så gö	r->5	
så ha	 ->4	n->3	r->6	
så he	l->8	t->1	
så hj	ä->4	
så ho	m->1	p->1	s->1	t->1	
så hu	r->3	
så hä	n->1	r->4	v->1	
så hå	l->1	
så hö	g->1	
så i 	A->1	S->1	T->1	b->1	d->4	e->5	f->2	k->2	l->1	n->1	r->1	s->1	v->2	
så ia	k->1	
så il	l->1	
så im	p->1	
så in	f->1	g->3	l->1	n->2	o->1	r->3	s->3	t->13	v->2	
så ja	g->2	
så ka	d->1	l->10	n->12	
så kl	a->3	
så ko	m->19	n->3	r->4	
så kr	i->4	ä->1	
så ku	n->2	
så kä	n->1	
så kö	r->1	
så li	g->1	s->1	t->3	
så ly	c->1	
så lä	m->1	n->13	t->2	
så lå	g->3	n->9	
så ma	n->1	
så me	d->13	l->1	r->3	
så mi	n->2	s->1	
så mo	t->1	
så my	c->38	
så må	n->15	s->13	t->2	
så mö	j->2	
så no	g->1	t->2	
så ny	s->1	
så nä	m->2	r->3	
så nå	g->4	t->1	
så nö	d->4	
så oa	c->2	
så oc	h->1	
så of	t->4	
så og	y->1	
så om	 ->7	t->1	
så or	s->1	
så pa	r->2	s->2	
så pe	n->1	
så pl	a->1	
så po	s->1	
så på	 ->11	m->2	p->2	v->1	
så ra	n->1	
så re	a->1	d->3	
så ri	k->2	
så rä	c->1	t->1	
så rå	d->1	
så rö	s->2	
så sa	d->1	m->3	n->2	t->1	
så se	 ->6	r->1	s->1	
så si	n->1	
så sj	ä->1	
så sk	a->11	e->3	o->1	u->5	y->1	
så sl	å->1	
så sm	i->1	å->5	
så sn	a->28	
så so	m->22	
så sp	e->1	
så st	a->3	o->8	r->4	ä->2	ö->3	
så sv	å->4	
så sä	g->11	k->5	r->1	t->13	
så så	 ->3	
så ta	 ->8	c->6	l->1	r->1	s->2	
så ti	l->17	
så to	g->1	
så tr	o->4	
så ty	d->1	
så tä	n->1	
så un	d->4	
så up	p->12	
så ut	 ->1	a->2	g->1	o->2	t->1	
så va	d->1	r->15	
så ve	m->1	r->2	t->1	
så vi	 ->4	a->1	c->1	d->10	k->12	l->11	s->2	t->1	
så vä	l->4	
så vå	r->3	
så zi	g->1	
så äg	n->1	
så än	 ->1	d->1	
så är	 ->33	
så åt	e->2	m->1	
så öp	p->1	
så öv	e->3	
så, a	t->2	
så, e	n->1	
så, f	r->1	ö->1	
så, h	e->2	
så, i	 ->2	
så, m	e->1	
så, n	u->1	
så, o	b->1	c->1	m->2	
så, s	o->1	å->1	
så, t	i->1	
så. D	e->1	
så.De	n->1	t->1	
så.I 	s->1	
så.In	t->1	
så.Ja	g->1	
så.Ni	 ->1	
så.Oc	h->1	
så.På	 ->1	
så: a	t->1	
sådan	 ->56	,->2	.->2	?->1	a->48	t->54	
såg a	t->7	
såg d	e->1	ä->1	
såg e	t->1	
såg i	n->1	
såg n	å->1	
såg o	m->1	
såg s	i->1	o->1	
såg u	t->2	
såg Ö	s->1	
sågs 	i->1	m->1	
sågs.	J->1	L->1	
sågve	r->1	
såhär	.->1	
sålde	r->2	
såled	e->40	
sålun	d->4	
sång 	s->1	
sånge	n->1	r->1	
sårba	r->3	
såret	,->1	
såsom	 ->32	
såte 	s->1	
såter	v->1	
såtgä	r->11	
såtgå	n->1	
såtil	l->1	
såvid	a->3	
såväl	 ->40	
sí är	 ->1	
södan	d->1	
söde 	u->1	
södra	 ->6	
sök a	t->4	
sök i	 ->5	
sök o	m->1	
sök s	o->1	
sök, 	o->1	s->1	
söka 	F->1	a->4	b->2	d->1	e->3	f->9	g->2	h->2	i->1	k->1	m->2	o->2	s->2	t->1	u->4	v->3	å->1	
söka,	 ->1	
sökan	d->7	
sökar	l->6	
sökas	 ->2	,->1	.->2	
söken	 ->1	
söker	 ->21	
söket	 ->4	
sökni	n->24	
sökt 	F->1	a->5	b->1	d->1	e->1	f->1	h->1	o->1	u->1	v->1	
sökte	 ->6	
sönde	r->7	
söner	 ->1	
sörja	 ->9	
sörjd	e->1	
sörje	r->2	
sörjn	i->4	
söver	g->1	s->12	t->1	v->1	
sövni	n->1	
t "EU	-->1	
t "Ku	l->2	
t "Kv	i->2	
t "Ol	j->1	
t "Po	r->1	
t "eg	e->1	
t "ek	o->1	
t "en	t->1	
t "eu	r->1	
t "ku	l->1	
t "ob	e->1	
t "re	f->1	s->1	
t (57	1->1	
t (80	9->2	
t (96	1->1	
t (B5	-->2	
t (CE	R->1	
t (EU	G->2	
t (FP	Ö->1	
t (IC	E->1	
t (IF	O->1	
t (SP	Ö->1	
t (ar	t->1	
t (de	 ->1	
t (fi	s->2	
t (hä	l->1	
t (i 	s->1	
t (in	r->1	
t (ko	n->1	
t (t.	e->1	
t (ty	v->1	
t (ÖV	P->1	
t , d	e->1	
t - a	l->2	t->2	v->3	
t - d	e->5	v->1	å->1	
t - e	l->1	n->2	t->1	v->1	
t - f	a->1	å->1	ö->4	
t - g	e->1	ö->1	
t - h	a->1	o->1	
t - i	 ->4	n->1	
t - j	a->4	
t - k	n->1	o->3	
t - m	e->2	o->1	
t - n	ä->2	å->1	
t - o	c->10	m->1	r->1	
t - p	r->1	
t - s	n->1	o->4	t->1	ä->2	å->3	
t - t	i->1	
t - u	t->1	
t - v	i->9	
t - ä	r->1	v->1	
t - å	t->2	
t - ö	p->1	v->1	
t -, 	m->1	u->1	
t -er	 ->1	
t 1 0	0->1	
t 1 u	t->1	
t 1, 	s->1	
t 10 	0->1	å->1	
t 11 	i->1	
t 12 	p->1	
t 13 	0->1	
t 180	 ->1	
t 194	8->1	
t 199	4->1	7->10	8->2	9->5	
t 2 i	 ->2	
t 200	1->1	
t 21:	a->1	
t 22 	r->1	
t 23,	7->1	
t 25 	p->2	
t 26 	"->1	
t 27 	f->1	
t 3 p	r->1	u->1	
t 39 	p->1	
t 4 i	 ->1	
t 4 l	i->1	
t 40 	p->1	
t 400	 ->2	
t 48 	ä->1	
t 5 0	0->1	
t 5, 	o->1	
t 5,5	 ->1	
t 50-	t->1	
t 6 o	m->1	
t 7 i	 ->1	
t 70 	p->1	
t 700	 ->2	
t 8 r	e->1	
t 80 	p->1	
t 88/	5->2	
t 9 f	a->1	
t 90 	d->1	
t 93 	p->1	
t 94/	7->1	
t 95 	m->1	
t 98 	m->1	
t : P	a->1	
t ABB	-->1	
t Ado	l->1	
t Aid	s->1	
t Akk	u->1	
t Ale	x->1	
t Alt	e->3	
t Ams	t->3	
t Ass	a->1	
t Aus	c->1	
t BNP	 ->1	
t Bar	a->1	n->1	ó->1	
t Ber	e->1	n->1	
t Bou	r->1	
t Bre	t->1	
t Bro	k->1	
t Bry	s->1	
t CEN	,->1	
t Cam	u->1	
t Cas	a->1	
t Cli	n->1	
t D k	r->1	
t Dal	a->2	
t Dan	m->4	
t De 	t->1	
t Dub	l->1	
t Dui	s->1	
t EG-	d->3	k->6	r->1	
t EG:	s->2	
t EIF	 ->1	
t EKS	G->1	
t ELD	R->1	
t EU 	a->1	b->1	p->1	r->1	s->2	u->1	ä->1	
t EU-	i->1	l->1	s->2	
t EU.	.->1	D->1	V->1	
t EU:	s->7	
t Ell	e->1	
t Equ	a->7	q->1	
t Eri	k->3	
t Eur	o->111	
t Eva	n->1	
t FEO	 ->1	
t FN-	u->1	
t FN:	s->1	
t FPÖ	 ->3	
t Flo	r->4	
t Fra	n->3	
t För	 ->1	e->4	
t Gar	g->1	
t Goe	b->1	
t Gre	k->3	
t Gru	p->1	
t Grö	n->1	
t Had	e->1	
t Hai	d->3	
t Heb	r->1	
t I T	u->1	
t ICE	S->1	
t INT	E->1	
t Int	e->2	
t Irl	a->1	
t Isr	a->4	
t Ita	l->3	
t Jon	c->3	
t Jör	g->3	
t Kar	a->1	
t Kir	g->1	
t Kos	o->2	
t Kou	c->2	
t Kul	t->3	
t Kyo	t->2	
t Lan	g->1	
t Lea	d->2	
t Mal	t->1	
t Mar	p->1	
t Mid	l->1	
t Min	i->1	
t Mon	t->1	
t Mor	a->1	b->1	g->1	
t Mün	c->1	
t Nat	o->1	
t OLA	F->3	
t Pat	t->1	
t Pet	e->1	
t Por	t->6	
t RIN	A->2	
t Ran	d->2	
t Rap	k->3	
t Rot	h->1	
t SEM	-->1	
t San	t->1	
t Sav	e->1	
t Sch	r->1	
t Sju	k->1	
t Sjö	s->1	
t Sok	r->1	
t Sou	l->1	
t Sto	r->3	
t Sud	r->1	
t Sve	r->1	
t TV-	k->1	
t The	a->3	
t Tib	e->1	
t Tod	i->1	
t Tot	a->2	
t Tur	k->14	
t UNM	I->1	
t Vat	a->1	
t Ver	s->1	
t Vod	a->1	
t Vär	l->1	
t Waf	f->1	
t Wal	l->1	
t Wul	f->1	
t abs	o->6	t->1	u->1	
t acc	e->12	
t ad 	h->1	
t add	i->1	
t ade	k->3	
t adm	i->2	
t age	r->16	
t aid	s->1	
t akt	a->1	e->1	i->8	u->7	
t aku	t->1	
t alb	a->1	
t ald	r->3	
t ali	b->1	
t all	 ->5	a->37	d->1	e->3	i->1	m->14	r->1	t->30	v->20	
t alt	e->2	
t amb	i->3	
t ame	r->3	
t ana	 ->1	l->9	
t and	e->1	r->62	
t anf	ö->5	
t ang	e->8	r->7	å->1	
t anl	e->2	i->1	
t anm	ä->2	
t ann	a->30	o->2	
t ano	r->2	
t anp	a->2	
t ans	e->10	j->2	l->6	t->8	v->66	å->2	ö->1	
t ant	a->61	i->1	o->8	
t anv	ä->31	
t ara	b->1	
t arb	e->102	
t arg	u->1	
t arr	a->2	e->1	
t art	i->15	
t arv	.->1	
t asy	l->3	
t att	 ->813	e->3	
t av 	"->1	-->1	1->3	A->1	B->3	D->1	E->23	I->1	J->1	K->3	M->1	P->1	T->1	V->2	a->35	b->11	c->1	d->119	e->60	f->48	g->9	h->5	i->6	j->1	k->14	l->7	m->17	n->7	o->9	p->16	r->18	s->20	t->6	u->7	v->18	ä->1	å->5	ö->2	
t ava	n->1	
t avb	r->2	
t avd	e->1	
t avf	a->4	
t avg	e->1	j->1	r->2	ö->11	
t avh	j->2	å->1	
t avl	ä->4	
t avs	e->22	i->1	k->13	l->11	t->10	ä->3	
t avt	a->17	v->1	
t avv	e->3	i->3	
t bad	 ->1	
t bak	 ->1	g->17	o->3	å->2	
t bal	a->1	
t ban	a->2	
t bar	a->18	n->2	
t bas	k->1	
t bax	a->1	
t be 	e->1	k->1	o->1	
t bea	k->10	
t bed	r->7	ö->4	
t bef	i->4	o->2	r->3	ä->6	
t beg	r->17	ä->9	å->3	
t beh	a->11	o->8	å->2	ö->26	
t bek	l->5	o->1	r->7	v->1	y->6	ä->24	
t bel	a->1	g->1	o->3	ä->2	
t bem	ö->4	
t ben	å->1	
t ber	 ->2	e->2	i->2	o->16	ä->5	ö->9	
t bes	i->1	k->7	l->42	t->23	v->9	ö->1	
t bet	a->10	o->10	r->14	y->21	ä->59	
t bev	a->12	i->23	
t bib	e->3	
t bid	r->24	
t bif	a->1	
t big	o->1	
t bil	a->3	d->8	i->3	l->2	m->1	t->3	v->1	ä->1	
t bin	d->7	
t bio	l->1	
t bis	t->9	
t bit	t->1	
t bl.	a->2	
t bla	n->6	
t ble	v->1	
t bli	 ->45	.->1	c->1	n->1	r->22	v->3	
t blu	n->1	
t bly	,->1	g->2	
t bo 	i->1	
t bog	s->1	
t bom	b->1	
t bor	d->12	t->5	
t bos	t->1	ä->1	
t bot	t->1	
t bra	 ->31	.->1	
t bre	t->5	v->5	
t bri	e->1	n->1	s->4	t->5	
t bro	k->1	m->4	t->4	
t bry	t->8	
t brä	n->2	
t brå	d->4	
t bud	g->7	s->4	
t byg	g->18	
t byr	å->3	
t bär	a->1	
t bäs	t->7	
t bät	t->22	
t båd	a->2	e->5	
t båt	a->1	
t bör	 ->34	j->26	
t cas	e->1	
t cem	e->2	
t cen	t->5	
t cha	n->2	
t cir	k->1	
t cit	e->1	
t civ	i->6	
t d) 	i->1	
t dag	e->1	o->6	s->3	
t dan	s->8	
t dat	u->9	
t de 	a->11	b->7	d->3	e->10	f->17	g->3	h->8	i->14	j->1	k->21	l->9	m->10	n->9	o->11	p->16	r->4	s->43	t->9	u->7	v->7	y->1	ä->10	å->4	ö->1	
t de,	 ->1	
t deb	a->11	
t dec	e->2	
t def	i->7	
t del	 ->3	a->12	e->2	t->8	
t dem	 ->9	,->1	.->1	o->16	
t den	 ->216	,->1	.->3	;->1	n->71	
t dep	a->1	
t der	a->5	
t des	s->50	
t det	 ->524	,->5	.->6	a->5	s->1	t->143	
t dia	l->1	
t dil	e->2	
t dip	l->1	
t dir	e->40	
t dis	c->2	k->36	
t div	e->1	
t dju	p->2	r->1	
t djä	r->3	v->1	
t doc	k->4	
t dok	u->11	
t dol	l->2	
t dom	a->1	e->1	i->1	s->7	
t dra	 ->14	b->9	g->1	m->2	r->2	s->2	
t dri	v->9	
t drå	p->1	
t drö	j->3	
t dub	b->2	
t dyk	a->1	
t dyn	a->2	
t dyr	a->2	t->1	
t däm	p->2	
t där	 ->23	,->1	.->2	f->9	i->3	m->3	v->1	
t då 	d->3	e->1	f->2	i->1	k->2	m->1	s->1	t->1	v->1	
t dål	i->5	
t dö 	i->1	
t död	a->2	
t döl	j->3	
t döm	a->6	
t dör	 ->1	
t e) 	i->1	
t e-m	a->1	
t ede	n->1	
t eff	e->20	
t eft	e->42	
t ege	n->12	t->19	
t egn	a->4	
t eko	l->2	n->22	
t el-	 ->1	
t ele	k->2	m->1	
t eli	m->1	
t ell	e->38	
t emb	a->1	
t eme	l->3	
t emo	t->5	
t en 	a->16	b->12	c->2	d->10	e->17	f->13	g->6	h->5	i->2	k->11	l->6	m->16	n->4	o->14	p->9	r->15	s->23	t->11	u->4	v->8	ä->2	å->2	ö->7	
t ena	 ->10	s->3	
t enb	a->5	
t end	a->28	
t ene	r->3	
t eng	a->8	
t enh	e->10	ä->6	
t eni	g->2	
t enk	e->25	l->5	
t enl	i->8	
t eno	r->6	
t ens	 ->2	a->1	k->1	
t ent	r->1	u->1	
t env	e->1	
t epo	k->1	
t er 	i->2	n->1	o->1	p->1	s->1	t->1	u->2	
t er,	 ->1	
t era	 ->4	
t erb	j->4	
t erf	a->3	o->1	
t erh	å->2	
t eri	n->3	
t erk	ä->13	
t ers	ä->6	
t ert	 ->7	
t eta	b->5	
t ett	 ->117	:->1	
t eur	o->48	
t eve	n->5	
t ex 	a->1	t->1	
t exa	k->6	m->1	
t exc	e->2	
t exe	m->30	
t exi	s->1	
t exp	a->3	e->6	
t ext	r->7	
t f.d	.->1	
t fai	l->1	
t fak	t->65	
t fal	l->34	
t fan	n->8	t->4	
t far	a->2	l->5	t->4	
t fas	c->1	t->27	
t fat	t->13	
t fed	e->1	
t fel	 ->4	,->1	.->2	a->4	
t fem	:->1	p->1	t->11	å->1	
t fen	o->1	
t fic	k->4	
t fin	a->17	l->4	n->198	s->2	
t fis	k->4	
t fjä	r->4	
t fle	r->21	x->6	
t fly	g->3	t->4	
t fod	e->1	
t fog	 ->1	
t fok	u->2	
t fol	k->7	
t fon	d->1	
t for	d->6	m->11	s->3	t->34	u->2	
t fot	f->1	
t fra	m->98	n->6	
t fre	d->11	
t fri	 ->1	a->2	g->2	h->9	t->1	
t fru	k->2	s->2	
t fry	s->1	
t frä	m->42	
t frå	g->24	n->97	
t ful	l->19	t->1	
t fun	d->1	g->14	k->1	n->1	
t fyl	l->1	
t fyr	a->2	
t fys	i->1	
t fän	g->1	
t fäs	t->2	
t få 	1->1	G->1	a->3	b->3	d->9	e->19	f->6	i->6	k->1	l->3	m->2	n->1	o->1	p->4	r->4	s->17	t->14	u->2	v->2	å->1	
t få.	E->1	G->1	
t fåg	e->1	l->2	
t får	 ->25	?->1	
t fåt	a->1	t->2	
t föd	s->1	
t föl	j->14	
t för	 ->603	,->1	?->1	a->13	b->60	d->30	e->96	f->32	g->1	h->30	i->1	k->15	l->10	m->9	n->9	o->8	r->4	s->236	t->19	u->9	v->23	ä->14	ö->2	
t gam	l->4	
t gan	s->4	
t gar	a->20	d->1	
t gav	 ->1	,->1	s->1	
t ge 	F->1	a->4	b->4	d->1	e->9	f->1	h->3	k->1	m->2	n->1	o->5	p->4	r->4	s->5	t->2	u->6	v->2	
t ge.	J->1	
t gem	e->43	
t gen	a->3	d->1	e->8	o->78	s->1	t->4	
t geo	g->2	
t ger	 ->11	,->1	
t ges	 ->1	
t get	t->2	
t gic	k->2	
t gil	t->1	
t giv	a->2	e->2	i->1	
t gjo	r->7	
t gla	d->6	
t glo	b->3	
t glä	d->11	
t god	 ->1	a->6	k->34	s->34	t->7	
t got	t->13	
t gra	n->15	t->8	v->1	
t gre	p->2	
t gri	p->4	
t gru	n->15	
t grä	l->2	
t grö	n->2	
t gyn	n->6	
t gäl	l->223	
t gär	n->1	
t gå 	e->1	f->3	g->2	h->1	i->10	l->1	m->2	o->1	s->2	t->3	u->2	v->2	
t gå.	O->1	
t går	 ->14	
t gåt	t->3	
t gör	 ->22	a->117	s->2	
t ha 	a->2	b->2	d->4	e->10	f->3	h->1	i->1	k->2	l->4	m->4	n->3	o->1	p->1	s->6	t->2	u->1	v->6	å->1	ö->1	
t ha,	 ->1	
t had	e->9	
t haf	t->4	
t hal	v->4	
t ham	n->3	
t han	 ->50	,->2	d->66	s->4	t->8	
t har	 ->205	,->3	
t hed	e->1	
t hel	a->8	h->1	l->3	s->1	t->14	
t hem	 ->2	.->1	l->5	
t hen	n->1	
t her	r->1	
t hes	 ->1	
t hin	d->10	n->1	
t his	t->4	
t hit	t->10	
t hjä	l->18	r->2	
t hon	 ->7	o->1	
t hop	p->7	
t hor	i->1	m->1	
t hos	 ->11	p->1	
t hot	 ->7	a->2	
t hug	g->3	
t hum	a->1	ö->1	
t hun	d->2	
t hur	 ->18	
t hus	 ->1	,->1	.->1	
t huv	u->3	
t hyc	k->2	
t hys	a->1	
t häl	s->1	
t hän	d->10	g->2	s->12	t->1	v->7	
t här	 ->62	,->1	.->2	i->2	v->1	
t häv	a->1	d->1	
t hål	 ->1	,->1	l->31	
t hån	 ->1	
t hår	d->4	t->3	
t hög	 ->5	a->3	e->1	r->3	s->3	t->8	
t höj	a->2	t->1	
t höl	l->2	
t hör	 ->9	a->11	d->1	n->3	
t i 2	0->1	
t i A	d->1	m->1	s->1	
t i B	e->3	i->1	r->1	u->1	
t i C	E->1	
t i D	u->2	
t i E	M->1	u->12	
t i F	e->1	r->4	ö->3	
t i G	a->1	
t i H	e->9	
t i I	r->2	s->1	t->2	
t i K	i->1	o->3	ä->1	
t i L	i->1	
t i M	a->1	e->2	i->1	
t i N	e->2	
t i P	e->1	o->3	
t i S	a->1	t->1	
t i T	a->8	
t i a	k->2	l->8	n->5	r->6	t->2	
t i b	e->6	i->2	r->1	ö->1	
t i d	a->17	e->67	i->6	o->1	
t i e	f->1	n->17	r->2	t->3	u->1	x->1	
t i f	a->1	e->2	o->3	r->23	u->1	y->1	ö->20	
t i g	e->5	o->3	r->1	å->2	
t i h	a->5	e->4	ä->1	ö->5	
t i j	u->2	ä->1	
t i k	a->3	o->6	r->5	u->1	
t i l	a->1	i->3	j->1	ä->1	
t i m	a->2	e->2	i->7	o->6	å->1	
t i n	o->1	ä->1	å->3	
t i o	c->5	f->1	l->1	m->1	r->2	
t i p	a->7	r->4	
t i r	a->1	e->2	i->1	ä->1	å->8	
t i s	a->15	e->1	i->26	j->3	l->4	n->1	o->2	t->9	y->2	å->1	ö->1	
t i t	i->7	o->1	r->1	
t i u	n->3	t->4	
t i v	a->2	e->2	i->9	ä->4	å->9	
t i Ö	s->4	
t i ä	m->1	n->1	
t i å	r->1	t->2	
t i ö	s->1	v->1	
t i.D	e->1	
t iak	t->1	
t ibl	a->6	
t ick	e->4	
t ide	a->1	n->4	o->1	
t idé	e->1	n->2	
t ifr	å->15	
t ige	n->9	
t igå	n->1	
t ill	a->1	e->1	
t ils	k->2	
t imm	i->3	
t imp	o->3	
t in 	f->1	i->3	m->1	p->3	s->1	
t inb	e->1	j->2	l->3	y->1	
t inc	i->2	
t ind	i->1	
t inf	e->1	i->1	l->7	o->14	r->1	ö->35	
t ing	a->3	e->18	r->8	å->2	
t inh	ä->1	
t ini	t->21	
t ink	l->1	
t inl	e->14	ä->2	å->1	
t inn	a->3	e->56	
t ino	m->46	
t inr	e->1	i->5	ä->22	
t ins	e->3	i->2	k->1	l->1	p->1	t->41	
t int	a->2	e->252	i->1	r->35	
t inv	a->1	e->3	o->2	ä->2	å->1	
t irl	ä->3	
t iro	n->1	
t irr	a->1	i->3	
t iso	l->4	
t ita	l->4	
t ja 	-->1	t->2	
t jag	 ->105	
t jap	a->1	
t job	b->1	
t jor	d->5	
t ju 	a->1	f->1	i->2	m->1	ä->2	
t jun	g->1	
t jur	i->7	
t jus	t->13	
t jäm	f->2	k->1	n->1	s->4	
t jär	n->1	
t kal	l->2	
t kam	m->4	p->2	
t kan	 ->98	,->1	d->1	s->8	
t kao	s->1	
t kap	i->6	
t kas	t->1	
t kat	a->1	
t kem	i->1	
t kla	g->3	r->43	s->6	u->1	
t klo	k->2	
t kly	f->1	
t kna	p->1	
t knu	s->1	
t kny	t->4	
t knä	c->1	
t koa	l->2	
t kol	l->9	
t kom	 ->4	m->310	p->23	
t kon	c->4	f->3	k->24	s->38	t->18	v->5	
t kop	i->1	
t kor	r->11	t->26	
t kos	t->14	
t kra	f->9	s->1	v->9	
t kri	g->4	m->1	n->2	s->1	t->13	
t kro	m->1	
t krä	n->2	v->50	
t kul	l->1	t->17	
t kun	d->7	n->60	s->1	
t kus	t->1	
t kva	l->9	n->1	r->5	
t kvi	n->4	
t kvä	v->2	
t kyl	i->1	
t käm	p->1	
t kän	d->1	n->5	s->11	t->1	
t kär	a->1	n->6	
t köl	 ->1	,->1	d->1	
t kön	s->1	
t köp	k->1	
t köt	t->2	
t lab	o->1	
t lad	e->2	
t lag	d->1	f->2	s->14	
t lan	d->54	t->1	
t lap	p->3	
t las	t->1	
t law	,->1	
t led	 ->1	a->23	e->3	
t leg	a->1	i->2	
t lek	t->1	
t lev	a->5	e->4	
t lib	e->1	
t lid	a->1	e->1	
t lig	g->15	
t lik	a->5	n->4	r->1	s->1	
t lil	l->4	
t lin	d->3	
t lis	t->1	
t lit	e->15	t->2	
t liv	 ->4	s->7	
t lju	s->2	
t lob	b->1	
t loc	k->1	
t log	i->4	
t loj	a->2	
t lok	a->1	
t lot	t->3	
t lov	a->1	
t lud	d->2	
t luf	t->1	
t lug	n->2	
t lut	a->1	h->1	
t lyc	k->12	
t lyd	a->1	
t lyf	t->2	
t lys	a->3	s->5	
t läg	e->7	g->58	l->1	r->2	
t läm	n->11	p->10	
t län	d->2	g->15	k->1	
t lär	 ->1	a->3	d->1	
t läs	t->1	
t lät	t->8	
t läx	a->1	
t låg	a->2	t->1	
t lån	g->13	
t låt	a->12	e->1	
t löf	t->2	
t lön	s->1	
t löp	a->5	e->2	t->1	
t lös	a->18	n->1	r->1	t->1	
t maj	o->4	
t mak	r->2	
t man	 ->206	,->6	a->1	d->4	t->1	
t mar	i->2	k->21	
t mas	s->2	
t mat	e->7	n->1	
t max	i->2	
t med	 ->268	,->1	a->3	b->16	d->17	e->4	f->2	g->5	l->23	v->11	
t mek	a->1	
t mel	l->39	
t men	 ->13	a->2	i->1	
t mer	 ->32	,->1	a->1	v->2	
t mes	t->7	
t met	o->1	
t mig	 ->71	.->1	
t mil	d->2	j->10	l->2	
t min	 ->37	a->2	d->1	i->12	n->5	o->2	s->26	u->3	
t mir	a->1	
t mis	s->16	
t mit	t->5	
t mix	.->1	
t mob	i->2	
t mod	 ->3	e->7	i->2	
t mog	e->1	
t mon	o->2	s->1	
t mor	d->1	
t mot	 ->45	a->1	i->6	o->1	s->12	t->2	v->4	
t mul	t->3	
t mun	t->2	
t mus	i->1	
t myc	k->89	
t myn	d->11	n->1	
t myt	i->1	
t män	g->1	n->10	
t mär	k->6	
t mät	a->1	
t måh	ä->1	
t mål	 ->16	,->1	e->7	i->3	
t mån	 ->1	a->2	g->17	
t mås	t->106	
t måt	t->1	
t möd	o->1	
t möj	l->47	
t mör	k->1	
t möt	a->3	e->5	
t nam	n->2	
t nar	k->2	
t nat	i->8	u->8	
t naz	i->2	
t ned	 ->7	e->1	l->1	s->1	
t neg	a->5	
t nek	a->1	
t ner	 ->3	
t ni 	a->3	b->4	d->2	e->1	f->3	h->6	i->4	j->1	k->4	l->1	n->2	o->1	p->2	r->1	s->8	t->2	u->2	v->1	ä->2	ö->1	
t ni,	 ->2	
t nio	 ->2	
t niv	å->3	
t nog	 ->7	,->1	.->1	a->6	g->5	
t nom	i->1	
t nor	d->4	m->2	
t not	e->3	
t nr 	1->1	
t nu 	3->1	b->2	e->1	f->5	g->6	h->1	i->2	k->1	n->3	o->1	p->1	r->1	s->4	ä->7	
t nu,	 ->3	
t nu.	.->1	V->1	
t num	e->1	
t nuv	a->10	
t ny 	k->1	
t nya	 ->23	
t nyb	i->1	
t nyd	a->1	
t nyk	t->2	
t nyl	i->5	
t nyn	a->1	
t nys	k->1	
t nyt	t->27	
t nyv	a->1	
t näm	n->6	
t när	 ->61	a->3	m->6	v->2	
t näs	t->8	
t nät	v->2	
t nå 	a->1	d->1	e->5	f->2	v->1	
t nåd	 ->1	
t någ	o->34	r->24	
t når	 ->1	
t nöd	v->29	
t nöj	a->1	d->2	e->1	
t nöt	k->1	s->1	
t oac	c->12	
t oav	s->1	
t obe	b->1	g->1	r->6	
t obs	e->1	
t och	 ->665	,->1	
t ock	s->58	
t odj	u->1	
t oef	t->1	
t oeg	e->1	
t oen	s->1	
t oer	h->2	
t off	e->16	
t oft	a->7	
t ofö	r->4	
t ogr	u->2	
t okl	a->2	
t okr	i->1	
t oku	n->1	
t ola	g->1	
t oli	k->2	
t olj	a->1	e->6	
t oly	c->6	
t olä	m->1	
t om 	1->1	E->7	G->1	a->31	b->3	d->42	e->19	f->5	g->1	h->9	i->7	k->12	l->1	m->14	n->2	o->3	p->2	r->9	s->12	t->5	u->11	v->20	Ö->1	ä->3	å->4	
t om,	 ->1	
t om.	A->1	D->2	E->1	J->1	
t omb	e->2	
t omd	ö->2	
t ome	d->5	
t omf	a->17	
t omh	u->1	
t omk	r->3	
t omo	r->2	
t omp	r->1	
t omr	å->42	ö->2	
t oms	t->3	ä->3	
t omv	a->1	ä->2	
t omö	j->5	
t ond	a->2	
t ont	 ->1	
t onö	d->3	
t opa	r->1	
t ope	r->2	
t opp	o->1	
t opr	a->1	o->1	
t opt	i->2	
t ord	 ->7	e->6	f->9	n->1	r->2	
t ore	a->1	d->1	
t org	a->10	
t ori	k->1	m->2	
t oro	a->11	l->2	n->1	s->1	
t ors	a->2	
t orw	e->1	
t orä	k->1	t->1	
t osa	n->1	
t oss	 ->48	,->1	?->1	
t osv	.->2	
t osy	n->1	
t osä	k->1	
t oti	l->5	
t oty	d->2	
t otä	n->1	
t ovä	l->1	s->1	
t oän	d->1	
t oöv	e->2	
t pak	e->1	
t pal	e->1	
t pap	p->1	
t par	 ->16	a->1	k->2	l->57	t->23	
t pas	s->5	
t pat	e->1	
t pea	n->1	
t pek	a->3	
t pen	g->9	s->1	
t per	 ->7	f->2	i->1	m->2	s->15	
t pes	t->2	
t pil	o->1	
t pla	c->6	n->14	s->1	t->2	
t plö	t->1	
t pol	i->39	
t pop	u->2	
t por	t->61	
t pos	i->29	
t pot	e->1	
t poä	n->3	
t pra	k->9	t->2	
t pre	c->4	j->2	m->2	r->1	s->5	
t pri	n->12	o->3	s->7	v->4	
t pro	b->32	c->3	d->9	f->1	g->21	j->11	n->1	t->5	v->6	
t prä	g->1	
t prö	v->2	
t pun	k->5	
t på 	1->1	2->1	3->1	5->1	A->1	B->1	C->1	E->2	I->5	a->29	b->5	d->42	e->38	f->34	g->14	h->1	i->7	k->7	l->2	m->11	n->4	o->8	p->6	r->11	s->17	t->7	u->1	v->14	ä->2	å->1	ö->1	
t på,	 ->3	
t på.	E->1	J->1	
t på:	 ->1	
t på?	J->1	
t påb	ö->3	
t påd	r->1	
t påg	i->2	å->3	
t påm	i->5	
t påp	e->8	
t pås	k->2	t->6	
t påt	a->1	v->2	
t påv	e->10	
t rad	e->1	i->2	
t rak	 ->1	r->1	t->2	
t ram	e->1	p->1	
t ran	d->1	
t rap	p->2	
t ras	h->1	i->1	
t rat	i->4	
t rea	g->4	
t red	a->16	o->1	s->1	
t ree	l->1	
t ref	l->4	o->15	
t reg	e->29	i->12	l->7	
t rek	l->2	o->3	
t rel	a->2	e->1	
t ren	s->3	t->4	
t rep	a->4	r->4	
t res	a->1	o->7	p->10	t->1	u->30	
t ret	r->6	
t rev	i->4	
t rid	a->1	
t rik	a->1	e->1	t->31	
t rim	l->7	
t rin	g->3	
t ris	,->1	k->5	
t ro 	i->1	
t rop	a->1	
t rub	b->1	
t rul	l->1	
t rum	 ->8	,->1	.->1	
t rut	t->1	
t ryk	t->4	
t räc	k->14	
t räd	d->4	s->1	
t räk	n->1	
t rät	t->47	
t råd	 ->2	a->2	e->42	f->3	g->1	s->2	
t råk	a->1	
t rör	 ->12	a->6	i->1	
t rös	t->38	
t röt	t->1	
t s.k	.->1	
t sad	e->7	
t sag	t->9	
t sak	 ->1	e->1	l->1	n->13	o->1	p->1	
t sal	u->1	
t sam	a->25	b->3	f->2	h->12	l->7	m->36	o->5	r->2	t->15	
t san	k->1	n->3	t->3	
t sat	s->3	t->2	
t se 	a->4	d->3	h->2	n->1	o->2	p->4	s->2	t->28	u->1	v->4	ä->1	ö->6	
t sed	a->11	
t seg	d->1	l->6	
t sek	e->1	r->1	t->1	
t sem	e->1	i->1	
t sen	a->15	f->1	t->2	
t ser	 ->8	b->4	i->3	v->1	
t ses	 ->1	
t set	t->27	
t sex	 ->5	
t sid	a->2	
t sif	f->1	
t sig	 ->60	,->2	.->3	n->1	
t sik	t->5	
t sin	 ->13	a->4	e->1	n->3	s->1	
t sis	t->7	
t sit	t->11	u->4	
t sju	 ->1	k->2	n->4	t->1	
t sjä	l->19	t->2	
t sjö	n->1	
t ska	 ->1	d->10	f->3	k->1	l->78	p->86	r->1	t->1	
t ske	 ->5	!->1	d->1	p->4	r->11	t->3	
t ski	c->5	l->5	n->1	p->1	
t skj	u->6	
t sko	g->1	l->1	
t skr	a->1	i->6	o->5	
t sku	l->97	
t sky	d->34	f->1	n->4	
t skä	l->10	m->1	r->4	
t skö	t->3	
t sla	g->9	
t sli	t->1	
t slu	k->1	t->21	
t slä	c->2	p->3	
t slå	 ->4	e->1	r->1	s->1	
t slö	s->2	
t smi	t->1	
t smä	r->1	
t små	 ->1	.->1	
t sna	b->17	r->3	
t snö	v->1	
t soc	i->20	
t sol	a->1	d->1	i->2	
t som	 ->515	,->2	
t sor	g->2	
t spa	n->4	r->4	
t spe	c->10	g->1	k->4	l->12	t->1	
t spo	n->1	t->1	
t spr	i->3	å->1	
t spå	r->2	
t spö	k->1	
t sta	b->2	d->4	g->1	n->4	r->25	t->21	
t ste	g->19	
t sti	f->1	g->2	m->2	
t sto	d->1	l->1	p->4	r->62	
t str	a->11	i->5	u->6	y->1	ä->8	
t stu	d->1	
t sty	c->1	m->1	r->7	
t stä	l->25	m->8	n->4	r->10	
t stå	 ->6	e->1	l->1	n->2	r->26	
t stö	d->135	r->25	t->3	
t sub	s->3	v->1	
t suc	c->1	
t sud	d->1	
t sun	d->1	
t suv	e->2	
t sva	g->5	r->30	
t sve	k->1	p->1	
t svå	r->19	
t syf	t->15	
t sym	p->3	
t syn	a->1	d->2	l->2	n->1	s->1	
t syr	i->1	
t sys	s->2	t->44	
t säg	a->36	e->6	s->1	
t säk	e->33	r->7	
t säl	j->1	
t säm	r->2	
t sän	d->3	k->4	
t sär	s->14	
t sät	e->1	t->175	
t så 	a->16	b->2	e->1	f->4	h->3	i->3	k->4	l->3	m->6	n->1	o->1	s->16	t->2	v->2	ä->2	
t så,	 ->1	
t så.	 ->1	D->1	
t såd	a->49	
t såg	 ->1	
t sål	e->3	
t sås	o->2	
t såv	ä->6	
t söd	r->1	
t sök	a->2	e->2	
t sör	j->2	
t t.o	.->1	
t ta 	A->1	a->3	b->2	d->8	e->7	f->6	g->1	h->12	i->11	l->1	m->3	o->2	p->1	s->6	t->4	u->24	v->2	ö->1	
t ta.	J->1	
t ta?	D->1	
t tab	u->1	
t tac	k->38	
t tag	 ->2	e->5	i->2	n->1	
t tak	 ->1	
t tal	a->24	
t tan	k->5	
t tap	p->1	
t tar	 ->10	
t tas	 ->5	
t tec	k->5	
t tek	n->2	
t tem	p->1	
t teo	r->1	
t ter	r->3	
t tex	t->2	
t the	 ->1	
t tib	e->1	
t tid	 ->4	,->1	e->2	i->15	p->1	s->8	t->1	
t til	l->368	
t tio	 ->1	
t tit	t->5	
t tju	g->1	
t tjä	n->4	
t tog	 ->1	
t tol	e->2	k->4	
t tom	r->2	
t ton	å->1	
t top	p->1	
t tor	v->1	
t tot	a->5	
t tra	d->2	g->1	m->1	n->8	u->1	
t tre	 ->4	:->1	d->21	v->1	
t tro	g->1	l->1	r->3	t->2	
t tru	p->1	s->1	
t try	c->2	
t trä	d->6	f->2	n->1	t->2	
t tuf	f->1	
t tun	g->3	
t tur	k->1	
t tus	e->1	
t tve	k->5	
t tvi	n->5	v->6	
t två	 ->9	:->1	n->1	
t tyc	k->7	
t tyd	l->30	
t tys	k->5	
t tyv	ä->2	
t täc	k->1	
t täm	l->2	
t tän	d->1	k->17	
t täp	p->2	
t tåg	,->1	e->1	
t tål	 ->1	
t ult	i->1	
t und	a->9	e->96	v->23	
t uni	k->1	o->11	
t upp	 ->21	,->3	.->2	b->1	d->12	e->9	f->19	g->6	h->8	k->3	l->4	m->17	n->37	r->23	s->7	t->6	v->3	
t ur 	U->1	b->1	d->1	e->2	m->1	p->1	s->1	
t ura	n->6	
t urh	o->1	
t urs	k->1	p->5	ä->1	
t urv	a->4	
t ut 	a->3	f->1	k->1	m->2	o->1	s->3	
t ut,	 ->9	
t ut.	 ->1	D->4	J->1	V->1	
t uta	n->19	r->18	
t utb	e->1	u->2	y->4	
t ute	s->8	
t utf	o->7	ä->3	ö->8	
t utg	i->1	j->1	å->2	ö->11	
t uth	ä->1	
t uti	f->3	
t utj	ä->3	
t utk	a->1	r->1	
t utl	a->1	ä->1	ö->1	
t utm	a->1	y->1	ä->15	
t utn	y->14	ä->3	
t uto	m->3	
t utp	e->1	l->1	r->1	
t utr	e->1	o->2	y->1	
t uts	a->3	e->2	k->20	l->2	t->2	ä->1	
t utt	a->24	j->1	r->28	ö->2	
t utv	a->1	e->27	i->20	ä->5	
t utö	k->8	v->5	
t vac	k->3	
t vad	 ->34	
t vag	t->1	
t vak	a->1	s->2	u->1	
t val	 ->4	,->1	.->1	d->7	u->2	
t van	a->1	l->4	
t var	 ->51	,->1	a->79	e->3	i->6	j->9	k->2	m->3	n->2	s->3	v->3	
t vat	t->4	
t ved	e->3	
t vem	 ->1	
t ver	k->48	
t vet	 ->7	a->4	e->6	t->1	
t vi 	1->1	a->17	b->34	d->11	e->7	f->23	g->16	h->46	i->66	j->3	k->41	l->3	m->30	n->7	o->14	p->5	r->9	s->42	t->8	u->10	v->12	ä->17	å->5	ö->2	
t vi,	 ->6	
t via	 ->3	
t vid	 ->47	,->2	.->2	a->2	h->1	m->1	t->25	
t vik	t->119	
t vil	a->1	j->13	k->12	l->84	
t vin	 ->1	n->3	s->2	
t vis	 ->6	.->1	a->28	e->4	s->31	t->1	
t vit	b->2	t->2	
t vol	u->1	
t vor	e->12	
t vra	k->1	
t väc	k->2	
t väg	 ->2	a->1	e->1	r->1	s->1	
t väl	 ->21	,->1	.->1	b->1	d->2	f->1	g->2	j->5	k->10	m->1	s->3	u->2	
t vän	d->6	l->1	s->1	t->7	
t vär	d->9	l->1	r->1	s->3	
t väs	e->7	
t väx	a->4	e->2	l->1	t->1	
t våg	a->1	
t vål	d->2	
t vår	 ->16	a->18	t->11	
t wor	s->1	
t ypp	e->1	
t ytt	e->15	r->19	
t zon	i->1	
t Öst	e->6	
t äck	l->1	
t äga	 ->17	
t äge	r->1	
t ägn	a->6	
t ämb	e->4	
t ämn	e->4	
t än 	a->5	b->1	d->3	e->4	f->1	i->3	m->2	p->1	s->2	v->1	ä->2	
t än,	 ->1	
t änd	a->5	r->55	å->1	
t änn	u->8	
t änt	l->2	
t är 	-->2	2->1	3->1	E->4	P->1	a->68	b->33	c->1	d->103	e->137	f->45	g->15	h->16	i->75	j->24	k->28	l->16	m->53	n->39	o->30	p->13	r->16	s->46	t->19	u->22	v->52	y->5	ä->7	ö->2	
t är,	 ->2	
t är.	.->1	
t är:	 ->1	
t ära	n->1	
t äre	n->5	
t ärl	i->1	
t äve	n->39	
t å e	n->3	
t åkl	a->1	
t åld	e->1	
t åli	g->4	
t ålä	g->2	
t år 	1->1	2->4	a->1	d->2	f->1	o->5	p->1	s->5	u->1	ä->1	
t år,	 ->4	
t år.	D->1	E->1	O->1	S->1	
t åre	t->1	
t årh	u->2	
t årl	i->1	
t års	b->1	
t åsi	k->1	
t åst	a->6	
t åt 	a->1	d->8	e->1	j->1	k->1	p->1	
t åta	 ->1	g->5	l->3	
t åte	r->50	
t åtf	ö->3	
t åtg	ä->10	
t åtm	i->3	
t åtn	j->1	
t åvi	l->1	
t öde	.->1	?->1	s->1	
t ögo	n->5	
t öka	 ->21	.->1	d->2	n->2	r->1	t->2	
t ökn	i->1	
t öl 	o->1	
t öms	e->1	
t öns	k->8	
t öpp	e->9	n->4	
t öst	e->15	
t öve	r->111	
t övr	i->2	
t! De	n->1	t->1	
t! Ja	g->2	
t! Nä	r->1	
t! So	m->1	
t! Va	d->1	
t!"Ja	g->1	
t!(Pa	r->1	
t!. (	F->1	
t!.(N	L->1	
t!Det	 ->1	
t!Där	f->1	
t!Her	r->3	
t!Jag	 ->1	
t!Kul	t->1	
t!Led	a->1	
t!Men	 ->1	
t!När	 ->1	
t!Pre	c->1	
t!Tvä	r->1	
t" (s	e->1	
t" gö	r->1	
t" me	d->1	
t" oc	h->1	
t" är	 ->1	
t", b	e->1	
t", d	e->1	
t", e	f->1	
t", s	o->1	
t".En	 ->1	
t".Ja	g->1	
t) (C	5->1	
t) C5	-->1	
t) ha	d->1	r->1	
t) på	 ->1	
t) so	m->1	
t) tä	c->1	
t), d	e->1	
t), s	o->1	
t), t	j->1	
t).De	t->1	
t).He	r->2	
t).Li	k->1	
t)Näs	t->1	
t, "e	n->1	
t, Co	s->1	
t, Da	g->1	
t, EG	-->1	
t, Ef	t->1	
t, Gi	l->1	
t, Ha	i->1	
t, II	 ->1	I->1	
t, In	g->1	
t, Jo	n->1	
t, La	 ->1	
t, Ob	e->1	
t, PV	C->1	
t, Sc	h->1	
t, So	a->1	
t, We	s->1	
t, Zi	m->1	
t, al	l->1	
t, an	n->1	s->2	v->1	
t, ar	r->1	t->1	
t, at	t->30	
t, av	 ->4	s->2	
t, be	d->1	g->3	t->1	v->2	
t, bl	.->3	i->1	
t, bo	r->1	
t, br	i->1	
t, by	r->1	
t, bö	r->6	
t, ci	v->1	
t, de	 ->4	c->1	l->4	m->4	n->9	t->20	
t, di	s->1	
t, dj	u->1	
t, dv	s->5	
t, dä	c->1	r->8	
t, då	 ->3	
t, ef	f->2	t->25	
t, el	l->6	
t, en	 ->14	e->1	l->4	
t, et	i->1	t->5	
t, ex	e->1	
t, fa	k->2	s->2	
t, fi	n->2	
t, fo	r->1	
t, fr	a->4	i->4	u->7	å->2	
t, fu	n->1	
t, få	r->3	
t, fö	r->39	
t, ge	n->4	
t, gi	v->1	
t, gl	ö->1	
t, gr	a->1	
t, gä	l->1	
t, gå	 ->1	r->3	t->1	
t, gö	r->2	
t, ha	 ->1	m->1	n->3	r->16	
t, he	l->1	r->20	
t, hj	ä->1	
t, ho	p->2	
t, hu	r->1	
t, hä	l->1	n->1	r->1	
t, hå	l->1	
t, i 	A->1	I->1	P->1	d->5	e->3	f->5	n->1	r->1	s->5	v->1	ö->2	
t, in	b->1	f->1	g->1	k->2	l->2	n->3	o->2	t->12	
t, ja	 ->1	g->3	
t, ju	s->3	
t, jä	m->2	
t, ka	l->3	n->8	
t, kl	a->1	
t, ko	m->12	n->3	
t, kr	a->1	i->1	ä->1	
t, ku	l->3	
t, kä	n->1	r->2	
t, la	d->1	
t, le	d->1	
t, li	k->4	t->1	
t, lä	g->1	m->1	
t, lå	n->1	t->1	
t, me	d->18	n->58	
t, mi	n->2	
t, mo	d->1	t->1	
t, my	c->3	
t, mä	n->1	
t, må	n->1	s->4	
t, na	r->1	t->3	
t, nä	m->8	r->8	
t, nå	g->1	
t, oa	n->1	v->1	
t, ob	e->1	
t, oc	h->109	k->1	
t, ol	i->1	
t, om	 ->19	d->1	e->1	f->1	v->1	
t, pa	r->1	
t, pe	r->1	
t, pl	a->1	
t, po	l->1	
t, pr	e->4	
t, på	 ->8	
t, ra	p->1	s->2	
t, re	g->1	s->1	
t, rä	d->1	t->2	
t, rå	d->2	
t, rö	r->1	
t, sa	m->3	
t, se	 ->1	d->2	t->1	x->1	
t, si	n->2	
t, sj	ä->1	
t, sk	a->6	r->1	u->2	
t, so	m->55	
t, sp	e->2	
t, st	a->1	r->1	å->1	
t, sä	k->28	r->7	
t, så	 ->22	v->3	
t, t.	e->1	
t, ta	c->3	
t, ti	l->6	
t, to	r->1	
t, tr	o->5	
t, tv	i->1	å->3	
t, ty	 ->3	v->1	
t, un	d->3	
t, up	p->2	
t, ur	 ->1	
t, ut	a->30	b->1	r->1	v->1	
t, va	d->4	l->1	r->8	
t, ve	k->1	m->1	
t, vi	 ->6	a->1	d->2	l->33	s->1	
t, vo	r->1	
t, vä	d->1	g->1	l->1	
t, vå	r->1	
t, än	d->2	
t, är	 ->17	a->1	
t, äv	e->13	
t, å 	a->1	
t, år	 ->1	
t, åt	e->2	
t, ök	a->1	
t, öp	p->1	
t- oc	h->3	
t-Exu	p->1	
t-ana	l->5	
t-ben	e->5	
t-frå	g->1	
t-sta	t->2	
t. (P	T->1	
t. 7 	l->1	
t. 7)	.->1	
t. Av	 ->1	
t. De	n->5	s->1	t->11	
t. Dä	r->1	
t. Et	t->1	
t. Fr	u->1	
t. He	r->1	
t. Hä	r->1	
t. I 	s->1	
t. In	g->1	t->1	
t. Ja	g->1	
t. Ko	s->1	
t. Me	n->1	
t. Of	f->1	
t. So	m->1	
t. Vi	 ->2	
t. Vå	r->1	
t. ai	d->1	
t.(Ar	b->1	
t.(FR	)->1	
t.(PT	)->1	
t.(Pa	r->1	
t.(Pr	o->1	
t.)An	d->1	
t.)Be	t->2	
t.)Fr	u->1	
t.)Re	f->1	
t.- H	e->1	
t.. (	E->2	
t..(D	A->1	
t...(	T->1	
t...F	r->1	
t..He	r->1	
t.199	8->1	
t.Acc	e->1	
t.Ald	r->1	
t.All	a->2	m->1	t->1	
t.Ans	v->1	
t.Anv	ä->1	
t.Ara	b->1	
t.Art	i->1	
t.Att	 ->2	
t.Av 	d->2	s->1	
t.Avs	l->6	
t.Ber	e->1	
t.Bet	r->1	ä->3	
t.Bil	l->1	
t.Bla	n->1	
t.Bor	d->1	
t.Bri	t->1	
t.Båd	a->2	
t.Dag	l->1	
t.De 	a->1	b->2	d->1	f->5	h->1	i->1	l->1	m->2	n->1	s->4	t->2	v->1	ä->1	å->1	
t.Del	s->1	v->1	
t.Den	 ->27	n->8	
t.Des	s->11	
t.Det	 ->141	s->1	t->28	
t.Dir	e->3	
t.Där	 ->1	f->15	v->1	
t.Då 	h->1	k->3	v->1	
t.EG-	d->1	
t.Eff	e->1	
t.Eft	e->6	
t.Eko	n->1	
t.En 	a->4	b->1	d->1	f->1	k->1	ö->1	
t.End	a->3	
t.Enl	i->6	
t.Erf	a->1	
t.Ett	 ->6	
t.Eur	o->10	
t.FPÖ	:->1	
t.Fel	a->1	
t.Fin	n->1	
t.Fle	r->1	
t.Flo	r->1	
t.Fra	m->5	n->1	
t.Fru	 ->10	
t.Frå	g->5	n->1	
t.Föl	j->2	
t.För	 ->25	d->3	e->4	s->4	u->1	v->2	
t.Gen	o->4	
t.Giv	e->1	
t.Gre	k->1	
t.Gru	p->1	
t.Han	 ->3	d->2	
t.Hel	a->1	
t.Her	r->48	
t.Hit	t->1	
t.Hur	 ->4	
t.Huv	u->1	
t.Här	 ->7	
t.I F	r->1	
t.I N	e->1	
t.I a	n->1	r->1	v->1	
t.I b	e->1	
t.I d	a->3	e->10	
t.I e	g->1	n->1	
t.I f	o->1	r->2	ö->1	
t.I k	o->1	
t.I l	i->1	
t.I m	o->2	
t.I n	ä->1	
t.I o	c->1	
t.I r	e->2	
t.I s	a->2	t->1	å->1	
t.I u	t->1	
t.I v	i->1	ä->1	å->3	
t.I ä	n->1	
t.Ibl	a->1	
t.Ing	e->1	
t.Inn	e->1	
t.Ins	a->1	
t.Int	e->2	
t.Ja 	t->1	
t.Ja,	 ->2	
t.Jag	 ->144	
t.Ju 	m->1	
t.Jus	t->1	
t.Kom	m->14	
t.Kon	k->3	s->1	
t.Kra	v->1	
t.Kul	t->2	
t.Kär	a->2	
t.La 	R->1	
t.Lik	s->1	
t.Lit	t->1	
t.Län	d->1	
t.Lån	 ->1	
t.Låt	 ->10	
t.Man	 ->14	
t.Mar	k->1	
t.Max	i->1	
t.Med	 ->7	a->1	b->1	g->1	l->1	
t.Mel	l->1	
t.Men	 ->39	
t.Mer	 ->1	
t.Mil	j->1	
t.Min	 ->7	a->4	s->1	
t.Mor	a->1	
t.Mot	 ->3	
t.Mån	g->1	
t.Nat	i->1	u->4	
t.Ni 	b->1	f->1	h->2	t->1	v->2	
t.Nu 	h->3	k->1	m->1	t->1	
t.Num	e->1	
t.Nuv	a->1	
t.När	 ->10	
t.Näs	t->1	
t.Någ	o->1	
t.Nöd	v->1	
t.OK,	 ->1	
t.Obe	r->1	
t.Och	 ->12	
t.Off	e->1	
t.Om 	d->3	j->1	k->1	m->2	n->2	s->1	u->1	v->5	
t.Ord	f->1	
t.Ork	a->1	
t.Oro	n->1	
t.PPE	-->1	
t.Par	l->8	
t.Plä	d->1	
t.Por	t->1	
t.Pre	c->1	
t.Pro	b->1	d->1	j->1	
t.Pun	k->1	
t.På 	d->3	g->1	m->1	s->2	
t.Rap	p->1	
t.Red	a->1	
t.Reg	e->1	
t.Res	u->1	
t.Rik	t->1	
t.Rät	t->1	
t.Sam	t->2	
t.San	n->1	
t.Sed	a->1	
t.Ska	l->1	
t.Sko	t->1	
t.Sku	l->1	
t.Slu	t->6	
t.Soc	i->1	
t.Som	 ->5	
t.Sta	b->1	t->3	
t.Sto	r->1	
t.Stö	d->2	r->1	
t.Syf	t->1	
t.Så 	d->1	h->1	j->2	k->1	l->2	s->1	v->1	
t.Såv	ä->1	
t.Tac	k->6	
t.Tan	k->1	
t.The	a->1	
t.Til	l->4	
t.Tre	 ->1	
t.Tro	t->2	
t.Tus	e->1	
t.Två	 ->1	
t.Ty 	i->1	u->1	
t.Tyv	ä->1	
t.Und	e->3	
t.Ung	e->1	
t.Uni	o->1	
t.Ur 	p->1	
t.Utb	i->1	
t.Utf	ö->1	
t.Uts	k->1	
t.Vad	 ->15	
t.Val	e->1	
t.Var	f->5	j->2	
t.Vi 	a->2	b->5	d->1	e->1	f->9	g->2	h->17	i->1	k->11	m->9	r->3	s->4	t->1	u->2	v->11	ä->5	
t.Vid	 ->2	a->1	
t.Vil	l->1	
t.Vis	s->2	
t.Väs	t->1	
t.Vår	 ->2	a->1	
t.ex.	 ->20	
t.o.m	.->7	
t.Änd	a->1	r->2	
t.Är 	d->1	
t.Äve	n->7	
t.Å a	n->2	
t.Å e	n->1	
t.År 	2->1	
t.Åre	t->1	
t.Åte	r->1	
t.Öka	d->1	
t.Öst	e->1	
t.Övr	i->1	
t: "D	e->2	
t: "M	i->1	
t: "a	l->1	
t: Ef	t->1	
t: Fr	i->1	
t: Ho	l->1	
t: Ja	g->2	
t: Un	i->1	
t: Ut	v->1	
t: Vi	 ->1	
t: at	t->1	
t: de	n->2	t->3	
t: en	 ->1	
t: et	t->1	
t: fr	å->1	
t: fö	r->1	
t: ha	n->1	
t: ja	g->2	
t: ka	n->1	
t: mi	n->1	
t: om	 ->2	
t: sy	s->1	
t: ta	n->1	
t: ut	b->1	
t: vi	 ->1	
t: vå	r->1	
t: ön	s->1	
t; Da	n->1	
t; al	l->1	
t; ar	t->1	
t; de	 ->1	t->4	
t; en	d->1	
t; fo	r->1	
t; fr	i->1	
t; un	d->1	
t; å 	e->1	
t? Me	d->1	
t? Rå	d->1	
t?. (	E->2	
t?.(E	N->2	
t?Ans	l->1	
t?Att	 ->1	
t?Av 	t->1	
t?De 	t->1	
t?Det	 ->3	
t?Ett	 ->1	
t?Eur	o->1	
t?Her	r->1	
t?Hur	 ->2	
t?I v	i->1	
t?Jag	 ->4	
t?Jo 	d->1	
t?Kom	m->1	
t?Kär	a->1	
t?Nej	,->2	.->1	
t?Ni 	k->1	n->1	
t?När	 ->1	
t?Och	 ->1	
t?Om 	i->1	
t?RIN	A->1	
t?Sku	l->2	
t?Tän	k->1	
t?Utg	i->1	
t?Vad	 ->1	
t?Vi 	b->1	
t?Vil	k->2	
t?Vis	s->1	
t?Är 	d->1	
tBetä	n->1	
tJag 	h->1	
tNäst	a->1	
ta - 	a->1	f->1	j->1	m->1	o->1	r->1	ä->1	
ta -,	 ->1	
ta 10	 ->1	
ta Al	t->1	
ta Am	s->1	
ta EG	-->5	
ta EU	:->1	
ta Eu	r->4	
ta FP	Ö->1	
ta Jö	r->1	
ta Ma	r->1	
ta Na	t->1	
ta Sh	e->1	
ta St	a->1	
ta ab	s->1	
ta ad	j->1	
ta ak	t->1	
ta al	l->6	t->1	
ta an	 ->1	b->1	d->1	g->1	n->1	s->10	t->1	v->5	
ta ar	b->8	g->1	
ta at	t->47	
ta av	 ->23	.->1	s->6	
ta ba	r->2	
ta be	d->1	f->1	g->5	h->9	k->1	l->1	s->12	t->64	v->1	
ta bi	b->3	d->2	l->4	n->1	s->1	
ta bl	i->7	
ta bo	r->4	
ta br	o->2	
ta bu	d->3	
ta bä	r->1	
ta bö	r->6	
ta ce	r->2	
ta ch	a->1	
ta da	g->3	t->1	
ta de	 ->22	b->3	c->2	f->1	l->24	m->9	n->22	r->2	s->8	t->27	
ta di	g->1	l->1	p->1	r->34	s->2	
ta dj	u->1	
ta do	k->6	
ta dr	i->1	o->1	
ta dä	r->1	
ta dö	r->1	
ta ef	f->3	t->3	
ta eg	e->1	
ta ek	o->2	
ta el	l->3	v->1	
ta em	o->9	
ta en	 ->46	b->1	d->1	h->2	o->1	v->1	
ta er	 ->5	b->3	f->3	
ta et	t->36	
ta ev	e->1	
ta ex	p->1	
ta fa	k->3	l->18	s->1	
ta fe	m->1	
ta fi	n->1	s->1	
ta fl	e->2	
ta fo	l->1	r->25	
ta fr	a->14	i->3	å->20	
ta fu	l->2	n->1	
ta få	 ->1	g->2	r->4	
ta fö	l->2	r->140	
ta ga	r->2	
ta ge	m->6	n->6	
ta gi	g->1	l->1	
ta gl	ö->1	
ta go	d->3	
ta gr	a->2	o->1	u->7	ä->1	
ta gä	l->9	
ta gå	n->21	
ta gö	r->2	
ta ha	l->1	n->36	r->30	
ta he	l->4	
ta hi	n->3	
ta hj	ä->1	
ta ho	m->1	n->1	s->1	t->1	
ta hu	r->2	s->1	
ta hä	n->31	v->1	
ta hå	l->2	
ta i 	D->2	E->1	a->2	b->1	d->11	e->7	f->3	g->2	l->2	m->3	n->2	o->3	p->1	r->1	s->3	t->1	u->2	v->4	y->2	ö->1	
ta id	é->1	
ta ig	e->3	
ta ih	j->1	
ta in	 ->3	d->1	f->1	i->8	l->3	n->12	o->2	s->3	t->20	v->2	
ta is	ä->1	
ta it	u->14	
ta jo	r->1	
ta ju	s->1	
ta ka	n->17	r->1	
ta kl	a->3	i->1	
ta ko	d->1	l->5	m->18	n->10	
ta kr	a->3	i->3	ä->4	
ta ku	n->1	
ta kv	a->2	i->1	
ta kä	l->1	n->1	r->3	
ta la	g->3	n->5	
ta le	d->1	g->1	
ta li	g->5	t->1	v->3	
ta lj	u->1	
ta lä	g->2	m->1	n->1	r->3	t->1	
ta lå	n->1	
ta ma	n->6	r->1	t->1	
ta me	d->70	n->3	r->3	t->2	
ta mi	g->6	l->2	n->1	s->1	t->4	
ta mo	b->1	d->1	n->1	t->8	
ta my	c->8	g->1	n->1	
ta mä	n->1	r->1	
ta må	l->5	n->4	s->19	
ta mö	j->17	t->4	
ta na	m->1	t->13	
ta no	g->2	r->2	
ta nu	 ->1	l->1	
ta ny	a->4	c->1	
ta nä	m->2	r->7	t->1	
ta nå	g->4	
ta oa	v->1	
ta ob	e->1	
ta oc	h->33	k->6	
ta oe	n->1	
ta of	f->1	
ta og	e->1	
ta ol	i->1	j->1	y->2	
ta om	 ->30	,->1	.->1	f->4	g->1	r->35	s->1	v->1	
ta on	d->1	
ta or	d->8	g->2	i->1	s->1	ä->1	
ta os	s->13	
ta pa	k->1	l->1	r->40	
ta pl	a->2	e->1	
ta po	l->5	s->1	
ta pr	a->3	e->4	i->3	o->38	
ta pu	n->38	
ta på	 ->43	,->1	.->1	m->1	p->2	s->1	
ta ra	m->2	n->12	p->3	
ta re	d->2	f->2	g->16	n->1	s->14	
ta ri	g->1	k->2	s->3	
ta ru	b->1	n->1	
ta rä	t->1	
ta rå	d->3	
ta rö	r->4	
ta sa	d->2	k->3	m->40	n->2	
ta se	 ->1	i->1	k->6	n->1	t->1	
ta si	d->2	f->1	g->29	n->5	t->7	
ta sj	u->1	ä->1	
ta sk	a->13	e->5	i->4	u->10	y->3	ä->2	
ta sl	a->10	u->3	
ta sm	u->1	å->2	
ta sn	a->1	
ta so	m->23	
ta sp	e->6	
ta st	a->20	e->5	o->6	r->6	y->1	ä->10	å->5	ö->6	
ta sv	a->1	å->1	
ta sy	f->2	n->5	s->4	
ta sä	g->3	k->1	s->1	t->20	
ta så	 ->3	n->1	
ta ta	g->1	l->5	n->2	r->1	s->2	
ta te	c->2	k->2	m->1	r->1	
ta ti	d->3	l->29	
ta tj	ä->1	
ta to	g->2	l->1	n->1	r->1	t->1	
ta tr	e->1	o->1	
ta tu	s->1	
ta tv	i->2	å->2	
ta ty	c->2	d->2	
ta tå	l->1	
ta un	d->4	i->3	
ta up	p->76	
ta ur	 ->3	a->1	
ta ut	 ->1	a->5	b->1	e->1	g->2	h->1	k->2	m->2	r->1	s->2	t->3	v->7	ö->1	
ta va	d->8	p->2	r->13	
ta ve	c->1	d->1	m->1	r->3	
ta vi	 ->5	d->2	k->5	l->15	s->5	
ta vo	r->1	
ta vä	g->1	k->1	s->2	
ta vå	l->1	r->4	
ta yt	t->2	
ta Ös	t->2	
ta äg	a->6	
ta äm	b->1	n->2	
ta än	d->11	t->1	
ta är	 ->163	,->3	.->1	e->2	
ta äv	e->4	
ta år	,->2	.->1	e->1	h->1	
ta ås	i->1	
ta åt	a->3	e->1	g->14	
ta ök	a->3	n->1	
ta öv	e->12	
ta!De	t->1	
ta!Fr	u->1	
ta, a	l->1	t->3	v->1	
ta, b	l->1	
ta, d	e->2	v->1	
ta, e	f->1	l->1	n->2	
ta, f	r->2	ö->7	
ta, h	a->2	e->2	u->2	
ta, i	 ->3	n->1	
ta, j	a->1	
ta, k	a->2	
ta, l	i->1	
ta, m	e->8	å->1	
ta, o	c->14	m->4	
ta, r	e->1	i->1	
ta, s	a->1	o->3	å->2	
ta, t	e->1	i->2	
ta, u	t->6	
ta, v	a->1	i->1	
ta. D	e->1	
ta. F	ö->1	
ta. V	a->1	
ta.(P	a->1	
ta.)F	r->1	
ta.- 	(->1	
ta.. 	H->1	
ta..(	N->1	
ta.An	n->1	
ta.Be	r->1	t->1	
ta.Co	r->1	
ta.De	 ->1	n->6	t->19	
ta.Dä	r->1	
ta.Då	 ->1	
ta.Ef	t->3	
ta.Em	e->1	
ta.En	 ->1	l->1	
ta.Fr	å->1	
ta.Fö	r->2	
ta.Ge	r->1	
ta.He	r->4	
ta.I 	d->1	f->1	l->1	r->1	s->1	
ta.In	o->1	t->1	
ta.Ja	g->12	
ta.Ko	m->1	
ta.Me	d->2	n->5	
ta.Nu	 ->1	
ta.Nä	r->1	
ta.Oc	h->2	
ta.Om	 ->2	
ta.Pr	e->1	o->1	
ta.På	 ->1	
ta.Se	d->1	
ta.Si	t->1	
ta.Sj	u->1	
ta.So	m->1	
ta.St	a->1	ö->1	
ta.Så	 ->1	
ta.To	p->1	
ta.Tr	o->1	
ta.Va	d->3	r->1	
ta.Vi	 ->11	
ta.Vå	r->1	
ta.Är	 ->1	
ta: I	 ->1	
ta: J	a->2	
ta: V	e->1	
ta: u	p->1	
ta: v	i->1	
ta; d	e->1	
ta; v	i->1	
ta?De	t->1	
ta?Ja	g->1	
ta?Nä	r->1	
ta?Vi	s->1	
taNäs	t->1	
taaff	ä->1	
tab s	k->1	
tabas	e->1	
tabeh	a->1	
tabel	 ->3	!->1	,->3	.->3	l->6	t->21	
tabil	 ->2	a->2	i->18	t->2	
tabla	 ->9	,->1	.->3	
table	r->13	
tabri	e->3	
tabu 	i->1	
tabul	a->1	
tack 	f->2	g->2	m->1	o->3	p->1	s->2	t->11	v->7	
tack,	 ->1	
tack.	H->1	J->1	
tacka	 ->84	r->21	
tacke	n->1	
tackl	a->1	
tacko	r->1	
tacks	a->9	
tad a	t->1	
tad f	e->1	ö->5	
tad m	e->2	o->1	
tad o	c->2	m->1	
tad p	å->2	
tad s	i->1	
tad ö	v->1	
tad, 	a->1	e->1	
tad."	M->1	
tad.(	S->1	
tad.D	e->1	
tad.F	r->1	
tad.H	e->3	
tad.J	a->1	
tad.M	e->1	ä->1	
tad.O	m->14	
tad.R	e->1	
tade 	"->1	E->1	O->1	a->8	b->3	d->3	e->8	f->5	g->1	i->4	j->1	k->1	m->6	o->3	p->6	r->1	s->4	t->2	u->2	v->2	å->1	
tade,	 ->3	
tade.	 ->1	E->1	T->1	
tadel	s->2	
tades	 ->13	,->1	
tadga	 ->14	,->1	d->1	n->10	r->2	
tadgo	r->1	
tadie	t->4	
tadiu	m->4	
tadko	m->24	
tadmi	n->2	
tadsb	e->1	
tadsc	e->1	
tadso	m->1	
tadsp	r->1	
tadt,	 ->1	
tafrå	g->10	
tag a	t->1	v->2	
tag b	e->1	
tag e	f->1	n->1	
tag f	r->2	ö->3	
tag g	ä->1	
tag h	a->4	e->1	
tag i	 ->5	,->1	n->5	
tag k	a->2	o->2	
tag l	e->1	i->1	
tag n	ä->1	
tag o	c->6	m->1	
tag p	å->3	
tag s	a->1	e->2	k->1	o->16	t->1	
tag t	i->1	
tag u	t->1	
tag v	i->2	
tag ä	r->3	
tag, 	e->3	f->2	m->3	n->1	o->3	s->4	t->1	u->2	v->1	
tag.A	v->1	
tag.D	e->3	ä->1	
tag.E	f->2	
tag.F	ö->1	
tag.I	 ->2	n->1	
tag.J	u->1	
tag.K	o->2	
tag.M	å->1	
tag.O	c->1	
tag.R	a->1	
tag.S	k->1	
tag.T	i->1	
tag.V	a->1	i->1	
tag?F	ö->1	
tagan	d->102	
tagar	a->2	e->48	l->3	n->16	v->1	
tagba	r->15	
tagel	s->1	
tagen	 ->34	,->6	.->5	:->1	;->1	s->21	
taget	 ->18	.->3	s->1	
tagit	 ->75	,->2	.->1	s->22	
tagli	g->5	
tagna	 ->8	,->1	t->1	
tagne	 ->7	r->1	s->1	
tagni	n->3	s->1	
tags 	f->1	p->1	v->1	
tagsa	m->3	v->1	
tagsb	e->1	
tagse	k->5	
tagsf	a->1	ö->2	
tagsg	r->2	
tagsi	n->1	
tagsj	u->2	
tagsk	o->1	
tagsl	i->1	
tagsm	ä->1	
tagsn	e->1	
tagsr	e->3	å->2	
tagss	t->3	
tagst	i->2	
tain,	 ->1	
taine	 ->1	
tains	a->2	t->22	
tak f	ö->1	
tak, 	a->1	v->1	
taka 	b->2	p->1	r->1	t->1	
takel	 ->2	
taket	 ->1	
takla	s->1	
takt 	m->6	o->1	ä->1	
takt.	M->2	
takte	r->12	
takti	k->2	s->2	
takul	ä->1	
tal -	 ->1	
tal a	v->4	
tal b	e->2	i->2	r->1	
tal d	e->1	
tal e	f->1	
tal f	o->1	r->4	å->1	ö->3	
tal h	a->1	ä->1	
tal i	 ->5	n->8	
tal k	o->2	v->2	
tal l	ä->2	
tal m	a->1	e->15	i->1	o->1	ä->1	å->2	
tal n	y->1	
tal o	c->6	m->7	
tal p	e->1	o->1	r->1	å->1	
tal r	e->3	i->1	o->1	
tal s	a->2	k->2	o->16	v->1	ä->1	
tal t	i->3	y->1	
tal u	p->1	t->1	
tal v	e->1	
tal ä	r->3	
tal å	s->1	
tal ö	v->3	
tal" 	m->1	
tal, 	g->1	h->1	o->2	s->1	v->1	
tal-F	i->3	
tal.D	e->1	
tal.E	n->1	
tal.F	ö->1	
tal.H	e->2	
tal.I	 ->1	
tal.J	a->1	
tal.K	a->1	o->1	
tal.S	a->1	
tal.V	i->1	
tal: 	O->1	
talFi	n->1	
tala 	K->1	a->3	b->2	d->2	e->5	f->4	h->1	i->2	k->1	m->14	n->1	o->41	r->1	s->18	t->3	u->3	v->3	ä->1	å->3	
tala"	;->1	
tala,	 ->3	
tala.	D->4	I->1	J->1	
tala?	D->3	
talad	 ->1	e->34	
talan	 ->1	.->1	d->52	g->1	s->2	
talar	 ->67	,->2	.->2	?->1	e->30	n->13	s->1	t->2	
talas	 ->10	,->1	
talat	 ->20	,->3	.->2	e->1	s->6	
talbe	l->1	
talbl	o->1	
talen	 ->11	,->1	.->3	
tales	m->2	ä->2	
talet	 ->44	,->9	.->5	s->3	
talfå	n->4	
talfö	r->1	
talie	n->36	
talig	 ->1	t->1	
talin	i->2	
talis	m->1	t->1	
talit	a->2	e->1	
talj 	o->1	ö->1	
talj,	 ->2	
talj.	V->1	
talja	n->1	
talje	r->26	
taljf	l->1	
taljk	o->2	
tall,	 ->1	
talld	e->1	
talle	r->9	
talli	n->1	
tallk	l->2	
talma	n->418	
talni	n->15	
talog	 ->2	
talri	k->4	
tals 	a->2	b->1	f->2	g->1	h->1	i->1	k->1	m->5	o->2	p->1	s->1	å->2	
tals.	D->1	
talsf	a->1	
talsk	a->3	u->1	
talsl	ö->1	
talsp	a->1	u->6	
talsr	u->1	
talss	t->1	
talsu	m->1	
talt 	2->1	9->1	a->1	f->1	s->1	t->1	
talt.	V->1	
talte	r->1	
talts	 ->1	
talvo	l->1	
talys	a->2	
tame-	f->1	
tamen	t->8	
tamin	a->1	e->1	
tamp 	i->1	
tan 1	0->2	7->1	
tan I	s->1	
tan a	l->1	n->2	r->1	t->61	v->2	
tan b	a->3	e->2	i->1	o->1	
tan d	a->1	e->29	r->2	ö->1	
tan e	f->1	l->1	n->11	r->1	t->3	
tan f	i->1	r->1	y->2	ö->7	
tan g	o->1	å->2	
tan h	a->2	e->2	i->1	ä->4	
tan i	 ->3	d->2	n->5	
tan j	a->1	
tan k	a->2	l->1	o->6	r->2	v->1	
tan m	a->2	e->3	i->2	o->1	å->1	ö->1	
tan n	o->1	u->1	å->8	
tan o	c->40	m->6	r->2	
tan p	a->1	r->1	u->1	å->15	
tan r	e->2	i->2	ä->1	
tan s	a->1	k->1	n->8	o->4	t->2	å->1	
tan t	e->1	i->2	v->34	
tan u	n->1	p->2	t->1	
tan v	a->1	e->1	i->4	ä->1	
tan ä	r->26	v->10	
tan ö	p->2	v->4	
tan, 	K->1	U->1	e->3	g->1	i->1	n->1	s->2	
tan.(	P->2	
tan.A	v->1	
tan.D	e->1	
tan.F	ö->1	
tan.H	e->1	
tan.J	a->4	
tan.M	e->1	
tan.S	å->1	
tan.T	a->1	
tan.U	t->1	
tan.V	i->3	
tan; 	d->1	
tan?Ä	r->1	
tana 	d->1	
tanbu	l->1	
tanda	 ->1	r->24	
tande	 ->102	,->5	.->4	f->6	h->1	l->2	n->2	r->2	t->34	
tanen	 ->2	.->1	
taner	 ->1	n->4	
tanfö	r->32	
tank-	 ->1	
tanka	r->16	
tanke	 ->48	,->2	b->1	f->1	g->1	n->11	p->1	r->4	
tankf	a->7	o->1	
tankr	a->5	e->2	
tanna	 ->5	r->2	t->3	
tanni	e->14	
tano 	o->1	
tans 	a->2	d->3	f->1	i->1	m->1	o->2	p->1	s->2	
tans,	 ->6	
tans.	M->1	
tans?	.->1	
tanse	n->3	r->5	
tansk	a->6	
tansl	a->1	
tansr	ä->22	
tansv	a->6	ä->7	
tant 	f->1	o->1	
tant,	 ->1	
tante	n->3	r->9	
tanti	e->2	s->1	
tanvä	n->1	
tapol	i->1	
tapp 	d->1	
tappa	 ->1	r->2	
tappe	n->1	r->3	
tar A	l->1	
tar E	u->1	
tar F	l->1	
tar a	k->1	l->3	n->2	t->13	v->2	
tar b	a->1	e->9	i->2	
tar d	e->27	ä->1	
tar e	f->3	m->3	n->9	t->3	x->2	
tar f	l->1	r->2	u->1	ö->14	
tar g	e->2	ä->1	å->1	ö->1	
tar h	a->2	e->1	i->1	ä->1	
tar i	 ->12	g->1	n->10	t->6	
tar j	a->9	u->2	
tar k	a->1	o->3	u->2	
tar l	ä->1	
tar m	a->2	e->10	i->14	o->2	
tar n	i->3	o->1	y->2	å->1	
tar o	a->1	c->10	f->1	l->1	m->9	s->2	
tar p	a->1	å->23	
tar r	i->1	ö->1	
tar s	i->16	k->1	l->2	o->6	t->3	ä->2	
tar t	i->30	r->1	v->2	
tar u	n->2	p->11	t->6	
tar v	a->1	e->3	i->12	ä->1	
tar y	t->1	
tar ä	n->1	r->1	
tar ö	v->3	
tar, 	P->1	f->1	n->1	o->2	u->1	
tar.D	e->3	
tar.F	ö->1	
tar.J	a->1	
tar.M	e->1	
tar.V	i->2	
tar.Ä	n->1	
tarbe	t->32	
tare 	a->9	b->2	f->2	h->1	i->1	k->4	o->3	p->1	r->1	s->3	t->2	u->1	ä->1	
tare,	 ->6	
tare.	F->1	K->1	P->1	
taren	 ->4	,->2	.->2	
tarer	 ->15	,->3	.->2	n->1	
tarhu	s->1	
taria	t->2	
tarik	e->9	
tarin	n->1	
taris	e->2	k->13	m->6	t->2	
tarit	e->3	
tariu	m->1	
tark 	e->1	f->2	k->2	o->1	p->3	s->1	v->1	
tark,	 ->1	
tarka	 ->13	,->1	r->6	s->5	
tarke	 ->1	
tarkl	a->1	
tarkt	 ->21	,->1	.->1	
tarlø	n->2	
tarma	d->4	t->6	
tarna	 ->9	,->1	.->4	?->1	s->4	
tarta	 ->4	d->1	r->2	s->2	t->2	
tarte	n->3	r->1	
tartp	l->1	
tarvl	i->1	
tas a	n->1	t->4	v->19	
tas b	e->1	l->1	o->3	
tas c	e->1	
tas d	e->6	ä->2	
tas e	l->1	n->5	t->2	x->1	
tas f	a->1	r->3	ö->5	
tas g	e->3	
tas h	ä->1	
tas i	 ->20	n->8	
tas j	u->1	
tas k	o->2	
tas l	e->3	
tas m	e->6	o->3	y->3	å->1	
tas n	a->1	e->1	i->1	u->1	ä->1	å->1	
tas o	c->3	m->4	
tas p	r->1	å->8	
tas r	ö->1	
tas s	e->1	k->1	o->8	ä->1	ö->1	
tas t	i->2	
tas u	n->4	p->12	r->1	t->3	
tas v	a->3	i->5	ä->1	
tas ä	n->1	r->1	v->1	
tas, 	e->1	f->2	i->1	l->1	m->1	o->1	s->1	v->1	ä->1	
tas. 	P->1	
tas.B	e->1	
tas.D	ä->1	
tas.F	ö->1	
tas.J	a->1	o->1	ä->1	
tas.O	m->1	
tas.P	a->1	e->1	å->1	
tas.V	a->1	i->2	
tas.Ä	n->1	
tasie	n->1	
tasif	u->1	
tasin	 ->1	
task 	f->1	
taspe	k->2	
tast 	m->1	
taste	 ->1	
tasti	s->9	
tastr	o->90	
tasäk	e->1	
tat -	 ->2	
tat a	l->1	t->6	v->9	
tat b	e->3	o->1	
tat d	e->7	ä->2	
tat e	m->3	n->2	r->1	t->5	
tat f	r->4	å->2	ö->13	
tat g	r->1	ö->1	
tat h	a->8	e->1	
tat i	 ->8	g->2	n->2	
tat k	o->2	
tat l	ä->3	
tat m	a->1	e->4	o->4	y->1	å->2	
tat n	ä->1	
tat o	c->9	m->6	s->3	
tat p	a->1	r->1	å->4	
tat r	å->1	
tat s	i->7	k->1	o->12	t->3	ä->1	å->3	
tat t	a->1	i->2	
tat u	n->4	p->1	t->1	
tat v	a->4	i->2	
tat ä	n->1	r->1	
tat å	t->1	
tat, 	d->1	e->2	i->1	k->2	l->1	m->1	o->4	p->1	s->1	u->1	v->1	
tat. 	F->1	O->1	
tat.B	e->1	
tat.D	e->7	ä->1	
tat.E	n->2	
tat.G	r->1	
tat.H	e->2	
tat.I	 ->3	
tat.J	a->4	
tat.K	o->2	
tat.L	ä->1	
tat.O	c->1	m->1	
tat.P	r->1	
tat.T	r->1	
tat: 	h->1	j->1	
tat?.	(->1	
tat?J	o->1	
tate 	c->2	
taten	 ->25	,->6	.->6	s->5	
tater	 ->60	,->10	-->1	.->16	;->1	?->1	a->40	n->209	s->3	
tatet	 ->26	.->3	
tatin	r->1	
tatio	n->33	
tatis	t->9	
tativ	 ->4	a->6	i->1	t->4	
tatli	g->100	s->1	
tator	l->1	
tats 	-->1	a->6	d->1	e->1	f->1	i->4	k->1	l->1	m->5	n->2	o->1	p->1	r->3	s->3	t->2	u->4	v->1	
tats,	 ->2	
tats-	 ->5	
tats.	D->2	K->1	
tatsb	a->2	
tatsk	a->1	
tatsm	a->2	i->2	
tatsn	i->4	
tatsp	r->1	
tatss	t->19	
tatta	c->1	v->7	
tatue	r->2	
tatur	e->2	k->1	
tatus	 ->4	.->1	?->1	e->1	f->1	
tatöv	e->6	
tatür	k->1	
tauen	,->1	
tauni	o->3	
taure	r->1	
tav o	c->1	
tav ö	k->1	
tavla	 ->4	"->2	n->1	
tavli	g->1	
tax-f	r->3	
taxer	i->1	
tbala	n->2	
tbank	e->4	
tbarh	e->1	
tbart	 ->2	
tbasi	s->1	
tbasu	n->1	
tbefo	g->2	
tbeho	v->1	
tbest	ä->4	
tbeta	l->7	
tbeva	k->1	
tbild	a->7	e->1	n->57	
tbloc	k->1	
tbok 	h->1	m->1	o->5	s->3	ä->2	
tbok,	 ->1	
tbok.	D->1	H->1	J->1	T->1	V->1	
tboke	n->35	
tboll	s->1	
tbran	s->1	
tbred	n->4	
tbrin	g->1	
tbud 	o->3	
tbuds	i->1	
tbure	t->1	
tbygg	n->2	t->1	
tbyta	 ->1	
tbyte	 ->10	,->1	t->5	
tc. o	c->1	
tc. Ä	m->1	v->1	
tc.De	t->1	
tc.En	 ->1	
tc?At	t->1	
tchan	d->1	
tcher	 ->1	
tdela	r->1	
tdeln	i->2	
tdemo	k->11	
tdera	 ->1	
tdikt	e->1	
tdire	k->1	
te (K	u->2	
te - 	a->1	d->1	i->1	k->1	m->1	n->1	p->1	ä->1	
te -,	 ->1	
te 19	9->1	
te Be	r->1	
te EM	U->1	
te EU	 ->1	:->1	
te Ek	o->1	
te Eu	r->8	
te FN	:->1	
te Fo	U->1	
te Is	r->1	
te Jo	n->1	
te Ou	v->1	
te Qu	e->1	
te ab	s->1	
te ac	c->11	
te ag	e->1	
te ak	t->1	
te al	l->42	
te an	 ->1	a->3	d->1	i->1	n->1	p->3	s->8	t->4	v->7	
te ar	b->4	g->1	
te as	p->1	t->1	
te at	t->76	
te au	t->4	
te av	 ->16	g->1	s->5	t->1	v->2	
te ba	r->91	
te be	a->2	d->5	f->4	g->5	h->11	i->1	k->3	r->2	s->8	t->11	v->3	
te bi	d->1	o->1	
te bl	a->1	e->1	i->25	u->2	
te bo	r->2	v->1	
te br	e->1	i->1	
te by	g->1	
te bä	r->2	
te bö	r->10	
te ce	n->1	
te ch	e->2	
te co	n->2	
te da	g->5	
te de	 ->12	b->1	c->2	f->1	g->1	l->6	m->2	n->21	s->6	t->41	
te di	r->2	s->1	
te do	c->5	
te dr	a->2	ö->1	
te dä	r->14	
te då	 ->3	
te dö	l->1	m->1	
te ef	t->2	
te ek	o->1	
te el	l->3	
te em	e->1	
te en	 ->15	b->9	d->10	g->1	i->1	s->8	
te ep	o->1	
te er	.->1	b->1	f->1	i->1	k->3	s->1	
te et	t->12	
te eu	r->2	
te ev	e->1	
te ex	 ->1	e->2	i->2	
te fa	k->1	l->5	n->3	s->7	t->2	
te fe	m->2	
te fi	c->1	n->23	
te fo	r->10	
te fr	a->3	e->1	i->1	ä->2	å->7	
te fu	l->1	n->6	
te fy	r->1	
te fä	s->1	
te få	 ->14	r->14	t->2	
te fö	l->2	r->84	
te ga	r->5	v->1	
te ge	 ->9	m->3	n->13	r->3	t->2	
te gi	v->1	
te gj	o->3	
te gl	ö->10	
te go	d->9	
te gr	a->3	u->1	
te gä	l->4	
te gå	 ->9	n->1	r->7	t->2	
te gö	m->1	r->29	
te ha	 ->11	d->9	f->1	l->2	n->12	r->75	
te he	l->48	m->1	r->1	
te hi	n->2	t->1	
te hj	ä->2	
te ho	n->2	p->1	t->1	
te hu	r->3	
te hä	n->3	r->3	
te hå	l->5	
te hö	g->1	l->1	r->4	
te i 	B->1	D->1	H->1	K->1	L->1	a->3	d->4	e->4	f->5	g->2	k->1	m->1	n->4	r->1	s->10	t->6	å->1	
te ia	k->2	
te if	r->3	
te ig	n->1	
te il	l->1	
te in	b->2	d->1	f->10	g->3	l->2	n->4	o->5	r->2	s->8	t->8	v->1	
te is	o->1	
te ja	g->9	
te jo	r->1	
te ju	 ->2	s->1	
te jä	m->1	
te ka	m->1	n->58	
te kl	a->3	
te kn	ä->1	
te ko	m->38	n->10	r->1	
te kr	a->3	i->2	o->1	ä->3	
te ku	n->18	
te kv	a->1	i->1	
te kä	n->4	
te kö	r->1	
te la	d->1	g->2	
te le	d->9	t->1	
te li	g->4	
te lu	r->1	
te ly	c->7	
te lä	g->2	m->3	n->30	r->1	t->3	
te lå	n->1	s->1	t->6	
te lö	n->1	p->1	s->5	
te ma	k->1	n->23	
te me	d->50	l->8	n->1	r->3	t->1	
te mi	g->1	n->18	s->3	
te mo	b->1	d->1	t->4	
te my	c->5	
te må	l->2	n->11	s->2	
te mö	j->6	t->1	
te na	t->4	
te ne	d->1	k->1	
te ni	 ->2	o->2	
te no	g->3	r->1	t->1	
te nu	 ->7	
te nä	m->2	r->3	
te nå	 ->1	g->26	r->1	
te nö	d->4	j->7	
te ob	e->1	
te oc	h->20	k->29	
te of	f->2	
te ol	j->1	o->1	
te om	 ->23	e->1	f->3	p->1	
te op	p->1	r->1	
te or	d->1	i->1	o->1	
te pa	l->1	r->3	
te pe	r->12	
te pl	a->2	
te po	l->1	s->1	
te pr	e->2	i->2	o->3	
te pu	n->2	
te på	 ->46	g->1	m->1	p->2	s->2	
te ra	m->6	p->3	s->2	t->1	
te re	a->4	d->3	f->1	g->19	s->6	
te ri	k->1	s->1	
te ru	b->1	
te rä	c->6	d->1	k->1	t->6	
te rå	d->11	
te rö	r->1	s->1	
te sa	g->2	k->2	m->6	n->2	t->1	
te se	 ->14	d->2	k->2	n->2	r->1	s->3	t->1	
te si	g->2	
te sj	ä->6	
te sk	a->26	e->7	i->3	j->2	u->15	y->3	ä->4	ö->1	
te sl	i->1	u->1	ä->1	
te sn	a->5	
te so	c->1	m->30	
te sp	e->1	ä->1	
te st	a->2	r->2	y->1	ä->5	å->6	ö->6	
te sv	a->2	e->1	å->1	
te sy	f->1	n->3	s->3	
te sä	g->10	k->2	l->1	n->1	r->2	t->9	
te så	 ->10	l->3	
te sö	k->1	r->3	
te ta	 ->28	c->1	g->6	l->7	n->1	r->3	s->3	
te te	c->1	k->2	n->1	
te ti	d->9	l->38	o->2	t->3	
te tj	a->1	
te to	p->1	
te tr	a->1	e->1	o->4	
te tu	m->3	
te tv	e->1	ä->1	
te ty	c->1	v->1	
te tä	c->6	n->2	
te un	d->9	i->3	
te up	p->39	
te ur	s->1	
te ut	 ->4	a->5	e->3	f->5	g->5	k->1	n->2	s->2	t->1	v->10	ö->2	
te va	d->5	l->1	r->55	
te ve	c->5	r->6	t->2	
te vi	 ->65	,->1	d->7	l->5	n->1	s->3	
te vo	r->2	
te vä	g->1	l->1	n->3	r->3	x->1	
te vå	n->1	r->2	
te äg	n->2	t->1	
te än	 ->2	.->1	d->9	n->2	t->3	
te är	 ->76	
te äv	e->5	
te ål	ä->1	
te år	e->16	
te ås	t->1	
te åt	 ->1	e->6	f->3	g->1	
te ök	a->4	
te ön	s->2	
te öp	p->2	
te öv	e->14	
te!De	t->1	
te!Me	n->1	
te, a	l->1	t->2	v->1	
te, d	e->2	
te, e	f->1	n->1	
te, f	ö->2	
te, g	a->1	
te, h	e->1	u->1	
te, i	 ->1	
te, k	a->1	o->1	
te, l	i->1	
te, m	e->2	
te, n	ä->1	
te, o	c->5	m->1	
te, p	r->1	
te, r	ö->1	
te, s	o->1	ä->1	
te, v	a->1	i->2	å->2	
te, ä	r->3	
te- o	c->1	
te-Le	 ->1	
te. D	e->1	
te.. 	P->1	
te.Ak	t->1	
te.An	n->1	
te.Be	s->1	
te.De	n->1	s->2	t->6	
te.Dä	r->1	
te.Fr	å->1	
te.Fö	r->2	
te.He	r->3	
te.I 	s->1	
te.Ja	g->5	
te.Ko	m->1	
te.Li	k->1	
te.Lä	g->1	
te.Lå	t->1	
te.Ma	l->1	
te.Me	n->1	r->1	
te.Ni	 ->1	
te.Om	 ->1	
te.På	 ->1	
te.Re	f->1	
te.Rå	d->1	
te.So	m->1	
te.Så	l->1	
te.Up	p->1	
te.Va	r->1	
te.Vi	 ->3	d->1	
te.Vå	r->1	
te.Å 	a->1	
te.År	 ->1	
te.Åt	g->1	
te: V	i->1	
te: v	a->1	
te?Fö	r->1	
te?Hu	r->1	
te?Hä	r->1	
te?I 	f->1	
te?So	m->1	
teate	r->1	
teau 	f->1	
teau,	 ->2	
tebas	e->1	
tebes	t->2	
tebet	a->12	
tebor	g->1	
tecke	n->15	
teckn	a->29	i->3	
tedel	 ->2	a->1	
tedt 	o->2	
tedt,	 ->2	
teend	e->3	
teenh	e->5	
teeri	n->1	
tefel	 ->1	
tefri	a->1	
tefrå	g->2	
teför	e->5	v->1	
teg a	t->1	
teg b	o->1	
teg f	r->6	ö->5	
teg g	j->1	
teg h	a->1	ä->1	
teg i	 ->13	
teg j	ä->1	
teg l	ä->2	
teg m	o->4	
teg n	ä->2	
teg o	c->2	
teg p	å->3	
teg s	o->7	
teg t	i->3	
teg u	n->1	
teg v	i->1	
teg, 	d->1	o->1	u->1	
teg.D	e->2	
tegen	 ->5	
teget	 ->1	,->1	
tegi 	f->5	h->1	i->1	k->1	m->1	o->2	s->4	t->2	
tegi,	 ->3	
tegi.	D->1	F->1	J->1	
tegie	r->14	
tegin	 ->5	.->2	s->1	
tegip	l->1	
tegis	k->17	
tegor	i->8	
tegra	t->16	
tegre	r->23	
tegri	t->3	
tegån	g->1	
tein.	J->1	
teinc	i->1	
teins	p->1	
teken	 ->1	s->1	
tekni	k->13	s->36	
tekno	l->3	
tekon	o->1	
tekti	o->4	
tel 2	.->1	
tel 4	 ->1	
tel i	 ->3	
tel o	m->1	
tela 	o->1	
tela,	 ->1	
telef	o->1	
telek	o->3	
telen	ä->1	
telev	e->1	i->1	
telig	e->1	
tell-	 ->3	
tella	m->1	
tellb	e->1	i->1	
telle	k->3	r->1	
tellf	ö->3	
telli	g->5	s->2	t->1	
tellm	y->1	
tellr	ä->4	
tellt	;->1	
teln 	"->1	
telse	 ->7	,->1	k->2	n->7	r->14	
telt.	D->1	
teläm	n->3	
telät	t->1	
tem -	 ->1	
tem a	l->1	v->2	
tem d	ä->3	
tem e	n->1	
tem f	u->1	ö->20	
tem g	r->1	
tem i	 ->3	n->2	
tem k	a->1	o->1	
tem m	e->8	o->1	å->1	
tem o	c->6	m->1	
tem p	å->3	
tem s	k->1	o->15	
tem ä	r->1	
tem ö	v->1	
tem, 	d->1	f->1	h->1	i->1	k->1	m->2	o->1	s->1	
tem. 	D->1	
tem.D	e->3	
tem.E	u->1	
tem.G	e->1	
tem.H	e->2	
tem.M	a->1	
tem.T	y->1	
tem.U	r->1	
tem: 	d->1	
tema,	 ->1	
temal	a->1	
teman	 ->3	.->1	n->1	
temat	 ->1	i->11	
tembe	r->15	
temen	 ->9	,->2	.->1	t->9	
temet	 ->49	)->1	,->6	.->12	?->1	
temot	 ->27	
tempe	r->4	
tempo	r->2	
temän	 ->17	,->1	.->1	d->3	n->12	s->3	
ten (	m->1	
ten -	 ->10	
ten 1	9->2	
ten A	B->1	n->1	r->1	
ten B	e->2	
ten I	 ->1	s->2	
ten L	o->1	
ten P	a->1	
ten R	e->1	
ten S	o->1	
ten a	l->1	n->2	t->61	v->69	
ten b	a->2	e->5	l->2	ä->1	
ten d	e->6	i->1	r->1	ä->1	å->1	ö->1	
ten e	f->4	l->3	n->3	t->1	u->1	
ten f	i->3	o->3	r->19	å->5	ö->59	
ten g	e->5	i->1	j->2	o->1	r->2	ä->9	ö->2	
ten h	a->20	e->2	o->5	y->1	å->1	ö->1	
ten i	 ->64	n->24	
ten j	u->1	
ten k	a->9	l->1	o->10	r->1	
ten l	i->1	ä->1	å->1	
ten m	a->2	e->23	i->2	o->2	y->2	å->10	ö->1	
ten n	a->1	e->1	u->1	y->2	ä->2	å->2	
ten o	c->53	f->1	l->1	m->55	u->1	
ten p	e->1	l->2	r->2	u->1	å->29	
ten r	e->2	u->1	ö->1	
ten s	a->2	e->1	j->2	k->25	l->1	o->15	p->1	t->10	y->1	ä->2	å->3	
ten t	a->2	i->20	o->3	r->2	
ten u	n->7	p->3	t->5	
ten v	a->8	e->3	i->18	ä->1	
ten ä	r->32	
ten å	r->1	t->5	
ten ö	k->2	v->7	
ten! 	E->1	J->1	M->1	N->1	
ten" 	s->1	
ten".	D->2	O->1	
ten) 	(->1	h->1	z->1	
ten, 	"->1	E->1	J->1	V->1	a->6	b->2	d->6	e->6	f->13	h->2	i->3	j->2	k->2	l->2	m->4	n->3	o->14	p->2	r->1	s->19	t->5	u->5	v->7	ä->4	
ten. 	J->1	L->1	
ten."	 ->1	
ten.A	l->2	r->2	
ten.D	e->43	ä->2	
ten.E	U->1	n->3	t->1	u->3	
ten.F	E->1	ö->8	
ten.H	a->1	e->6	ä->2	
ten.I	 ->2	n->2	
ten.J	a->16	
ten.K	a->2	o->4	
ten.L	å->1	
ten.M	a->1	e->7	o->1	ä->1	å->1	
ten.N	a->1	i->2	u->1	
ten.O	c->6	m->4	r->1	
ten.P	r->1	
ten.R	ä->1	
ten.S	i->1	l->2	o->1	t->1	y->1	ä->2	å->1	
ten.T	h->1	y->2	
ten.U	n->1	
ten.V	a->1	i->16	
ten.Ä	r->1	
ten.Å	 ->2	
ten.Ö	g->1	
ten: 	d->1	j->1	
ten; 	a->1	f->1	
ten?J	a->1	
ten?K	o->1	
tenFr	å->1	
tenHe	r->1	
tenNä	s->1	
tena 	e->1	i->3	m->3	
tenar	:->1	n->2	
tenbe	t->4	
tenda	 ->1	
tende	l->1	n->11	r->2	
tendr	a->1	
tendö	v->1	
tenen	 ->1	
tener	 ->7	-->10	N->1	
tenfö	r->2	
tenhe	t->3	
tenko	l->1	
tenlö	s->1	
tenpr	o->1	
tenre	n->1	s->1	
tens 	V->1	a->1	b->10	f->4	g->2	h->3	i->1	j->1	k->4	l->2	m->2	n->3	o->8	p->3	r->6	s->8	t->1	u->4	v->5	ä->1	å->1	ö->1	
tens,	 ->4	
tens.	I->1	J->1	
tensb	e->1	
tense	r->1	
tensi	f->3	t->1	v->8	
tensk	a->72	
tent 	e->1	o->1	s->1	
tenta	 ->2	t->5	
tenti	a->3	e->3	o->1	
tenvä	g->8	
teore	t->2	
tepol	i->1	
tepro	d->1	
ter (	i->1	
ter -	 ->14	
ter 1	9->1	
ter A	m->2	
ter B	a->2	
ter C	o->1	
ter E	G->1	h->1	r->1	u->2	x->1	
ter F	a->1	
ter G	A->1	a->2	o->1	u->2	
ter H	e->1	
ter J	o->1	
ter K	i->1	
ter L	i->1	
ter M	a->2	
ter O	F->1	s->1	
ter S	e->2	
ter T	a->2	
ter a	c->1	k->2	l->2	n->7	r->2	t->68	v->27	
ter b	a->3	e->8	i->1	l->1	o->1	r->1	ö->1	
ter d	e->52	i->1	o->2	r->1	y->1	ä->4	å->1	
ter e	f->2	g->2	l->10	n->15	t->8	x->1	
ter f	a->1	i->2	o->2	r->20	u->1	å->6	ö->36	
ter g	e->5	r->2	å->3	ö->3	
ter h	a->21	o->2	u->2	y->1	ä->1	å->1	
ter i	 ->55	g->2	n->23	
ter j	a->7	o->1	ä->1	
ter k	a->6	l->1	o->13	r->1	v->1	ä->1	
ter l	a->1	e->1	i->2	u->1	y->1	ä->1	å->2	
ter m	a->2	e->22	i->12	o->5	y->1	å->6	ö->1	
ter n	a->1	i->1	ä->5	å->1	
ter o	c->103	l->1	m->19	r->3	s->7	
ter p	l->1	r->1	å->32	
ter r	e->4	ä->1	å->1	ö->3	
ter s	a->5	e->2	i->7	k->18	n->1	o->94	p->1	t->7	v->1	å->9	
ter t	a->5	i->28	o->2	r->5	
ter u	n->5	p->5	r->1	t->7	
ter v	a->14	e->1	i->12	ä->3	å->2	
ter Ö	s->1	
ter ä	n->7	r->19	v->3	
ter å	r->5	t->1	
ter ö	k->1	n->1	v->10	
ter! 	D->4	E->1	J->1	L->1	P->1	S->1	T->1	U->1	V->1	
ter!J	a->1	
ter!M	y->1	
ter!V	i->1	
ter" 	s->1	
ter",	 ->1	
ter) 	o->2	
ter, 	a->3	b->7	d->10	e->7	f->7	g->4	h->2	i->6	j->2	k->2	m->9	n->3	o->12	p->1	r->2	s->20	t->6	u->5	v->5	ä->1	
ter-b	i->1	
ter-k	o->1	
ter-n	a->1	
ter. 	D->1	E->1	M->1	S->1	
ter.)	 ->1	
ter..	(->1	
ter.A	v->1	
ter.B	e->1	
ter.D	e->33	o->1	ä->1	
ter.E	U->2	n->4	t->4	u->2	
ter.F	r->4	ö->7	
ter.H	a->1	e->2	ä->1	
ter.I	 ->2	n->1	
ter.J	a->21	
ter.K	o->4	
ter.L	å->3	
ter.M	e->7	i->1	
ter.N	ä->3	
ter.O	c->1	m->2	r->1	
ter.P	a->2	u->1	å->1	
ter.S	a->1	l->2	o->1	t->1	å->1	
ter.T	a->2	e->1	i->3	
ter.U	n->1	
ter.V	a->3	i->12	
ter.Ä	n->1	v->2	
ter.Å	 ->2	
ter: 	A->1	I->1	f->1	
ter; 	a->1	d->1	
ter?B	o->1	
ter?D	e->1	
ter?H	e->1	
ter?T	a->1	
terHe	r->1	
tera 	-->2	F->1	I->1	a->38	b->3	d->39	e->23	f->10	g->2	h->3	i->5	k->6	l->1	m->9	n->1	o->13	p->8	r->5	s->5	t->1	u->2	v->9	ä->2	ö->2	
tera,	 ->5	
tera.	B->1	D->2	F->1	H->2	I->1	J->4	L->2	M->2	V->1	
terad	 ->9	,->2	.->1	e->36	
teral	 ->1	a->6	t->1	
teran	-->1	b->8	d->16	v->18	
terar	 ->102	,->1	.->4	e->4	
teras	 ->51	,->2	.->11	
terat	 ->30	,->1	.->1	o->2	s->8	u->9	
terbe	t->3	
terbi	l->1	
terda	m->41	
terdö	r->1	
terer	ö->1	
terfa	r->1	
terfi	n->3	r->2	
terfr	å->8	
terfu	n->2	
terfö	l->3	r->8	
terga	v->2	
terge	 ->1	r->2	s->1	
tergi	f->2	v->6	
tergr	u->1	
tergå	t->1	
terha	n->5	
terhä	m->2	
terhå	l->2	
teri 	o->1	
teria	l->23	
terie	l->4	r->20	s->1	t->3	
terig	e->19	
teril	 ->1	
terim	s->8	
terin	 ->1	f->4	g->77	r->2	s->8	t->1	ä->3	
teris	e->2	
terko	m->7	
terkr	ä->1	
terle	v->3	
terli	g->56	
terly	s->2	
terlä	m->3	
terme	r->3	
termi	d->9	
termö	t->2	
tern 	(->1	-->1	d->1	e->1	g->1	h->1	i->1	k->3	m->1	n->1	o->6	r->1	s->2	t->1	u->1	v->2	ä->1	
tern,	 ->2	
tern.	)->1	D->4	H->1	J->2	Ö->1	
tern/	N->2	
terna	 ->339	"->1	,->68	.->70	:->3	;->1	?->4	s->75	t->91	
terne	r->1	t->10	
ternf	r->1	
terni	v->1	
terns	 ->5	
ternt	 ->3	.->1	
terom	r->1	
terpa	r->1	
terpo	s->2	
terpr	e->1	
terra	n->2	
terre	g->3	s->1	z->1	
terri	k->130	t->17	
terro	r->10	
terrå	d->14	
ters 	a->3	b->4	i->1	k->1	r->2	u->1	v->1	
ters-	b->1	
tersa	m->1	t->3	
terse	n->1	
tersk	a->4	r->1	
terso	m->190	
tersp	e->3	
terst	 ->18	a->15	r->12	ä->13	å->14	
tert 	o->2	
terta	 ->2	g->6	n->3	s->1	
tertr	a->1	ä->1	
tertä	n->1	
terup	p->34	
terve	n->7	r->1	
tervi	n->66	
tervj	u->3	
tervu	n->2	
tervä	n->3	r->1	
teråt	 ->1	
tes 3	,->1	
tes a	l->1	v->3	
tes e	n->1	
tes i	 ->4	h->1	n->1	
tes m	e->1	o->1	
tes t	i->1	
tes u	p->1	
tes, 	e->1	
tes- 	o->1	
tes.F	l->1	
tes.K	o->1	
tes.O	m->1	
tes.V	i->1	
tesat	s->1	
tesek	t->2	
tesen	 ->1	
tesgå	 ->2	s->1	
tesis	k->3	
teslu	t->17	
teslö	t->2	
tess 	n->1	o->1	r->1	s->1	
tessb	e->5	
tesse	n->2	
tessh	ä->1	
test 	f->1	m->1	n->1	
test,	 ->1	
testa	n->2	
teste	n->1	r->5	
testä	n->4	
testå	e->1	
tesys	t->1	
tet (	f->1	
tet ,	 ->1	
tet -	 ->7	
tet 1	9->2	
tet K	u->1	
tet M	o->1	
tet a	c->1	l->2	n->10	r->1	t->43	v->48	
tet b	a->2	e->8	l->3	ä->1	ö->6	
tet c	h->1	i->1	
tet d	e->9	i->2	r->1	ä->2	å->2	
tet e	f->3	l->3	n->3	x->1	
tet f	a->1	i->1	o->2	r->8	u->1	å->2	ö->144	
tet g	e->4	i->1	o->7	r->3	ö->2	
tet h	a->34	e->1	o->2	ä->2	ö->1	
tet i	 ->43	b->1	n->29	
tet j	u->3	
tet k	a->8	o->16	r->4	u->3	
tet l	a->1	e->1	i->1	y->1	ä->5	
tet m	e->45	o->4	ä->1	å->9	
tet n	o->1	u->4	ä->1	
tet o	c->74	f->1	k->1	m->29	r->3	
tet p	o->1	å->14	
tet r	e->3	å->1	ö->1	
tet s	a->1	e->4	i->1	j->1	k->11	n->1	o->17	p->3	t->7	ä->3	å->5	
tet t	i->10	v->1	y->1	ä->1	
tet u	n->3	p->2	t->4	
tet v	a->2	e->2	i->11	ä->2	
tet ä	n->3	r->22	v->2	
tet å	t->1	
tet!H	e->1	
tet",	 ->1	
tet".	J->1	
tet, 	C->1	G->1	I->1	a->6	d->10	e->5	f->1	g->2	h->3	i->6	k->5	m->10	n->2	o->10	p->1	r->1	s->10	t->1	u->2	v->9	ä->2	å->1	ö->1	
tet- 	o->1	
tet. 	D->1	
tet.)	A->1	B->2	
tet..	.->1	
tet.B	r->1	
tet.D	e->24	ä->2	å->1	
tet.E	f->1	n->1	u->2	
tet.F	l->1	r->2	ö->4	
tet.H	a->1	e->5	i->1	
tet.I	 ->3	
tet.J	a->15	
tet.K	o->2	u->1	
tet.L	i->1	
tet.M	a->2	e->2	
tet.N	ä->1	
tet.P	o->1	
tet.R	ä->1	
tet.S	o->1	å->2	
tet.T	a->1	
tet.V	a->1	i->7	å->1	
tet.Ä	v->1	
tet: 	"->1	d->1	e->1	ö->1	
tet?D	e->1	
tet?H	e->1	u->1	
tet?N	ä->1	
tet?Ä	r->1	
teten	 ->44	,->4	.->6	:->1	s->1	
teter	 ->9	.->1	n->9	s->1	
tetis	k->2	
tets 	-->1	a->5	b->10	d->8	e->1	f->11	g->3	h->2	k->2	l->8	m->3	o->17	p->2	r->6	s->15	t->9	u->5	v->1	y->3	ä->2	ö->2	
tets-	 ->1	
tetsa	r->2	
tetsb	e->3	
tetsf	i->1	r->1	
tetsg	a->1	
tetsh	a->2	
tetsk	l->1	r->2	
tetsn	o->1	
tetso	m->1	
tetsp	a->4	r->15	
tetsr	e->3	
tetss	a->1	p->1	
teuro	p->9	
text 	a->1	f->1	i->1	k->1	l->1	o->2	s->5	
text,	 ->5	
text.	M->1	
texte	n->17	r->10	
tfall	e->7	
tfara	n->89	
tfart	y->1	
tfasn	i->3	
tfatt	a->2	
tfede	r->1	
tflag	g->1	
tfler	 ->1	
tflir	t->1	
tflyt	t->1	
tform	a->15	n->26	
tfors	k->1	
tfram	t->1	
tfråg	a->1	n->7	o->8	
tfull	 ->2	a->8	t->5	
tfäll	i->8	
tfärd	a->12	i->8	
tfäst	e->2	
tfång	a->1	
tfölj	a->9	d->1	e->1	t->1	
tför 	a->1	b->3	d->5	e->1	f->3	h->1	k->1	l->4	m->4	o->12	s->9	t->2	
tföra	 ->14	.->2	n->1	s->1	
tförb	u->1	
tförd	,->1	a->1	e->2	r->3	
tföre	b->1	
tförf	a->2	
tförk	l->7	
tförl	i->3	u->1	
tföro	r->6	
tförs	 ->3	l->1	t->1	
tfört	 ->4	,->2	s->7	
tförä	n->4	
tgavs	 ->1	
tgick	 ->1	
tgift	e->11	s->5	
tgilt	i->8	
tgivi	t->1	
tgivn	a->1	
tgjor	d->4	
tgrup	p->7	
tgärd	 ->13	,->6	.->5	;->1	a->3	e->207	s->10	
tgå e	n->1	
tgå f	r->2	
tgå t	i->1	
tgå.D	ä->1	
tgå.N	ä->1	
tgåen	d->14	
tgång	 ->2	a->1	e->4	s->11	
tgår 	f->2	h->1	i->2	j->1	o->2	
tgåvo	r->1	
tgör 	"->1	3->1	8->1	a->1	d->6	e->15	f->2	g->3	h->1	i->1	k->1	m->1	n->2	p->1	r->1	s->3	t->2	u->1	v->1	y->1	
tgör,	 ->1	
tgör.	D->1	
tgöra	 ->11	n->2	
tgörs	 ->2	
th Sc	h->1	
th ha	r->1	
th nä	m->1	
th oc	h->1	
th, o	r->1	
th-Be	h->7	
thand	l->1	
thant	e->1	
thar 	e->1	v->1	
thar"	 ->1	
thava	r->1	
the R	o->1	
the c	i->1	
the i	m->1	
then 	f->2	h->1	
then,	 ->1	
thens	 ->2	
ther"	 ->1	
thera	n->1	
thet 	o->1	s->1	
thet.	D->1	
thete	n->1	
thets	n->1	
thies	 ->2	
thom 	P->3	
thu o	c->1	
thuse	f->3	
thusg	a->4	
thy o	c->1	
thäls	n->1	
thärd	a->1	l->3	
thåll	a->8	e->1	n->1	s->1	
thöra	n->1	
ti - 	a->1	
ti an	s->1	
ti de	l->1	t->1	
ti fr	å->1	
ti fö	r->9	
ti gj	o->1	
ti ha	r->3	
ti he	m->1	
ti i 	E->1	d->1	e->1	s->1	Ö->1	
ti ig	e->1	
ti in	g->2	n->1	
ti ko	m->2	
ti kr	ä->1	
ti me	d->2	
ti oc	h->11	
ti om	 ->1	
ti på	 ->2	
ti sn	a->1	
ti so	m->7	
ti så	 ->1	
ti ti	l->2	
ti up	p->1	
ti va	d->1	
ti åt	e->1	
ti! J	a->1	o->1	
ti! U	p->1	
ti" s	o->1	
ti, M	i->1	
ti, b	r->1	
ti, d	e->2	
ti, e	n->1	
ti, k	a->1	
ti, l	i->1	
ti, m	e->1	
ti, o	c->1	
ti, p	r->1	
ti, s	k->1	o->1	
ti, ä	r->1	v->1	
ti-ge	m->1	
ti-ir	l->1	
ti-ra	s->1	
ti...	(->1	
ti.De	 ->1	n->1	t->1	
ti.Ef	t->1	
ti.En	 ->1	
ti.Fo	l->1	
ti.Ha	i->1	
ti.He	r->1	
ti.Hä	r->1	
ti.I 	k->1	
ti.Ja	g->1	
ti.Ka	n->1	
ti.Ku	l->1	
ti.Mi	n->1	
ti.Vi	 ->1	
tial 	m->1	
tial,	 ->1	
tial.	F->1	
tian 	1->1	
tiati	v->80	
tibed	r->1	
tibet	a->10	
tical	 ->1	
tice 	d->4	
tiche	r->1	
tick 	i->1	
ticke	t->1	
tickp	r->3	
tid E	U->1	
tid a	l->1	n->2	t->24	v->2	
tid b	a->1	e->3	l->2	ä->1	ö->4	
tid c	a->1	
tid d	e->5	r->1	ä->1	å->3	
tid e	f->1	n->4	t->3	
tid f	i->2	r->1	u->1	y->1	å->2	ö->11	
tid g	j->2	ö->1	
tid h	a->11	e->1	i->1	ä->1	ö->2	
tid i	 ->5	n->9	
tid j	a->1	
tid k	a->5	l->1	o->1	r->2	
tid l	a->1	ä->2	
tid m	e->2	i->1	o->1	y->1	ä->1	å->1	
tid n	a->2	o->1	ä->1	å->1	
tid o	c->4	e->1	m->1	p->1	
tid p	r->1	å->3	
tid r	ä->1	å->1	
tid s	e->1	j->1	k->3	l->1	o->4	t->2	y->1	ä->1	å->2	
tid t	a->3	i->4	v->1	
tid u	n->2	
tid v	a->2	i->4	
tid y	r->1	
tid ä	n->2	r->8	v->1	
tid å	t->3	
tid, 	d->1	e->1	f->1	h->1	i->2	m->1	o->4	p->1	v->3	ä->1	
tid..	 ->1	
tid.D	e->5	
tid.F	ö->1	
tid.K	o->1	
tid.M	a->1	
tid.N	ä->1	
tid.O	m->1	
tid.S	o->1	
tid.T	a->1	i->1	
tid.V	i->1	
tid: 	d->1	
tida 	E->1	a->1	b->3	d->1	e->2	f->3	h->1	k->1	p->1	r->1	s->2	t->4	v->1	å->1	
tidem	o->1	
tiden	 ->74	,->7	.->31	:->1	?->2	s->3	
tider	 ->3	,->2	
tidig	a->80	t->72	
tidli	g->4	
tidni	n->6	
tidpu	n->10	
tidsa	r->4	
tidsb	e->2	
tidsd	i->3	u->1	
tidsf	r->10	ö->1	
tidsg	r->1	
tidsi	n->2	
tidsm	ä->2	
tidso	r->1	
tidsp	e->10	l->5	
tidsr	a->5	y->2	
tidss	k->1	y->1	
tidså	l->2	t->1	
tidsö	d->1	
tidta	b->6	
tie- 	o->1	
tiebö	r->1	
tiede	p->2	
tielf	t->1	
tiell	 ->1	a->9	
tiemi	n->3	
tient	 ->1	e->3	
tier 	f->7	h->2	m->1	o->3	r->1	s->2	u->1	
tier,	 ->2	
tiera	d->1	t->2	
tieri	n->4	
tiern	a->12	
tiet 	(->3	e->1	o->1	r->1	
tiet)	 ->1	,->2	.->1	
tiet,	 ->4	
tietn	i->3	
tiets	 ->16	
tieur	o->1	
tieäg	a->2	
tifas	c->3	
tific	e->13	i->2	
tifie	r->16	
tifik	a->4	
tifiq	u->1	
tifol	k->1	
tifon	d->2	
tifrå	g->1	n->17	
tifta	 ->4	n->5	r->5	t->1	
tiftn	i->113	
tig -	 ->1	,->1	
tig b	e->2	r->1	
tig d	e->6	i->1	
tig e	x->1	
tig f	r->10	u->2	ö->8	
tig g	l->1	r->2	
tig h	j->1	ä->2	
tig i	.->1	n->3	
tig j	u->1	
tig k	a->1	o->2	r->1	u->1	
tig l	e->1	ö->2	
tig m	e->1	i->2	å->1	ö->1	
tig o	c->10	r->1	
tig p	o->1	u->7	å->2	
tig r	a->1	e->3	o->8	
tig s	a->1	e->1	i->1	t->1	
tig t	e->1	i->3	r->1	
tig u	p->1	t->4	
tig å	t->3	
tig ö	k->1	v->1	
tig, 	b->1	f->1	g->1	l->1	o->1	s->2	u->1	
tig.D	e->4	
tig.I	 ->1	
tig.J	a->3	
tig.M	a->1	e->1	
tig.N	a->1	
tig?J	o->1	
tiga 	"->1	-->1	E->1	a->7	b->10	d->5	e->5	f->26	i->14	k->4	l->2	m->5	n->2	o->11	p->2	r->4	s->13	t->7	u->1	v->6	ä->4	
tiga,	 ->6	
tiga.	A->1	O->1	V->1	
tigad	,->1	.->2	e->7	
tigan	d->2	
tigar	e->17	
tigas	 ->2	t->46	
tigat	 ->8	,->2	
tigdo	m->12	
tiger	 ->2	.->1	n->1	
tigge	r->1	
tighe	t->182	
tigit	 ->1	.->1	
tigli	g->4	
tigma	t->1	
tigt 	-->1	R->1	a->66	b->4	d->3	e->2	f->18	g->2	h->3	i->7	k->3	l->1	m->9	n->4	o->14	p->2	r->1	s->13	t->4	u->3	v->3	y->1	ä->2	
tigt,	 ->17	
tigt.	A->1	D->1	E->1	F->2	J->1	L->1	N->1	S->1	V->4	
tihop	,->1	
tiint	r->1	
tik -	 ->2	
tik J	ö->1	
tik a	n->1	v->4	
tik e	g->1	l->1	n->1	
tik f	i->1	r->1	å->1	ö->16	
tik h	a->2	u->1	ö->1	
tik i	 ->6	n->1	
tik k	a->2	u->1	
tik m	e->5	o->3	å->2	ö->1	
tik n	ä->1	
tik o	c->25	m->2	r->1	
tik p	å->2	
tik r	e->1	ö->1	
tik s	o->28	
tik t	i->1	
tik u	n->1	p->1	
tik v	a->1	i->2	
tik ä	r->4	
tik ö	v->1	
tik!O	m->1	
tik" 	o->1	
tik, 	d->6	e->2	f->2	h->1	i->1	m->1	n->2	o->1	s->2	t->10	v->3	
tik..	(->1	
tik.D	e->6	ä->1	å->1	
tik.E	n->1	u->1	
tik.F	r->1	ö->1	
tik.H	a->1	i->1	ä->1	
tik.I	 ->1	
tik.J	a->1	
tik.M	e->1	
tik.R	e->1	i->1	
tik.T	v->1	
tik.V	i->2	
tik.Ä	v->1	
tik?H	e->1	
tik?V	a->1	
tika 	f->2	i->1	
tikab	e->1	
tikaf	r->1	
tikal	a->3	
tikan	 ->1	
tikap	r->1	
tikas	m->1	
tikel	 ->93	,->2	
tiken	 ->77	,->20	.->27	?->2	H->1	s->17	
tiker	 ->8	.->1	n->6	s->1	
tikla	r->15	
tikol	o->1	
tikom	r->6	
tikra	t->1	
tikry	p->2	
tiks 	m->1	
til -	 ->1	
til m	e->1	
til n	ä->1	
tilat	e->1	
tiled	a->1	
tiler	a->1	
tilis	m->1	
till 	"->1	-->1	1->5	2->4	3->2	4->1	5->1	7->3	8->2	9->4	A->1	B->5	C->2	D->1	E->32	F->7	G->2	K->13	L->2	M->3	N->2	O->1	P->5	R->1	S->7	T->5	V->1	W->4	a->298	b->37	c->1	d->267	e->187	f->133	g->31	h->45	i->22	j->5	k->64	l->13	m->72	n->33	o->48	p->30	r->53	s->144	t->26	u->22	v->59	y->5	Ö->1	ä->10	å->10	ö->3	
till!	H->1	
till,	 ->17	
till.	A->1	D->5	E->1	F->1	H->2	I->2	R->1	S->1	
till:	 ->1	
till?	D->1	H->1	J->1	
tilla	 ->1	
tillb	a->52	r->4	
tilld	e->12	r->1	
tille	r->3	
tillf	o->6	r->27	ä->97	ö->13	
tillg	o->1	r->2	ä->21	å->25	
tillh	a->43	e->2	ö->8	
tillk	o->6	ä->9	
tillm	ä->2	ö->3	
tilln	ä->6	
tillr	ä->77	
tills	 ->42	,->2	.->3	?->1	a->31	e->13	k->5	l->1	t->22	v->3	ä->4	
tillt	a->3	r->8	
tillv	a->1	e->84	i->1	ä->28	
tillä	g->20	m->174	
tillå	t->45	
tima 	f->1	i->1	o->2	s->1	
tima,	 ->1	
tima.	H->1	
timal	 ->2	a->1	
timat	u->1	
timer	a->4	i->1	
timet	e->1	
timis	t->4	
timit	e->6	
timma	r->6	
timme	 ->5	
timt 	i->1	o->2	
timt,	 ->1	
timul	a->4	e->7	
timög	e->1	
tin a	t->2	
tin b	e->1	
tin f	ö->2	
tin h	a->1	
tin i	n->1	
tin m	o->1	
tin o	c->3	
tin s	o->2	å->1	
tin v	u->1	
tin, 	f->1	m->1	
tin.A	l->1	
tin.F	ö->2	
tin.H	e->1	
tin.O	m->1	
tina 	a->1	f->1	o->3	s->1	
tina-	I->1	
tinaf	l->1	r->1	
tinas	 ->1	
tinat	i->5	
tindu	s->2	
tinen	,->1	t->5	
tiner	 ->6	
tinez	 ->1	
ting 	-->1	a->9	b->1	d->1	f->6	g->1	h->5	k->3	l->1	m->8	n->1	o->1	p->1	s->11	t->1	u->1	v->4	ä->4	å->2	
ting,	 ->4	
ting.	D->4	
tinga	r->12	
tinge	l->1	n->10	t->2	
tingf	o->1	
tinie	r->4	
tinkt	e->1	i->2	
tinmä	s->1	
tinne	h->1	
tinno	v->1	
tinos	 ->2	,->2	
tinot	t->1	
tinri	k->2	
tins 	a->1	p->1	s->2	v->1	
tinsk	 ->1	a->7	
tinue	r->2	
tinve	s->1	
tio f	a->1	
tio g	r->1	å->2	
tio m	i->2	
tio s	i->1	
tio ä	n->1	
tio å	r->7	
tioel	v->1	
tiofe	m->1	
tion 	(->5	-->3	1->5	5->1	A->1	I->1	a->22	b->3	d->6	e->1	f->17	g->4	h->5	i->23	j->1	k->5	m->11	n->3	o->42	p->9	s->45	t->18	u->3	v->7	ä->4	
tion"	 ->1	
tion,	 ->36	
tion.	 ->1	1->1	B->1	D->11	E->2	F->2	H->5	I->5	J->8	K->1	M->3	N->1	O->2	S->3	T->2	V->8	Å->1	
tion:	 ->3	
tion;	 ->1	
tion?	 ->1	J->1	K->1	
tiona	l->46	
tiond	e->1	
tione	l->274	n->180	r->306	
tioni	s->5	
tions	 ->1	-->2	a->12	b->2	d->1	f->18	h->8	i->1	k->11	l->1	m->5	n->1	p->10	r->3	s->14	t->2	u->3	v->1	
tiopi	e->3	
tiosj	u->1	
tiota	l->6	
tiotu	s->1	
tipen	d->1	
tipro	g->2	
tique	 ->1	s->1	
tiref	o->1	
tis d	ä->1	
tis e	l->1	
tis i	n->1	
tis r	a->1	
tis t	i->1	
tis u	t->1	
tis å	t->1	
tis, 	d->1	
tis.D	e->1	
tisda	g->2	
tisek	t->2	
tisem	i->3	
tiser	a->15	i->2	
tish 	P->1	
tisk 	a->2	b->6	d->8	f->5	g->3	h->1	i->5	k->8	l->4	m->4	n->3	o->5	p->6	r->8	s->16	t->5	u->9	v->2	ö->1	
tisk,	 ->2	
tisk-	s->1	
tisk.	 ->1	H->1	I->3	J->1	M->1	
tiska	 ->308	,->7	.->1	
tiskt	 ->148	!->1	,->6	.->6	
tism 	i->1	o->1	
tism,	 ->2	
tism.	D->1	H->1	N->1	
tispl	i->1	
tisti	k->6	s->3	
tisys	t->1	
tit a	r->1	t->1	
tit e	t->1	
tit f	ö->1	
tit m	o->1	
tit s	i->2	
titat	i->4	
titel	n->1	
titet	 ->4	,->1	.->1	s->2	
titie	-->1	d->2	m->3	
titio	n->1	
titru	s->1	
tits 	a->1	f->1	n->1	p->1	u->4	
titt 	p->2	
titta	 ->13	n->1	r->6	
titue	r->1	
titut	i->158	
tityd	 ->4	.->1	
tiv (	K->1	
tiv -	 ->3	
tiv 9	3->1	4->2	6->5	
tiv E	n->1	
tiv a	n->3	t->2	v->1	
tiv b	a->1	e->1	
tiv d	e->2	i->2	
tiv e	f->1	k->2	n->4	
tiv f	a->1	r->4	å->2	ö->9	
tiv g	e->1	
tiv h	a->7	j->1	
tiv i	 ->5	m->1	n->7	
tiv k	a->3	o->7	
tiv l	a->2	e->1	i->3	ö->1	
tiv m	e->2	i->1	o->1	å->1	
tiv o	c->8	m->21	p->1	
tiv p	o->1	å->7	
tiv r	e->1	i->1	o->1	
tiv s	a->1	e->2	k->2	n->1	o->25	t->7	y->3	å->4	
tiv t	i->14	r->1	
tiv u	t->3	
tiv v	e->1	i->4	ä->1	
tiv ä	n->1	r->5	
tiv å	t->2	
tiv ö	v->1	
tiv, 	9->1	a->1	b->1	d->3	e->1	h->1	i->1	j->1	l->1	m->2	n->1	o->5	s->3	u->1	
tiv. 	V->1	
tiv..	H->1	
tiv.A	t->1	
tiv.B	l->1	
tiv.D	e->4	å->1	
tiv.E	n->1	
tiv.F	ö->4	
tiv.I	 ->1	n->1	
tiv.L	å->1	
tiv.M	e->1	
tiv.O	m->1	
tiv.R	i->1	
tiv.S	å->1	
tiv.V	i->1	
tiv.Y	t->1	
tiv: 	F->1	v->1	
tiv; 	a->1	
tiv?F	ö->1	
tiv?N	e->1	
tiva 	a->4	b->8	c->1	d->3	e->5	f->8	h->2	i->5	k->9	l->1	m->3	n->1	o->12	p->8	r->9	s->9	t->9	v->3	å->4	ö->1	
tiva,	 ->4	
tiva.	A->1	H->1	V->1	
tivan	d->1	
tivar	e->11	
tivas	t->1	
tivat	i->1	
tivav	t->7	
tivbe	t->1	
tive 	E->1	a->1	b->2	d->1	f->1	k->2	l->1	m->2	p->3	t->1	
tiven	 ->8	,->2	.->1	s->1	
tiver	a->14	i->3	
tivet	 ->69	,->10	.->14	s->7	
tivfö	r->4	
tivis	e->3	m->1	
tivit	e->38	
tivli	s->2	
tivri	k->1	
tivrä	t->4	
tivt 	-->1	a->9	b->4	d->1	e->1	f->5	h->1	i->5	k->3	m->4	n->1	o->15	p->4	r->4	s->29	t->6	u->1	v->1	y->1	ä->1	å->2	ö->1	
tivt,	 ->7	
tivt.	 ->1	D->2	E->1	I->1	P->1	Ä->1	
tiös 	d->1	u->1	
tiös,	 ->1	
tiösa	 ->5	.->1	r->2	
tiöst	 ->1	
tja a	l->4	r->1	
tja c	h->1	
tja d	e->4	i->1	
tja i	 ->1	
tja o	c->1	
tja s	a->1	i->1	t->3	
tjade	 ->2	s->2	
tjand	e->9	
tjar 	a->1	d->1	m->1	
tjas 	a->1	f->3	i->1	s->1	
tjat 	m->1	
tjata	 ->1	
tjock	 ->1	a->1	
tjugo	 ->2	f->1	n->1	
tjust	 ->1	
tjämn	a->3	i->2	
tjämt	 ->2	.->1	
tjäna	 ->4	d->1	r->16	
tjäns	t->123	
tjänt	 ->2	a->27	
tjära	.->1	
tjärn	a->2	
tkant	e->1	
tkast	 ->9	,->1	e->5	
tkate	g->1	
tklas	s->1	
tkom.	D->1	
tkomm	e->1	i->17	
tkomp	e->1	
tkoms	t->1	
tkonc	e->1	
tkonk	u->1	
tkont	r->16	
tkost	n->2	
tkrav	e->1	
tkrig	 ->1	
tkräv	a->1	e->2	
tkubi	k->1	
tkust	e->2	
tkväl	l->1	
tkäll	a->1	
tkött	 ->2	s->1	
tlagt	s->1	
tland	 ->3	,->3	.->2	e->4	s->3	
tlant	e->4	i->1	k->1	
tle o	c->2	
tle ä	r->1	
tle.V	i->1	
tlekt	y->1	
tler 	d->1	s->1	ä->1	
tler,	 ->1	
tler-	r->1	
tlers	 ->1	
tlevn	a->1	
tlig 	a->2	b->2	d->8	f->5	i->5	k->6	n->2	o->3	p->3	r->2	s->12	t->7	u->6	å->1	
tlig,	 ->1	
tlig.	G->1	J->1	O->1	V->1	
tlig?	D->1	
tliga	 ->180	,->4	.->3	/->1	
tlige	n->137	
tligg	j->8	ö->9	
tligh	e->37	
tligt	 ->72	,->2	.->7	
tlinj	e->76	
tlist	a->2	
tlova	d->1	t->2	
tlägg	 ->1	a->1	e->1	s->1	
tlämn	a->1	i->1	
tländ	e->12	s->3	
tlänn	i->1	
tlåta	n->2	
tlös.	D->1	
tlösa	 ->1	
tlösh	e->2	
tlöst	 ->1	
tmakt	e->1	
tmana	 ->1	
tmani	n->21	
tmarg	i->1	
tmark	n->1	
tmatc	h->1	
tmede	l->1	
tmedl	e->1	
tmer 	i->1	
tmins	t->27	
tmiss	b->1	
tmonn	ä->1	
tmynd	i->3	
tmynn	a->1	
tmäng	d->2	
tmärk	e->1	s->1	t->30	
tmäss	i->1	
tmäti	g->1	
tmåls	d->1	
tna a	t->1	
tna b	a->1	e->1	
tna d	e->1	ö->1	
tna e	n->1	
tna f	å->1	
tna h	a->1	
tna i	 ->1	
tna m	å->1	
tna o	c->2	m->16	
tna p	å->1	
tna s	ä->1	
tna t	i->2	o->2	
tna v	e->1	
tna, 	d->1	m->1	n->1	
tna. 	J->1	K->1	
tna.D	ä->1	
tna.E	f->1	
tna.S	l->1	
tna.U	n->1	
tnad 	a->1	e->1	f->3	k->1	m->1	s->2	t->1	
tnad.	J->1	
tnad;	 ->1	
tnade	n->13	r->62	
tnads	-->4	/->1	b->4	e->4	f->5	i->2	p->1	u->1	
tnar 	a->1	d->1	i->4	o->2	
tnas 	g->1	p->1	
tnas.	D->1	
tne o	m->1	
tne t	i->1	
tnen 	o->1	
tnen,	 ->1	
tnen.	J->1	
tner 	-->1	i->3	o->3	
tner.	D->1	
tner?	K->1	
tnern	a->1	
tners	h->1	k->17	
tness	 ->1	
tnet 	f->1	i->1	o->1	v->1	
tnet.	 ->1	N->1	
tning	 ->221	)->1	,->42	.->44	:->1	;->2	?->1	a->68	e->165	s->103	
tnisk	 ->3	a->8	t->3	
tnjut	e->1	
tnytt	i->1	j->41	
tnämn	a->3	d->2	i->3	
tnät 	s->1	
to - 	d->1	
to ac	c->1	
to fö	r->3	
to ha	r->1	
to hå	r->1	
to i 	f->1	
to ka	n->1	
to oc	h->1	
to om	 ->1	
to sa	d->1	
to så	 ->1	
to ti	l->1	
to vi	k->1	
to öp	p->1	
to-an	a->1	
to-pr	o->1	
to.Ja	g->1	
to.Vi	 ->1	
to/Oi	l->1	
toakt	i->1	
toana	l->1	
tobak	,->1	s->1	
tobas	e->1	
tober	 ->8	
tobet	ä->1	
tockh	o->3	
tod a	t->2	v->2	
tod b	ö->1	
tod d	e->2	
tod e	f->2	
tod f	r->1	ö->2	
tod i	 ->1	
tod j	a->1	
tod m	e->2	y->1	
tod n	y->1	
tod p	r->1	å->1	
tod s	k->1	o->5	
tod ä	r->1	
tod å	t->1	
toden	 ->2	,->1	.->1	
toder	 ->8	,->1	.->2	n->1	
todon	t->1	
tog 1	9->1	
tog b	e->1	
tog d	e->3	
tog e	n->2	t->2	
tog h	e->1	ä->1	
tog i	 ->3	
tog k	o->3	
tog l	a->4	ä->1	
tog m	a->1	å->1	
tog n	i->1	
tog o	c->1	m->1	
tog p	a->1	
tog r	e->3	å->1	
tog s	t->1	
tog u	p->9	
togam	 ->1	,->1	
togen	a->1	t->1	
togs 	-->1	a->4	b->1	e->1	i->2	k->2	m->3	o->2	s->1	u->3	
togs,	 ->2	
tokol	l->26	
tol b	e->1	
tol d	ä->1	
tol i	 ->1	
tol o	c->1	
tol s	o->2	
tol v	i->1	
tol.D	e->1	
tol.E	t->1	
tolar	 ->12	,->1	.->2	n->8	s->2	
tolen	 ->27	,->5	.->6	s->8	
toler	a->11	e->7	
tolik	.->1	:->1	e->2	
tolka	 ->2	r->5	s->4	t->1	
tolkn	i->14	
tolpe	 ->1	
tolsa	v->1	
tolsb	u->1	
tolsf	a->1	ö->1	
tolsk	a->4	
tolsp	r->1	
tolss	y->1	
tolst	v->1	
tolsu	t->1	
tolsv	ä->1	
tolt 	ö->6	
tolta	 ->3	
tolth	e->2	
tolv 	å->1	
tom P	P->1	
tom a	l->5	n->2	t->7	v->1	
tom b	e->4	l->1	o->1	ö->3	
tom d	e->3	r->1	
tom e	f->1	t->1	
tom f	a->1	i->1	ö->5	
tom g	e->2	o->1	
tom h	a->3	ä->1	
tom i	 ->2	n->3	
tom k	a->1	o->4	r->2	u->1	
tom m	e->2	i->1	å->4	
tom n	å->2	
tom o	a->1	c->1	m->3	
tom p	o->1	å->2	
tom r	e->4	
tom s	i->1	k->2	t->3	
tom t	i->3	r->1	
tom v	i->5	
tom ä	r->4	v->1	
tom!T	r->1	
tom) 	o->1	
tom, 	d->1	f->1	h->1	n->1	s->1	
tom.V	i->1	
tomat	i->8	
tomen	e->3	
tomeu	r->3	
tomfo	r->1	
tomma	 ->1	
tomor	d->7	
tomru	m->2	
tområ	d->6	
tomst	å->2	
ton 5	7->1	
ton a	n->1	v->2	
ton f	ö->3	
ton i	 ->3	
ton k	o->1	
ton m	e->7	i->2	
ton o	c->2	l->3	
ton p	e->1	
ton s	o->1	t->2	
ton t	i->1	
ton v	e->1	
ton å	r->2	
ton, 	e->1	
ton-H	a->1	
ton. 	D->1	
ton.H	e->1	
ton.V	a->1	
ton/å	r->2	
ton? 	D->1	
tona 	a->8	d->5	e->2	h->1	i->1	n->1	o->1	s->1	t->4	v->2	
tonad	e->6	
tonar	 ->6	,->1	
tonas	 ->1	
tonat	 ->2	,->2	.->1	i->1	
tonde	 ->2	.->1	
tone 	a->2	b->1	d->1	e->1	f->1	g->1	h->1	i->5	j->1	k->2	l->1	n->4	o->1	r->1	s->1	t->1	v->2	
tonen	 ->1	
toner	 ->1	,->1	
tongi	v->1	
tonhu	n->1	
tonin	g->1	
tons 	b->1	p->1	r->1	v->1	
tonvi	k->4	
tonår	i->1	
top-s	h->1	
topil	o->1	
topp 	f->7	p->1	
toppa	 ->4	d->1	r->1	s->4	
toppe	n->3	
toppm	ö->10	
topro	t->2	
tor a	n->2	r->1	v->2	
tor b	e->11	i->2	r->2	ö->1	
tor c	h->1	
tor d	e->11	j->1	ä->1	ö->1	
tor e	l->1	n->1	r->1	u->1	
tor f	a->1	r->2	ö->6	
tor g	e->1	r->1	
tor h	a->1	j->3	ä->2	
tor i	 ->2	n->2	
tor j	o->2	
tor k	a->2	o->1	
tor l	i->1	
tor m	a->6	e->2	ä->2	å->2	
tor o	c->3	m->2	r->2	
tor p	o->2	r->1	
tor r	e->5	o->1	
tor s	o->6	y->1	
tor t	i->2	j->1	
tor u	n->1	p->5	t->10	
tor v	a->1	i->3	
tor ä	r->1	
tor ö	v->1	
tor, 	i->1	k->1	m->1	n->2	o->2	s->3	
tor.A	l->1	
tor.D	e->1	
tor.J	a->3	
tor.O	c->1	
tor.R	e->1	
tor.T	y->1	
tora 	a->9	b->6	d->5	e->5	f->47	g->7	h->2	i->7	k->3	m->4	n->1	o->10	p->12	r->3	s->17	t->5	u->3	v->4	å->3	
tora,	 ->2	
tora.	E->1	M->1	V->1	
tora?	A->1	
torat	 ->3	,->2	e->13	
torbr	i->14	o->1	
torcy	k->4	
torde	 ->1	
tordr	i->2	
tore 	i->1	
toren	 ->1	
torer	 ->29	,->2	.->4	n->7	
toret	 ->1	
torfö	r->2	
torga	n->1	
torha	v->1	
torhe	t->1	
toria	 ->6	,->2	.->2	
torie	l->5	n->7	r->5	t->3	
torik	 ->1	,->1	.->1	e->1	
torin	d->2	g->1	o->7	
toris	e->2	k->31	
torit	a->1	e->4	
toriu	m->10	
torka	,->1	p->1	
torkn	i->1	
torlä	r->1	
torm 	v->1	
torm,	 ->1	
torma	r->20	
torme	n->6	
tormf	ä->1	
torn 	-->2	b->1	e->2	f->3	i->2	k->1	o->5	s->3	u->1	ä->2	
torn)	.->1	
torn,	 ->12	
torn.	D->4	F->3	H->1	K->1	M->1	
torn?	A->1	
torna	 ->2	.->1	?->1	
torne	t->1	
torns	 ->4	
torpe	t->2	
torpo	l->1	
tors 	s->1	
torsa	n->1	
torsd	a->8	
torsi	n->1	
torsk	a->2	r->1	
torsl	a->2	
torsö	v->1	
tort 	a->12	b->1	e->2	f->1	g->1	h->1	i->5	k->1	m->4	n->1	p->1	s->6	t->4	u->1	
torta	m->1	
torte	r->1	
torty	r->1	
torve	n->4	
tos b	e->9	
tos e	n->1	
tos f	ö->1	
tos k	l->1	
tos o	r->1	
tos v	ä->1	
total	 ->3	a->14	b->2	f->5	i->2	s->1	t->6	v->1	
town 	a->1	ä->1	
town,	 ->1	
toxis	k->1	
tpart	 ->1	.->1	e->1	i->5	s->1	
tpeka	s->1	
tpens	i->1	
tperi	o->10	
tplan	 ->1	.->1	e->1	
tplat	t->1	
tplån	a->1	i->1	
tpoli	t->3	
tpost	 ->6	.->1	e->3	
tprat	.->1	
tpres	s->1	
tprio	r->1	
tprob	l->1	
tprog	r->1	
tproj	e->1	
tprot	o->1	
tpräg	l->1	
tpunk	t->3	
tra A	t->1	
tra E	u->3	
tra F	r->1	
tra J	e->1	
tra T	y->1	
tra a	r->1	
tra b	a->1	å->1	
tra c	e->1	
tra d	e->13	
tra f	ö->4	
tra g	e->2	ä->1	
tra h	e->1	
tra i	 ->1	n->1	
tra k	a->1	o->5	v->1	
tra l	e->1	i->1	
tra m	e->1	i->3	ä->1	
tra o	c->2	r->1	s->1	
tra p	r->1	
tra r	å->1	
tra s	i->6	o->2	t->2	y->1	ä->2	
tra t	e->1	i->1	r->1	
tra u	t->1	
tra v	ä->1	
tra ö	g->1	
tra, 	ä->1	
trad 	a->2	i->1	k->1	s->1	
trade	 ->2	
tradi	t->19	
traff	 ->2	,->1	-->2	a->4	b->1	l->1	p->2	r->28	
trafi	k->9	
trage	d->4	
tragi	s->6	
traka	s->1	
trako	p->5	
trakt	 ->2	.->1	:->1	a->24	e->1	i->1	
tral 	b->1	d->1	f->1	p->1	r->2	s->1	
tral-	 ->6	
tral.	F->1	H->1	
trala	 ->12	,->1	s->6	t->1	
tralb	a->8	
trale	r->1	u->1	
tralf	ö->1	
trali	b->1	s->25	
tralt	 ->6	,->1	
tram 	t->1	
tramn	i->2	
tramp	 ->2	
tran 	t->1	
trand	e->37	
trans	e->1	i->6	p->106	
traor	d->1	
trape	r->1	
trapp	o->1	
trapr	o->1	
trar 	a->1	d->1	e->2	f->2	h->1	k->2	m->1	o->5	r->1	s->1	t->3	v->1	
trar,	 ->3	
trar.	R->1	
trar:	 ->1	
trarn	a->6	
trars	 ->1	
tras 	a->2	d->1	f->1	m->1	o->3	
tras.	E->1	P->1	
trasa	s->1	
trasb	o->5	
trasm	a->1	
trass	l->1	
trast	e->2	
trat 	o->1	s->1	v->1	
trate	g->63	
trati	o->26	v->18	
trats	 ->2	
traum	a->1	
trava	r->1	
trave	n->1	
trax 	a->1	e->1	i->1	
tre a	l->3	n->4	t->3	
tre b	a->1	e->2	
tre d	i->1	u->1	
tre e	k->1	
tre f	j->1	r->4	u->1	ö->7	
tre g	e->1	r->3	å->2	
tre h	a->1	
tre i	 ->1	n->1	
tre k	a->1	l->1	o->7	v->1	
tre l	a->1	
tre m	e->1	i->4	o->1	y->2	å->10	ö->2	
tre o	c->5	m->5	v->1	
tre p	r->1	u->1	å->1	
tre r	e->4	ä->1	
tre s	a->3	e->3	m->1	o->1	t->4	y->1	ä->9	
tre t	i->5	j->1	
tre u	p->1	
tre v	e->3	i->3	
tre ä	n->6	
tre å	r->3	
tre ö	n->1	
tre, 	D->1	i->1	o->1	s->1	ä->1	
tre.E	n->1	
tre.I	 ->1	
tre.J	a->2	
tre.P	r->1	
tre.T	i->1	
tre: 	b->1	
trea 	o->1	
treal	 ->1	,->1	
tream	i->8	
treck	 ->1	
treda	 ->2	n->1	
tredd	 ->1	
tredj	e->72	
tredn	i->4	
trege	r->1	
tregi	o->1	
trekl	a->1	
trela	t->1	
trema	 ->2	
tremh	ö->14	
tremi	s->10	
tremt	 ->4	
tremå	n->1	
trend	 ->1	
trepr	e->3	i->2	
trera	 ->13	d->3	r->5	s->3	t->4	
treri	n->3	
tres 	l->2	v->1	
tress	a->21	e->99	
tresu	l->3	
tret 	(->1	i->1	
treta	n->1	
trett	i->2	o->3	
trevl	i->3	
tri b	e->1	
tri d	i->1	
tri i	 ->1	
tri o	c->2	
tri s	o->6	
tri, 	t->2	u->1	
tri- 	o->1	
tribu	t->1	
trich	t->6	
trici	t->1	
trid 	m->8	s->1	
trida	 ->2	
tridd	 ->2	
tride	n->1	r->7	
tridi	g->1	
tridl	i->1	
triel	l->6	
trier	 ->2	
trifr	å->4	
trike	s->19	
trikt	 ->8	.->1	a->12	i->4	
trili	k->1	
trilj	o->1	
trilo	b->1	
trin 	a->3	b->1	e->2	f->5	h->1	i->4	k->3	l->1	m->1	o->5	p->1	s->8	v->2	ä->2	
trin!	H->1	
trin,	 ->15	
trin.	 ->2	D->3	H->1	I->1	J->1	N->1	S->2	V->3	
trin:	 ->1	
trin?	P->1	
tring	 ->10	,->2	.->2	a->6	e->3	s->1	
trins	 ->9	
trio 	u->1	
triot	i->1	
tripo	l->2	
tris 	i->1	k->2	
tro a	t->4	
tro d	e->1	
tro m	å->1	
tro n	å->2	
tro p	å->2	
tro t	i->1	
tro ä	r->1	
tro.V	i->1	
troak	t->12	
trodd	e->3	
trodu	c->2	k->4	
troen	d->58	
trof 	-->1	a->1	e->2	f->5	h->2	i->3	k->1	l->1	o->2	s->4	u->1	ä->1	
trof,	 ->4	
trof.	D->2	E->1	J->1	
trofa	l->1	
trofd	r->1	
trofe	n->20	r->31	
trofh	j->1	
trofs	i->1	t->3	
troge	n->1	t->1	
trojk	a->1	
trol,	 ->1	
trol.	M->1	
trole	u->1	
troli	g->11	
troll	 ->44	!->1	,->6	-->1	.->17	:->1	a->1	e->82	f->1	m->4	o->2	s->3	u->14	v->1	
tron 	a->1	
troni	k->1	s->8	
trono	d->3	m->1	
tropa	s->2	
tror 	-->1	a->80	d->8	e->1	f->1	g->1	i->10	j->23	k->2	m->4	n->4	o->5	p->1	s->2	u->1	v->2	ä->4	
tror,	 ->1	
tros 	m->1	s->1	
trota	 ->2	
trotn	i->2	
trots	 ->46	
trott	 ->2	,->1	s->1	
troux	-->1	
trove	r->4	
trovi	c->1	
trovä	r->14	
truer	a->5	
truki	t->1	
trukt	i->30	u->153	ö->3	
trum 	f->3	i->1	m->1	å->1	
trum!	M->1	
trum,	 ->2	
trume	n->52	t->2	
trunt	a->3	p->1	
trupp	e->3	
trust	a->1	b->1	e->4	n->3	
trutt	e->1	
tryck	 ->24	,->2	.->1	a->23	b->1	e->19	l->13	n->3	s->3	t->12	
trygg	a->2	h->6	
tryk.	H->1	
tryka	 ->23	,->2	s->4	
tryke	r->2	
tryks	 ->2	
trymm	e->11	
tryps	.->1	
trä u	t->1	
trä ö	v->1	
träck	a->2	e->1	n->28	t->1	
träd 	b->1	f->1	h->1	u->1	
träd,	 ->1	
träd.	D->1	
träda	 ->10	,->1	n->10	r->57	
trädd	 ->1	a->2	e->7	
träde	 ->15	.->3	H->1	P->1	l->5	n->4	r->15	s->9	t->12	
träds	 ->2	
träff	a->115	l->2	
tränd	e->2	
träng	 ->3	a->17	d->1	e->5	n->35	t->5	
träni	n->1	
träpr	o->1	
träsk	.->1	
träto	r->1	
trätt	 ->11	a->2	e->1	
träva	 ->4	d->4	n->15	r->4	s->3	t->1	
trävi	g->1	
tråda	r->3	
tråde	n->1	
trået	.->1	
tråki	g->3	
trålk	a->1	
tråln	i->3	
tråls	k->1	
trång	 ->1	m->1	
trögh	e->1	
tröjo	r->1	
trök 	b->1	
trök,	 ->1	
tröks	,->1	
tröm 	a->2	b->1	i->1	
tröm,	 ->1	
tröm:	 ->1	
trömm	a->3	e->4	
trömn	i->6	
trösk	e->3	
tröst	 ->1	
trött	a->2	
ts "B	i->1	
ts "g	e->1	
ts (u	n->1	
ts - 	a->1	b->1	e->1	f->1	h->1	i->1	o->3	
ts 80	 ->1	
ts Ba	l->1	
ts Eu	r->1	
ts Le	i->1	
ts Sp	a->2	
ts ab	s->1	
ts al	l->15	
ts am	b->2	
ts an	d->2	g->2	s->4	t->1	
ts ar	b->4	t->2	
ts at	t->23	
ts au	k->1	
ts av	 ->68	s->1	
ts be	f->1	g->2	h->2	k->1	s->20	t->1	v->1	
ts bi	d->2	
ts bo	r->1	
ts bu	d->2	
ts bä	t->1	
ts ce	n->1	
ts co	s->1	
ts de	 ->4	l->8	m->1	n->3	r->1	t->14	
ts di	m->1	p->1	r->10	s->2	
ts do	m->2	
ts dä	r->3	
ts ef	f->2	t->1	
ts eg	e->2	
ts el	l->3	
ts en	 ->3	d->1	h->1	o->1	
ts er	f->1	
ts et	t->1	
ts ex	k->1	
ts fa	l->1	s->2	
ts fe	m->1	
ts fi	l->1	
ts fj	o->1	
ts fl	e->1	
ts fo	n->1	r->1	
ts fr	a->22	e->2	i->1	ä->1	å->4	
ts fu	l->1	n->1	
ts få	 ->3	
ts fö	r->57	
ts ge	m->11	n->6	
ts gi	l->3	
ts go	d->1	
ts gr	a->1	u->13	ä->1	
ts gå	n->1	
ts gö	r->2	
ts ha	n->1	r->1	v->1	
ts hi	s->2	t->2	
ts hj	ä->1	
ts ho	s->2	
ts hu	v->1	
ts hä	n->2	r->8	
ts hå	l->1	r->1	
ts i 	A->1	D->1	E->2	F->2	K->3	S->2	T->1	b->1	d->8	e->3	f->3	g->1	h->1	l->1	m->2	n->2	o->2	r->4	s->4	t->1	v->2	ö->1	
ts ik	r->1	
ts in	 ->2	g->1	i->2	n->2	o->3	r->2	t->3	
ts ka	n->1	
ts kl	.->2	a->1	
ts ko	m->2	n->1	r->1	
ts kr	a->2	e->1	
ts ku	s->1	
ts kä	r->1	
ts la	g->1	n->1	
ts le	d->6	g->1	
ts li	n->1	v->1	
ts lo	g->2	
ts lö	f->1	
ts ma	k->1	
ts me	d->19	l->1	n->2	r->1	
ts mi	l->2	n->2	
ts mo	n->1	t->4	
ts my	c->1	
ts må	l->2	s->1	
ts mö	j->3	t->2	
ts ne	d->3	g->1	
ts nu	 ->1	v->1	
ts ny	a->1	l->1	
ts nä	r->1	
ts nå	g->3	
ts oc	h->39	
ts oh	ö->1	
ts oi	n->1	
ts ol	i->1	
ts om	 ->6	
ts or	d->16	o->1	s->1	
ts ot	i->1	
ts pa	r->1	
ts pe	r->2	
ts pl	e->1	
ts po	l->2	r->2	
ts pr	i->4	o->2	
ts pu	b->1	n->1	
ts på	 ->18	
ts re	g->6	k->2	s->7	
ts ri	k->2	
ts rä	t->6	
ts rå	d->1	
ts sa	m->1	
ts se	d->3	s->2	
ts si	d->2	f->1	s->1	t->1	
ts sk	r->1	u->2	
ts sl	u->5	
ts so	l->1	m->6	
ts sp	ö->1	
ts st	r->4	ä->2	å->7	ö->2	
ts su	v->2	
ts sv	å->1	
ts sy	n->4	
ts sä	r->1	
ts så	 ->1	
ts ta	l->3	
ts te	x->1	
ts ti	d->1	l->36	o->1	
ts tj	ä->1	
ts tr	o->3	
ts un	d->9	
ts up	p->20	
ts ut	 ->4	.->4	a->1	f->1	i->1	s->3	t->1	v->1	
ts va	d->2	p->1	r->2	
ts ve	r->2	t->1	
ts vi	d->5	s->1	
ts vä	g->1	r->1	
ts yt	t->3	
ts än	d->2	n->3	
ts är	 ->4	
ts ål	d->1	
ts ås	i->1	
ts åt	 ->2	e->1	
ts ön	s->1	
ts öv	e->2	r->1	
ts!Fö	r->1	
ts, S	t->1	
ts, a	l->1	t->2	
ts, b	e->2	
ts, d	ä->2	
ts, e	f->1	l->1	n->1	t->1	
ts, f	ö->1	
ts, h	a->1	
ts, i	 ->1	n->2	
ts, m	e->4	å->1	
ts, n	ä->3	å->1	
ts, o	c->5	
ts, p	å->1	
ts, s	o->1	å->3	
ts, t	r->2	
ts, u	n->1	p->1	
ts, v	a->1	i->3	å->1	
ts, ä	r->1	
ts, å	t->2	
ts- o	c->12	
ts-be	l->1	
ts.An	h->1	
ts.Be	t->1	
ts.De	 ->1	n->4	t->11	
ts.Dä	r->2	
ts.Då	 ->2	
ts.Ef	t->1	
ts.En	 ->2	d->1	l->1	
ts.Er	t->1	
ts.Fa	c->1	
ts.He	r->1	
ts.Ho	p->1	
ts.I 	d->1	
ts.Ja	g->5	
ts.Ko	m->1	n->1	s->1	
ts.Me	n->1	
ts.Mi	n->1	
ts.Nä	r->1	
ts.Ra	p->1	
ts.Re	a->1	
ts.Sl	u->2	
ts.So	m->1	
ts.Så	 ->1	
ts.Ta	c->1	
ts.Vi	 ->2	l->1	
ts.Än	n->1	
ts: v	a->1	
ts?Fr	å->1	
ts?Ko	m->1	
tsa a	l->1	
tsa m	e->1	
tsa p	å->4	
tsa s	ä->1	
tsakt	 ->2	.->1	e->2	
tsam 	b->1	t->1	v->1	
tsam,	 ->1	
tsamh	e->6	
tsamm	a->9	
tsamt	 ->5	.->1	
tsana	l->3	
tsand	a->4	e->1	
tsanl	ä->4	
tsar 	i->1	k->1	n->1	p->2	r->1	
tsar.	S->1	
tsarb	e->1	
tsarg	u->1	
tsas 	k->1	m->1	o->1	s->1	
tsasp	e->3	
tsat 	n->1	
tsats	 ->15	e->43	f->1	
tsatt	 ->11	,->1	a->14	s->1	
tsavb	r->1	
tsavt	a->1	
tsban	k->2	
tsbas	.->1	e->1	
tsbeh	a->2	
tsbek	ä->3	
tsbes	k->1	l->4	t->1	
tsbet	ä->1	
tsbud	g->1	
tsbör	d->5	
tscen	t->1	
tscer	t->1	
tsche	 ->1	f->3	
tsdeb	a->1	
tsdok	u->4	
tse d	e->1	
tse e	n->2	
tse f	r->4	
tse m	y->1	
tse o	c->1	m->1	
tse v	i->1	
tse.E	n->1	
tseda	n->3	
tsedd	a->1	
tseen	d->1	
tsekt	o->2	
tsel 	o->4	
tsel.	D->1	
tsen 	E->1	a->7	b->4	h->1	m->4	t->1	v->2	ä->2	
tsen!	N->1	
tsen,	 ->1	
tsen.	 ->1	J->1	K->1	
tsen;	 ->1	
tsenh	e->3	
tser 	-->1	a->2	b->2	f->12	i->5	k->1	m->2	o->3	p->3	s->8	u->1	v->3	å->1	ö->2	
tser,	 ->7	
tser.	-->1	D->2	E->1	F->1	J->2	K->1	
tsern	a->20	
tses 	d->1	f->1	
tses.	A->1	
tsett	 ->3	s->1	
tsfat	t->11	
tsfie	n->1	
tsfla	g->15	
tsfor	d->1	m->1	u->1	
tsfrå	g->10	
tsfån	g->1	
tsför	d->4	e->1	f->1	h->1	k->2	l->2	o->1	
tsgar	a->3	
tsgiv	a->8	
tsgre	n->2	
tsgru	p->5	
tsgrä	n->1	
tshan	d->2	
tshjä	l->2	
tsiff	r->2	
tsiga	 ->1	
tsikt	e->1	i->4	
tsins	a->2	p->1	t->2	
tsitu	a->2	
tska 	e->1	
tskaf	f->1	
tskal	:->1	
tskam	p->1	
tskan	 ->1	
tskap	e->1	i->1	
tskil	l->3	
tskip	n->7	
tskla	u->1	
tskli	m->1	
tskoe	f->1	
tskol	l->1	
tskon	c->1	t->1	
tskot	t->163	
tskra	f->4	v->1	
tskri	d->1	s->2	t->1	
tskul	t->1	
tskyd	d->8	
tslag	 ->2	,->1	.->1	e->1	i->1	n->12	s->2	
tsled	a->28	
tslig	 ->17	a->75	h->13	t->29	
tslin	g->2	
tsliv	e->2	
tslog	 ->1	s->1	
tslop	p->2	
tsläg	e->3	
tsläm	n->2	
tslän	d->1	
tsläp	p->9	
tslå 	E->1	a->1	k->1	n->1	v->1	
tslår	 ->4	
tslås	 ->7	.->1	
tslös	a->6	h->37	
tsmak	t->2	
tsman	n->1	
tsmar	k->12	
tsmed	e->1	
tsmet	o->3	
tsmin	i->2	
tsmyn	d->10	
tsmän	g->1	n->1	
tsmål	 ->1	s->1	
tsnin	g->4	
tsniv	å->6	
tsnor	m->6	
tsnät	e->1	
tsoff	e->2	
tsoly	c->1	
tsomr	å->5	ö->1	
tsord	n->13	
tsorg	a->3	
tsos 	o->2	
tsos,	 ->1	
tsosä	k->2	
tspak	t->4	
tspar	k->1	
tsper	i->1	s->1	
tspla	n->7	t->4	
tspol	i->7	
tspra	x->1	
tspri	n->72	o->1	
tspro	b->2	c->5	d->1	g->4	t->1	
tspår	 ->1	,->1	
tsram	e->1	
tsrap	p->2	
tsrea	k->1	
tsreg	e->3	i->1	l->1	
tsris	k->1	
tsrub	r->1	
tsrum	 ->1	
tsrut	i->1	
tsrät	t->4	
tsråd	 ->1	.->1	e->2	g->14	
tssan	k->1	
tssek	r->1	t->4	
tssif	f->2	
tsski	p->3	
tsskä	l->2	
tsspr	å->1	
tssta	d->1	t->9	
tssty	r->5	
tsstö	d->19	
tssyn	e->1	
tssys	t->22	
tssäk	e->21	
tstag	a->40	
tstak	,->1	
tstat	i->10	u->1	
tstid	 ->2	,->1	e->4	s->3	
tstil	l->40	
tstjä	n->1	
tstra	d->1	m->2	
tstru	k->1	
tsträ	c->28	v->2	
tstyc	k->3	
tstäl	l->53	
tstän	k->2	
tstån	d->10	
tstår	 ->2	
tståt	t->1	
tstöd	 ->1	e->1	
tstöt	t->1	
tsuga	r->1	
tsutb	i->2	y->3	
tsuts	k->2	
tsvag	 ->1	
tsvan	s->1	
tsvar	a->15	i->2	
tsven	t->1	
tsver	k->1	
tsvil	j->1	l->4	
tsväs	e->4	
tsynp	u->1	
tsyst	e->1	
tsäga	 ->1	n->1	
tsäge	l->8	
tsäke	r->8	
tsätt	 ->1	a->46	e->42	n->56	s->7	
tså E	u->1	
tså a	n->1	t->3	v->1	
tså b	i->1	r->1	
tså d	e->2	
tså e	n->3	t->1	
tså f	r->2	å->1	ö->2	
tså g	e->1	
tså i	 ->1	n->10	
tså k	o->1	
tså l	ä->1	
tså m	y->1	å->1	
tså p	o->1	å->1	
tså r	e->2	ä->1	
tså s	a->1	e->2	i->1	j->1	t->3	ä->1	å->2	
tså t	a->2	i->3	
tså v	a->3	e->1	i->1	
tså, 	f->1	h->1	
tsågs	 ->1	.->2	
tsåtg	ä->2	
tt "P	o->1	
tt "o	b->1	
tt (5	7->1	
tt (9	6->1	
tt - 	d->1	g->1	i->1	k->1	n->1	o->1	s->1	v->2	å->1	ö->1	
tt 19	9->3	
tt 23	,->1	
tt 25	 ->1	
tt 40	 ->1	
tt 50	-->1	
tt 70	 ->1	
tt 8 	r->1	
tt 80	 ->1	
tt 98	 ->1	
tt Al	t->1	
tt Am	s->3	
tt Ba	r->3	
tt Be	r->1	
tt Bo	u->1	
tt Br	y->1	
tt CE	N->1	
tt Da	n->3	
tt EG	-->8	:->2	
tt EI	F->1	
tt EK	S->1	
tt EL	D->1	
tt EU	 ->5	-->1	.->1	:->6	
tt Er	i->1	
tt Eu	r->79	
tt Ev	a->1	
tt FE	O->1	
tt FN	-->1	:->1	
tt FP	Ö->1	
tt Fl	o->2	
tt Fö	r->1	
tt Gr	e->1	
tt Ha	i->1	
tt IC	E->1	
tt IN	T->1	
tt Ir	l->1	
tt Is	r->3	
tt It	a->1	
tt Jö	r->3	
tt Ko	u->2	
tt Ky	o->1	
tt Ma	l->1	r->1	
tt Na	t->1	
tt OL	A->3	
tt Pa	t->1	
tt Po	r->2	
tt RI	N->1	
tt Ra	n->1	
tt Ro	t->1	
tt Sa	n->1	
tt So	k->1	
tt St	o->1	
tt Th	e->2	
tt To	t->1	
tt Tu	r->13	
tt Vä	r->1	
tt ab	s->1	
tt ac	c->5	
tt ad	 ->1	d->1	e->2	
tt ag	e->14	
tt ak	t->7	
tt al	d->2	l->51	t->2	
tt am	b->1	e->2	
tt an	a->7	d->6	f->4	g->4	m->1	n->18	o->2	p->2	s->40	t->41	v->20	
tt ar	b->53	g->1	r->1	t->3	
tt as	y->1	
tt at	t->72	
tt av	 ->26	a->1	f->2	g->8	h->1	l->2	s->24	t->10	v->4	
tt ba	l->1	n->1	r->5	
tt be	 ->2	a->8	d->5	f->7	g->19	h->18	k->29	l->3	m->4	n->1	r->6	s->44	t->42	v->29	
tt bi	b->3	d->16	f->1	l->13	n->2	o->1	s->1	
tt bl	.->1	a->3	i->43	u->1	y->1	
tt bo	 ->1	g->1	m->1	r->2	s->2	t->1	
tt br	a->20	e->8	i->4	o->7	y->7	ä->2	å->1	
tt bu	d->3	
tt by	g->15	r->1	
tt bä	r->1	t->11	
tt bå	d->4	
tt bö	r->24	
tt ce	n->3	
tt ci	t->1	v->1	
tt da	g->7	t->2	
tt de	 ->171	,->1	b->7	c->1	f->1	l->15	m->9	n->207	r->4	s->41	t->545	
tt di	a->1	l->2	p->1	r->25	s->29	v->1	
tt dj	u->2	ä->2	
tt do	k->5	m->9	
tt dr	a->14	i->9	å->1	ö->1	
tt du	b->2	
tt dy	k->1	n->1	
tt dä	m->2	r->6	
tt då	l->1	
tt dö	 ->1	d->1	l->2	m->6	
tt e-	m->1	
tt ef	f->17	t->9	
tt eg	e->14	
tt ek	o->5	
tt el	-->1	i->1	l->6	
tt em	b->1	
tt en	 ->91	a->2	b->3	d->7	e->2	g->1	h->13	k->1	l->2	o->4	s->1	
tt ep	o->1	
tt er	a->1	b->2	f->2	h->1	i->2	k->5	s->3	t->4	
tt et	a->4	t->33	
tt eu	r->11	
tt ev	e->3	
tt ex	a->1	c->1	e->19	i->1	p->3	t->1	
tt fa	k->4	l->4	n->2	r->4	s->13	t->6	
tt fe	d->1	l->2	m->2	
tt fi	n->18	s->1	
tt fl	e->14	y->5	
tt fo	d->1	k->1	l->6	n->1	r->31	t->1	
tt fr	a->22	e->7	i->3	u->1	y->1	ä->28	å->17	
tt fu	l->12	n->11	
tt fy	l->1	r->1	
tt få	 ->88	.->1	t->1	
tt fö	l->8	r->333	
tt ga	m->1	n->2	r->19	
tt ge	 ->51	.->1	m->28	n->55	
tt gi	v->2	
tt gl	o->1	ä->1	
tt go	d->17	t->9	
tt gr	a->14	e->1	i->4	u->5	
tt gy	n->4	
tt gä	l->5	
tt gå	 ->24	.->1	
tt gö	r->107	
tt ha	 ->43	,->1	d->1	l->3	m->1	n->52	r->2	
tt he	d->1	l->7	m->5	n->1	
tt hi	n->4	s->3	t->4	
tt hj	ä->17	
tt ho	n->7	p->2	s->2	t->2	
tt hu	g->3	m->1	n->1	r->3	s->1	v->3	
tt hy	c->1	s->1	
tt hä	n->8	r->2	v->2	
tt hå	l->25	n->1	r->2	
tt hö	g->6	j->2	r->11	
tt i 	2->1	A->1	C->1	E->1	L->1	a->8	b->1	d->14	e->4	f->5	g->4	j->1	k->4	m->4	o->4	p->3	s->6	t->2	v->3	Ö->1	ä->1	
tt i.	D->1	
tt ia	k->1	
tt ib	l->3	
tt ic	k->1	
tt id	e->4	é->2	
tt if	r->6	
tt ig	e->3	å->1	
tt im	m->2	p->1	
tt in	 ->5	b->1	c->1	d->1	f->29	g->21	h->1	i->10	l->14	n->12	o->6	r->21	s->28	t->49	v->3	
tt ir	l->2	o->1	r->2	
tt is	o->2	
tt it	a->1	
tt ja	 ->1	g->84	p->1	
tt jo	b->1	r->3	
tt ju	 ->1	n->1	r->2	s->3	
tt jä	m->4	
tt ka	m->4	n->14	p->3	t->1	
tt kl	a->17	o->2	y->1	
tt kn	u->1	y->2	ä->1	
tt ko	l->6	m->166	n->47	p->1	r->12	s->9	
tt kr	a->9	i->7	ä->16	
tt ku	l->9	n->51	s->1	
tt kv	a->4	i->3	ä->2	
tt kä	n->1	r->5	
tt kö	l->3	p->1	
tt la	g->9	n->35	p->3	s->1	
tt le	d->16	g->3	v->7	
tt li	d->1	g->3	k->3	l->1	n->3	s->1	t->3	v->8	
tt lj	u->1	
tt lo	c->1	g->1	k->1	
tt lu	d->2	g->2	t->1	
tt ly	c->8	f->2	s->5	
tt lä	g->43	m->10	n->1	r->3	t->2	
tt lå	g->1	n->1	t->12	
tt lö	p->2	s->19	
tt ma	j->4	n->205	r->15	s->1	t->2	x->2	
tt me	d->62	k->1	l->2	r->11	t->1	
tt mi	g->4	l->11	n->36	r->1	s->6	t->1	x->1	
tt mo	b->2	d->4	g->1	n->1	r->1	t->16	
tt mu	l->2	s->1	
tt my	c->45	n->12	
tt mä	n->8	r->2	t->1	
tt må	l->16	n->5	s->3	
tt mö	j->5	r->1	t->6	
tt na	r->1	t->4	z->1	
tt ne	d->1	g->2	k->1	
tt ni	 ->42	,->2	v->3	
tt no	g->2	m->1	r->3	
tt nu	 ->2	m->1	
tt ny	a->2	d->1	k->2	l->1	n->1	t->23	
tt nä	m->1	r->17	s->5	t->1	
tt nå	 ->10	g->19	
tt nö	d->1	j->2	t->1	
tt oa	c->1	
tt ob	e->3	
tt oc	h->38	k->15	
tt od	j->1	
tt oe	f->1	r->1	
tt of	f->7	t->1	ö->2	
tt og	r->1	
tt ok	r->1	u->1	
tt ol	j->4	y->2	ä->1	
tt om	 ->30	b->2	e->4	f->11	h->1	k->1	o->1	p->1	r->26	s->4	v->2	
tt on	ö->2	
tt op	a->1	e->1	p->1	r->1	
tt or	d->12	g->7	o->5	s->1	ä->1	
tt os	s->5	v->1	
tt ot	i->1	
tt oä	n->1	
tt oö	v->1	
tt pa	l->1	p->1	r->64	s->3	
tt pe	a->1	k->1	n->5	r->12	s->1	
tt pi	l->1	
tt pl	a->8	
tt po	l->15	p->1	s->9	ä->3	
tt pr	a->4	e->8	i->10	o->45	ö->2	
tt pu	n->1	
tt på	 ->43	.->1	b->1	g->1	m->3	p->5	s->6	t->1	v->8	
tt ra	d->1	m->2	n->1	p->2	s->1	t->1	
tt re	a->3	d->3	f->14	g->30	l->1	n->4	p->4	s->26	t->3	v->4	
tt ri	d->1	k->18	m->2	n->1	s->1	
tt ro	 ->1	p->1	
tt ru	m->1	t->1	
tt ry	k->1	
tt rä	c->1	d->5	k->1	t->14	
tt rå	d->25	
tt rö	r->1	s->31	t->1	
tt s.	k->1	
tt sa	g->1	k->3	l->1	m->49	n->1	t->2	
tt se	 ->50	d->2	g->3	k->2	m->2	n->3	r->5	x->1	
tt si	f->1	g->8	n->2	s->2	t->4	
tt sj	u->2	ä->10	
tt sk	a->79	e->6	i->8	j->5	o->1	r->5	u->3	y->27	ä->4	ö->2	
tt sl	a->3	i->1	u->12	ä->3	å->4	ö->1	
tt sm	å->1	
tt sn	a->7	
tt so	c->8	l->3	m->46	r->1	
tt sp	a->2	e->11	r->2	å->2	ö->1	
tt st	a->23	e->13	i->3	o->24	r->12	u->1	y->6	ä->19	å->9	ö->66	
tt su	b->1	c->1	d->1	
tt sv	a->13	e->1	
tt sy	f->2	m->1	n->2	r->1	s->25	
tt sä	g->26	k->22	l->1	n->4	r->6	t->32	
tt så	 ->20	d->40	v->3	
tt sö	k->1	r->2	
tt t.	o->1	
tt ta	 ->84	.->1	?->1	c->17	g->2	k->1	l->10	n->1	p->1	s->4	
tt te	c->2	m->1	r->1	
tt th	e->1	
tt ti	d->13	l->135	t->4	
tt tj	ä->3	
tt to	l->5	r->1	t->3	
tt tr	a->5	e->3	o->2	u->1	y->1	ä->5	
tt tu	n->1	r->1	s->1	
tt tv	e->2	i->4	å->2	
tt ty	c->3	d->11	
tt tä	c->1	n->10	p->2	
tt tå	g->2	
tt ul	t->1	
tt un	d->65	i->10	
tt up	p->83	
tt ur	 ->5	h->1	s->1	v->3	
tt ut	 ->1	a->18	b->1	e->5	f->13	g->2	i->2	j->3	k->1	l->1	m->11	n->12	o->1	p->1	r->3	s->5	t->30	v->46	ö->8	
tt va	c->2	d->4	k->2	l->2	r->66	
tt ve	d->2	r->22	t->4	
tt vi	 ->381	,->6	d->36	k->17	l->12	n->4	s->26	t->1	
tt vr	a->1	
tt vä	c->2	g->3	l->15	n->10	r->3	s->1	x->4	
tt vå	l->1	r->21	
tt wo	r->1	
tt yp	p->1	
tt yt	t->18	
tt zo	n->1	
tt äg	a->17	n->4	
tt äm	b->2	
tt än	 ->3	d->34	n->1	
tt är	 ->18	,->1	e->3	
tt äv	e->20	
tt å 	e->3	
tt åk	l->1	
tt ål	d->1	
tt år	 ->17	,->1	.->2	h->1	s->1	
tt ås	i->1	t->5	
tt åt	 ->1	a->4	e->36	f->2	g->5	m->2	
tt öd	e->1	
tt ög	o->1	
tt ök	a->22	
tt öm	s->1	
tt ön	s->3	
tt öp	p->9	
tt ös	t->1	
tt öv	e->53	
tt, E	G->1	
tt, a	t->3	
tt, b	e->1	l->1	
tt, d	e->1	i->1	
tt, e	f->3	l->2	n->2	
tt, f	a->1	r->3	å->1	ö->4	
tt, g	i->1	ä->1	ö->1	
tt, h	a->2	e->1	ä->1	
tt, i	 ->4	
tt, k	a->2	r->1	u->1	
tt, l	i->1	
tt, m	e->4	
tt, n	ä->1	
tt, o	c->9	m->2	
tt, p	å->1	
tt, r	e->1	
tt, s	i->1	k->1	o->3	å->4	
tt, t	a->1	i->2	r->2	v->3	
tt, u	r->1	t->1	
tt, v	i->4	
tt, ä	v->3	
tt, å	r->1	
tt. D	e->2	
tt. I	n->1	
tt..(	D->1	
tt...	(->1	
tt.Al	l->2	
tt.Be	t->1	
tt.De	 ->2	n->5	s->1	t->20	
tt.Dä	r->2	
tt.En	 ->2	
tt.Er	f->1	
tt.Fö	r->7	
tt.He	r->9	
tt.I 	a->1	f->1	u->1	v->1	
tt.Ja	g->13	
tt.Ko	m->3	
tt.Lå	t->4	
tt.Ma	n->1	
tt.Me	n->7	
tt.Mi	l->1	n->1	
tt.Mo	r->1	t->1	
tt.Na	t->1	
tt.Ni	 ->1	
tt.Nä	r->1	
tt.Ob	e->1	
tt.Om	 ->1	
tt.Or	o->1	
tt.PP	E->1	
tt.Pa	r->3	
tt.Sl	u->1	
tt.So	m->1	
tt.St	a->1	
tt.Sy	f->1	
tt.Ta	c->1	
tt.Ut	f->1	
tt.Vi	 ->5	d->1	s->1	
tt.Äv	e->3	
tt: "	D->2	
tt: H	o->1	
tt: j	a->1	
tt: o	m->1	
tt: s	y->1	
tt?An	s->1	
tt?De	t->1	
tt?Om	 ->1	
tt?Sk	u->1	
tt?Vi	l->1	
ttBet	ä->1	
tta -	 ->5	,->1	
tta A	l->1	
tta E	G->5	U->1	u->2	
tta F	P->1	
tta a	b->1	l->2	n->7	r->5	t->22	v->18	
tta b	a->2	e->63	i->2	l->3	o->1	u->1	ä->1	ö->4	
tta c	e->2	
tta d	a->1	e->31	i->33	j->1	o->6	r->2	ä->1	
tta e	f->2	k->2	l->1	n->27	r->2	t->19	v->1	x->1	
tta f	a->16	i->2	l->2	o->3	r->5	å->5	ö->60	
tta g	e->3	i->1	l->1	o->2	r->4	ä->3	
tta h	a->22	e->1	i->1	o->1	u->1	ä->5	å->1	
tta i	 ->21	n->37	
tta k	a->16	o->15	r->5	v->1	ä->2	
tta l	a->5	e->2	i->6	j->1	ä->1	
tta m	a->4	e->33	i->7	o->2	y->6	ä->2	å->20	ö->2	
tta n	a->3	o->2	u->1	y->2	ä->4	å->2	
tta o	a->1	b->1	c->20	e->1	l->1	m->43	n->1	r->6	s->2	
tta p	a->40	l->2	o->2	r->31	u->1	å->23	
tta r	e->9	i->1	u->1	ä->1	å->2	
tta s	a->31	e->5	i->10	j->1	k->27	l->9	m->1	o->13	p->6	t->21	y->8	ä->10	å->3	
tta t	a->4	e->2	i->12	o->2	r->1	v->2	y->2	å->1	
tta u	n->3	p->4	r->2	t->17	
tta v	a->13	e->1	i->16	o->1	å->3	
tta y	t->2	
tta ä	m->2	n->6	r->149	v->3	
tta å	r->3	s->1	t->5	
tta ö	k->3	v->3	
tta!D	e->1	
tta!F	r->1	
tta, 	a->2	b->1	d->1	e->1	f->7	h->5	i->2	k->2	m->8	o->11	s->1	t->3	u->1	v->2	
tta. 	F->1	
tta.(	P->1	
tta..	(->1	
tta.A	n->1	
tta.B	e->2	
tta.C	o->1	
tta.D	e->19	å->1	
tta.E	f->3	n->2	
tta.F	r->1	ö->1	
tta.G	e->1	
tta.H	e->3	
tta.I	 ->5	n->1	
tta.J	a->8	
tta.K	o->1	
tta.M	e->6	
tta.N	u->1	ä->1	
tta.O	c->1	m->2	
tta.P	r->2	å->1	
tta.S	e->1	o->1	t->2	å->1	
tta.T	o->1	
tta.V	a->3	i->7	å->1	
tta.Ä	r->1	
tta: 	J->1	
tta?J	a->1	
ttack	 ->2	e->1	
ttad 	f->1	ö->1	
ttade	 ->16	,->1	.->2	s->3	
ttag.	V->1	
ttaga	n->7	r->4	
ttage	l->1	
ttagi	t->3	
ttagn	i->2	
ttala	 ->21	d->13	n->51	r->8	s->1	t->4	
ttan 	o->2	
ttan.	D->1	
ttand	e->66	
ttant	,->1	
ttar 	E->1	F->1	a->6	b->5	d->12	e->6	f->2	i->2	j->3	k->2	n->1	o->1	p->5	r->1	s->4	t->3	u->3	v->3	ä->1	
ttar.	Ä->1	
ttare	 ->13	,->2	.->1	n->2	
ttarh	u->1	
ttarn	a->5	
ttas 	a->15	b->2	d->3	e->7	f->2	g->1	i->10	m->3	p->3	s->1	u->1	v->2	ä->1	
ttas,	 ->4	
ttas.	 ->1	J->1	P->1	V->1	
ttat 	a->1	e->5	f->3	h->1	l->1	m->2	o->1	s->3	u->1	v->2	
ttat.	E->1	
ttats	 ->12	,->1	.->1	
ttavl	a->7	
tte O	u->1	
tte d	e->2	
tte i	 ->2	
tte j	ä->1	
tte m	å->1	
tte o	c->1	m->1	
tte p	e->10	
tte r	a->2	e->4	
tte ö	v->2	
tte, 	m->1	
tte- 	o->1	
tte-L	e->1	
tteba	s->1	
ttebe	s->2	t->12	
ttede	l->1	
ttefr	i->1	å->1	
ttefö	r->1	
ttegå	n->1	
ttein	c->1	s->1	
tteli	g->1	
ttels	e->3	
ttelä	t->1	
tten 	-->1	I->1	a->28	b->1	e->2	f->5	g->4	h->7	i->6	k->2	m->7	n->3	o->25	p->3	s->8	t->7	u->5	v->5	ä->3	ö->1	
tten!	 ->2	
tten)	 ->1	
tten,	 ->27	
tten.	"->1	A->1	D->5	E->2	F->3	H->3	I->1	J->4	K->1	M->3	N->1	O->2	R->1	S->4	T->2	V->3	
tten;	 ->2	
tten?	K->1	
ttenF	r->1	
ttenH	e->1	
ttend	e->1	r->1	
ttenf	ö->2	
ttenl	ö->1	
ttenp	r->1	
ttenr	e->2	
ttens	 ->10	
ttent	a->5	
ttenv	ä->8	
ttepo	l->1	
tter 	a->14	d->11	e->7	g->2	h->1	i->4	j->1	k->3	l->2	m->6	n->1	o->13	p->1	r->1	s->10	t->2	u->1	v->4	Ö->1	ä->3	
tter,	 ->3	
tter.	D->1	J->1	
ttera	 ->11	n->6	r->1	s->6	t->11	
tterd	a->2	ö->1	
tteri	 ->1	e->2	n->5	
tterl	i->55	
ttern	a->4	
ttero	m->1	
tterr	a->2	
tters	k->1	t->33	
tterv	ä->1	
ttes 	3->1	a->1	i->3	u->1	
ttes.	O->1	V->1	
ttesa	t->1	
ttesy	s->1	
ttet 	,->1	-->1	a->11	d->4	e->2	f->85	g->2	h->5	i->4	k->4	l->1	n->1	o->6	p->1	s->2	u->1	v->1	ä->3	
ttet,	 ->9	
ttet.	D->2	H->1	I->2	J->3	M->1	V->2	
ttet:	 ->1	
ttets	 ->7	
ttfra	m->1	
ttful	l->1	
ttfär	d->7	
ttför	s->1	
ttgör	a->1	
tthål	l->9	
tti g	j->1	
ttich	e->1	
ttide	n->1	
ttig 	f->2	o->1	r->1	u->1	å->1	ö->1	
ttiga	 ->16	,->2	d->9	n->1	r->3	s->4	t->8	
ttigd	o->12	
ttigh	e->103	
ttigt	 ->3	,->1	
ttill	g->2	s->44	v->1	
ttin,	 ->1	
ttinn	e->1	
ttiof	e->1	
ttiot	a->1	
ttisk	 ->1	-->1	a->12	t->2	
ttit 	a->1	
ttity	d->5	
ttja 	a->5	c->1	d->5	i->1	o->1	s->5	
ttjad	e->4	
ttjan	d->9	
ttjar	 ->3	
ttjas	 ->6	
ttjat	 ->1	
ttjän	t->25	
ttkri	g->1	
ttkvä	l->1	
ttlan	d->5	
ttle 	o->2	ä->1	
ttle.	V->1	
ttlig	a->1	t->1	
ttmät	i->1	
ttmål	s->1	
ttna 	d->1	e->1	p->1	
ttna.	 ->1	
ttnad	e->1	
ttnar	 ->7	
ttnas	 ->2	.->1	
ttne 	o->1	t->1	
ttnen	 ->1	,->1	.->1	
ttnet	 ->4	.->2	
ttnin	g->287	
tto a	c->1	
tto f	ö->1	
tto-a	n->1	
ttoan	a->1	
ttolk	a->1	
tton 	m->1	o->1	v->1	å->1	
ttona	t->1	
ttond	e->2	
ttone	r->1	
ttons	 ->1	
ttor 	o->1	
ttork	n->1	
ttorn	a->1	
ttra 	E->1	a->1	b->2	d->13	f->2	g->3	i->1	k->5	l->2	m->4	o->2	s->9	t->2	
ttrad	 ->4	e->2	
ttraf	i->1	
ttrak	t->1	
ttran	d->33	
ttrar	 ->6	
ttras	 ->5	.->2	
ttrat	 ->2	s->2	
ttre 	a->6	b->2	d->1	e->1	f->6	g->3	h->1	i->1	k->6	l->1	m->5	o->5	r->4	s->14	t->5	u->1	v->1	ä->6	
ttre,	 ->3	
ttre.	E->1	I->1	J->2	P->1	T->1	
ttret	a->1	
ttrin	g->21	
ttryc	k->72	
tträd	a->5	
tts a	l->1	n->1	t->1	v->5	
tts b	e->1	
tts f	r->1	ö->8	
tts g	e->1	
tts h	ä->1	
tts i	 ->4	
tts k	o->1	
tts m	e->1	o->1	
tts n	u->1	
tts o	c->1	
tts p	å->1	
tts u	n->2	p->1	t->2	
tts v	a->1	
tts ö	v->1	
tts, 	m->1	n->1	t->1	
tts- 	o->1	
tts.D	e->3	
tts.E	n->1	
tts.I	 ->1	
tts.N	ä->1	
tts.R	a->1	
ttsak	t->4	
ttsbe	h->2	k->3	t->1	
ttsde	b->1	
ttsfr	å->1	
ttsfö	r->1	
ttshj	ä->2	
ttsin	s->2	
ttska	f->1	
ttski	p->7	
ttsku	l->1	
ttsli	g->130	n->2	
ttslä	g->3	
ttsmy	n->1	
ttsmå	l->1	
ttsof	f->2	
ttsom	r->1	
ttsor	d->3	
ttsos	ä->2	
ttspa	r->1	
ttspr	a->1	i->1	o->1	
ttsre	g->2	
ttsru	b->1	
ttsse	k->1	
ttssk	i->3	
ttsst	a->9	
ttssy	s->20	
ttssä	k->20	
ttsti	l->2	
ttstj	ä->1	
ttstr	a->1	
ttsvä	s->4	
ttvik	t->2	
ttvil	l->1	
ttvis	 ->6	.->1	a->50	o->3	t->12	
ttysk	l->2	
ttänk	a->1	
tté -	 ->2	
tté e	l->1	
tté f	ö->3	
tté h	a->1	
tté m	e->1	
tté s	o->2	
ttéer	.->1	n->3	
ttéfö	r->2	
ttén 	(->2	f->3	i->1	k->1	l->1	o->11	s->2	v->1	ä->1	
ttén,	 ->4	
ttén.	H->1	M->1	
ttén?	V->1	
tténs	 ->11	
ttésy	s->2	
ttömd	,->1	
ttömm	a->3	
ttömt	 ->1	
tu me	d->20	n->1	
tuali	s->1	
tuati	o->129	
tud 7	 ->1	
tuden	t->2	
tuder	a->3	
tudie	 ->1	b->1	p->1	r->6	
tuell	 ->7	.->3	a->31	t->14	
tuera	 ->2	r->1	
tuff 	n->1	
tuffa	r->1	
tugal	 ->15	,->4	s->7	
tugis	i->70	
tugor	,->1	
tugue	s->1	
tulat	i->6	
tuler	a->33	
tulla	r->2	
tullf	ö->1	
tullg	å->1	
tum a	t->56	
tum d	å->1	
tum f	ö->3	
tum i	n->1	
tum m	å->1	
tum o	c->3	
tum s	k->1	o->4	
tum ä	r->4	
tum å	s->1	
tum, 	b->1	m->1	o->1	
tum.D	e->1	
tum.I	 ->1	
tum.V	i->2	
tumet	 ->2	.->1	
tumma	 ->3	
tunc 	d->1	
tund 	(->2	s->6	
tunda	n->2	
tunde	n->6	r->1	
tung 	a->1	b->1	o->1	p->2	u->1	
tunga	 ->1	,->1	n->1	
tungm	e->6	
tungr	o->1	
tungt	 ->1	,->1	
tunis	m->1	t->1	
tunne	l->3	
tunnl	a->2	
tur -	 ->2	
tur 2	0->20	
tur b	a->1	e->2	
tur d	e->1	r->1	ä->1	
tur e	t->1	
tur f	o->1	ö->6	
tur g	e->1	
tur h	o->1	
tur i	 ->2	n->2	
tur k	a->1	
tur o	c->7	
tur p	å->1	
tur s	k->1	o->7	
tur u	n->1	t->1	
tur v	e->1	i->1	
tur ä	r->4	
tur, 	(->1	G->1	a->2	h->1	l->1	m->3	o->3	s->1	t->2	u->3	å->1	
tur- 	o->2	
tur.D	e->3	
tur.F	o->1	
tur.N	i->1	
tur.O	m->1	
tur.T	y->1	
tur.V	i->3	
tur?M	e->1	
tura.	D->1	
turak	t->1	
turan	s->1	
turar	b->1	v->5	
turbe	s->1	
turel	l->40	
turen	 ->37	,->5	.->4	?->1	s->7	
turer	 ->12	,->4	.->4	a->6	i->9	n->6	s->1	
turfo	n->58	r->1	
turfö	r->2	
turhi	s->1	
turie	n->1	
turis	m->20	t->4	
turk-	d->1	
turka	r->2	t->13	
turki	s->6	
turli	g->102	
turmä	s->1	
turnä	t->1	
turnö	d->1	
turom	r->2	
turpo	l->16	
turpr	o->4	
turre	f->1	
turse	k->5	
turst	ö->3	
turut	g->1	s->1	v->1	
turve	t->1	
turåt	g->1	
tus a	v->1	
tus e	n->1	
tus q	u->2	
tus.D	e->1	
tus?O	c->1	
tusen	 ->3	,->1	d->3	t->10	
tusfö	r->1	
tusia	s->3	
tutio	n->158	
tutsk	o->12	
tutvi	d->2	
tvakt	e->1	
tvald	 ->1	
tvape	n->1	
tvara	n->2	
tvaro	r->1	
tveck	l->238	
tveka	 ->2	d->1	n->15	r->3	t->2	
tvekl	ö->1	
tveks	a->5	
tverk	 ->11	,->1	.->2	?->1	a->8	e->6	
tvers	i->1	
tvety	d->7	
tvidg	a->36	n->71	
tvikt	 ->1	n->3	s->2	
tvill	i->2	
tvin 	o->1	
tving	a->32	
tvis 	G->1	a->18	b->8	d->4	e->2	f->3	g->6	h->8	i->16	k->3	l->2	m->8	o->15	p->3	r->2	s->12	t->2	u->3	v->2	ä->13	ö->1	
tvis,	 ->6	
tvis.	 ->1	E->1	M->1	S->1	
tvisa	 ->19	,->8	.->14	?->1	n->6	r->3	
tviso	r->3	
tvist	 ->13	e->6	
tvive	l->33	
tvivl	a->10	
tvung	e->5	n->6	
tvänl	i->1	
tvärd	e->33	
tvärl	d->1	
tvärp	o->2	
tvärs	 ->1	
tvärt	o->14	
tvätt	 ->1	,->2	.->1	a->1	
två a	k->1	l->1	s->2	v->6	
två b	e->2	o->1	
två d	a->1	e->1	
två e	l->2	t->1	u->2	x->2	
två f	a->3	i->1	l->1	o->1	r->4	ö->13	
två g	r->1	å->1	
två h	a->1	u->1	
två i	n->2	r->1	
två j	o->1	
två k	o->2	r->1	ä->1	
två l	a->1	i->1	
två m	i->4	y->1	å->2	ö->1	
två n	e->1	y->1	
två o	l->1	r->1	
två p	e->1	r->3	u->8	
två r	e->1	ö->1	
två s	a->3	e->2	k->2	m->1	t->3	ä->1	
två t	i->5	r->2	y->1	
två u	n->1	p->1	t->1	
två v	e->1	i->4	
två y	t->1	
två å	r->7	s->1	
två.B	r->1	
två: 	d->2	
tvåhu	n->1	
tvång	 ->1	s->5	
ty Eu	r->1	
ty de	n->1	t->3	
ty i 	h->1	
ty na	t->1	
ty nä	r->1	
ty på	 ->2	
ty vi	 ->2	
ty är	 ->1	
ty-pr	o->1	
tycka	 ->1	,->1	s->1	
tycke	 ->7	.->3	n->1	r->59	t->1	
tyckl	i->5	
tycks	 ->8	
tyckt	e->7	
tyd g	e->1	
tyd i	 ->1	
tyd s	o->1	
tyd t	i->1	
tyd.S	a->1	
tyda 	m->1	
tydan	d->16	
tydde	 ->2	s->1	
tydel	s->73	
tyder	 ->22	,->1	:->1	
tydig	 ->1	a->3	h->4	t->3	
tydli	g->124	
tyg d	e->1	
tyg f	r->1	å->1	ö->3	
tyg i	 ->4	
tyg m	e->3	
tyg n	ä->1	
tyg o	b->1	c->1	m->1	
tyg s	o->14	å->1	
tyg u	n->2	t->1	
tyg),	 ->1	
tyg, 	d->1	s->1	u->1	
tyg.E	n->1	
tyg.F	ö->1	
tyg.V	a->1	i->1	
tyg; 	m->1	
tyg?D	ä->1	
tyga 	a->2	d->1	g->1	i->1	o->1	s->2	v->1	y->1	
tygad	 ->16	e->5	
tygan	d->5	
tygar	 ->1	
tygel	l->1	s->4	
tygen	 ->3	,->3	s->7	
tyget	 ->6	s->1	
tygsb	e->1	
tygsi	n->1	
tygss	k->7	t->1	ä->1	
tygst	a->1	
tygsä	g->1	
tympa	d->1	
tympn	i->2	
tynan	d->1	
tynga	n->1	
tyngd	 ->2	p->4	
tynge	r->1	
tyngs	t->2	
typ C	a->1	
typ a	v->18	
typ f	å->1	
typ, 	d->1	l->1	
typ.D	e->1	
typ.E	f->1	
typen	 ->12	
typer	 ->3	n->1	
typfa	l->1	
typgo	d->1	
tyr a	l->1	
tyr.E	f->1	
tyra 	d->2	e->1	f->1	g->1	h->1	m->1	u->1	ä->1	
tyran	d->4	
tyrar	 ->5	
tyras	 ->1	.->1	
tyre 	s->1	
tyre,	 ->1	
tyrek	o->3	
tyrel	s->7	
tyren	,->1	
tyret	 ->1	s->2	
tyrka	 ->7	,->1	.->1	n->4	
tyrke	f->1	p->1	
tyrko	r->2	
tyrni	n->7	
tyrs 	a->2	
tyska	 ->20	,->1	
tyskl	a->2	
tyskt	 ->2	
tyst 	m->3	
tyvär	r->30	
tz i 	B->1	
tz oc	h->1	
tz so	m->1	
tz, p	å->1	
tz. E	u->1	
tzida	k->2	
täcka	 ->5	n->4	
täcke	r->10	
täckn	i->1	
täcks	 ->4	.->1	;->1	
täckt	 ->3	s->2	
täda 	u->1	
tädat	 ->1	
täder	 ->7	,->2	.->1	n->7	
tädes	 ->1	,->1	
täkts	a->3	b->1	f->1	
tälla	 ->78	,->1	.->1	n->32	r->4	s->20	
tällb	a->1	
tälld	 ->5	a->22	e->17	h->23	
tälle	 ->2	,->1	l->7	n->3	r->41	t->50	
tälli	g->6	
tälln	i->70	
tälls	 ->18	.->2	
tällt	 ->13	,->1	.->1	s->7	
tämd 	a->1	i->1	o->1	t->1	v->1	
tämda	 ->7	,->1	
tämde	 ->5	
tämdh	e->1	
tämli	g->3	
tämma	 ->18	,->1	n->5	
tämme	l->122	r->37	
tämmi	g->4	
tämni	n->2	
tämpe	l->1	
tämpl	i->1	
täms 	u->1	
tämt 	a->2	f->2	i->1	o->1	p->1	s->4	t->1	ö->1	
tämt,	 ->3	
tän e	n->1	
tända	n->6	
tändi	g->107	
tändl	i->1	
tänga	 ->1	s->1	
tängd	e->1	
tänge	r->1	
tängn	i->6	
tängt	 ->1	
tänk 	t->1	
tänka	 ->28	,->1	n->288	s->1	
tänkb	a->3	
tänke	r->36	
tänkl	i->5	
tänks	a->2	
tänkt	 ->5	.->1	a->3	e->3	
täppa	 ->3	
täppe	r->1	
tär a	n->1	t->1	
tär f	ö->1	
tär o	c->2	
tär v	ä->1	
tär, 	a->1	
tär.R	a->1	
tära 	d->1	h->1	k->2	m->1	o->1	u->5	
tären	 ->2	
tärer	 ->1	,->1	
tärka	 ->22	,->1	n->2	s->3	
tärke	r->3	
tärkn	i->6	
tärks	 ->2	.->3	
tärkt	 ->7	a->1	s->1	
tärt 	b->1	p->1	
täta,	 ->1	
tätar	e->1	
täten	 ->2	
täthe	t->1	
täv m	e->1	
tävja	s->1	
tävla	d->1	r->1	
tävli	n->1	
tå al	l->1	
tå at	t->11	
tå av	 ->4	
tå de	 ->1	t->2	
tå en	a->1	
tå fo	l->1	
tå fr	i->1	å->7	
tå fö	r->12	
tå hu	r->2	
tå i 	k->1	p->1	s->1	v->1	
tå in	f->1	
tå kl	a->3	
tå kv	a->1	
tå ny	a->1	
tå nä	r->1	
tå oc	h->2	
tå om	 ->1	
tå so	m->1	
tå ti	l->1	
tå ut	 ->2	
tå va	r->4	
tå, a	t->1	
tå, f	ö->1	
tå, s	t->1	
tå.FP	Ö->1	
tå.Ju	s->1	
tå: å	 ->1	
tådd 	m->1	
tådda	 ->1	
tåeli	g->6	
tåels	e->8	
tåend	e->32	
tåg e	l->1	
tåg, 	v->1	
tåget	 ->1	
tågkr	a->1	
tågol	y->1	
tål a	t->1	
tålam	o->2	
tålfö	r->5	
tålge	m->1	
tålig	a->1	h->1	
tålin	d->25	
tålse	k->5	
tålst	i->1	
tålve	r->5	
tånd 	a->5	d->2	e->7	f->7	h->2	i->5	k->2	m->3	n->1	o->7	p->1	s->5	t->4	v->1	ä->1	å->1	
tånd,	 ->8	
tånd.	 ->1	A->1	D->3	F->1	H->1	J->1	V->2	
tånd?	.->1	J->1	
tånda	r->5	
tånde	l->1	n->10	t->19	
tåndi	g->1	
tåndp	u->97	
tånds	 ->1	d->12	p->2	r->1	s->1	t->2	
tår a	l->1	t->13	v->11	
tår d	e->12	ä->1	
tår e	n->2	r->3	t->1	
tår f	a->1	o->3	r->7	ö->9	
tår g	i->1	
tår h	a->1	e->6	ä->1	ö->1	
tår i	 ->22	g->1	n->21	
tår j	a->2	u->1	
tår k	l->8	o->2	
tår l	e->1	i->1	
tår m	e->1	i->2	o->1	y->3	
tår n	a->1	ä->1	
tår o	c->2	
tår p	a->1	å->13	
tår s	k->1	o->1	
tår t	i->4	
tår u	n->1	
tår v	a->3	e->1	i->4	
tår ä	v->1	
tår å	t->1	
tår ö	p->1	v->1	
tår, 	i->1	k->1	s->1	
tår.D	e->2	
tår.H	e->1	
tåret	 ->9	,->1	
tås d	ä->1	
tås f	a->1	
tås k	o->1	
tås s	k->1	
tås u	p->1	
tås v	a->1	
tåt",	 ->1	
tåtgä	r->3	
tått 	-->1	E->1	K->1	a->4	d->2	f->2	h->1	i->2	j->1	k->1	m->1	p->2	t->3	u->1	v->2	ä->1	å->1	
tått,	 ->1	
tått.	F->1	
tåtts	 ->1	
té - 	o->2	
té el	l->1	
té fö	r->3	
té ha	r->1	
té me	d->1	
té so	m->2	
téer.	D->1	
téern	a->3	
téför	f->2	
tén (	C->2	
tén f	ö->3	
tén i	 ->1	
tén k	o->1	
tén l	a->1	
tén o	c->3	m->8	
tén s	a->1	i->1	
tén v	i->1	
tén ä	r->1	
tén, 	k->1	o->1	u->1	v->1	
tén.H	u->1	
tén.M	e->1	
tén?V	i->1	
téns 	a->2	g->6	r->2	s->1	
tésys	t->2	
tête 	o->3	
tónio	 ->1	
töd -	 ->2	
töd a	n->1	v->4	
töd b	i->1	
töd d	e->2	ä->1	
töd e	f->1	n->2	
töd f	r->7	ö->19	
töd g	e->1	
töd h	a->1	o->1	
töd i	 ->5	b->1	n->5	
töd k	a->4	o->1	
töd l	ö->1	
töd m	e->2	å->3	
töd o	c->12	m->4	
töd p	e->1	r->1	å->5	
töd s	k->1	o->18	å->1	
töd t	i->43	
töd v	a->1	i->3	
töd ä	n->2	
töd å	t->2	
töd ö	k->1	
töd, 	d->1	e->1	m->1	o->3	s->7	u->1	
töd."	J->1	
töd..	(->1	
töd.A	t->1	
töd.D	e->9	å->1	
töd.E	u->1	
töd.F	ö->2	
töd.H	a->1	e->4	
töd.I	 ->2	
töd.J	a->2	
töd.M	o->1	
töd.N	i->1	
töd.O	r->1	
töd.R	e->1	
töd.S	å->1	
töd.T	r->1	
töd.U	t->1	
töd.V	i->2	
töd.Ä	n->1	v->1	
töd.Å	 ->1	r->1	
töd; 	d->1	
töd?-	 ->1	
tödde	 ->1	s->1	
töden	 ->23	,->2	.->4	s->3	
töder	 ->56	,->1	.->1	
tödet	 ->27	,->1	.->2	s->2	
tödja	 ->62	.->2	s->7	
tödje	r->1	
tödme	d->1	
tödmo	t->1	
tödni	v->1	
tödpo	l->1	
tödra	m->2	
töds 	a->5	e->1	g->1	j->1	
tödsp	o->1	
tödsy	s->4	
tödåt	g->5	
töka 	a->1	d->1	f->1	h->1	o->1	u->1	
tökad	 ->1	
tökan	d->1	
tökas	 ->1	.->1	
tökat	 ->1	
tökni	n->1	
töld,	 ->1	
tömd,	 ->1	
tömma	n->3	
tömme	r->1	
tömt 	s->1	
tör b	a->1	
tör i	 ->1	
tör k	o->1	
tör m	å->1	
tör s	y->1	
tör, 	m->1	
töra 	s->2	
töras	 ->2	!->1	
törda	 ->1	
törde	s->2	
törel	s->5	
tören	 ->1	,->1	s->1	
törer	 ->6	,->3	.->4	n->10	
törin	g->2	
törni	n->5	
törre	 ->75	
törs 	a->1	
törs,	 ->1	
törsk	å->1	
törso	m->1	
törst	 ->2	.->1	a->34	
törtn	i->1	
törts	 ->2	
töta 	p->1	
tötan	d->1	
tötar	 ->1	
töter	 ->1	
tötes	t->1	
tötfå	n->1	
tött 	B->1	F->1	d->2	p->2	s->1	u->1	v->1	ä->1	
tötta	,->1	t->1	
tötts	 ->1	
töva 	e->2	n->1	p->1	s->2	t->1	
tövan	d->1	
tövar	 ->3	
tövas	 ->4	
töver	 ->14	s->6	v->1	
tövni	n->1	
türkd	a->1	
u - a	l->1	
u 34 	s->1	
u Ahe	r->2	
u Ang	e->1	
u Ber	g->1	
u Egy	p->1	
u Eri	k->1	
u Fra	g->1	
u Lyn	n->1	
u McN	a->1	
u Mor	a->1	
u Pei	j->1	
u Plo	o->1	
u Red	i->3	
u Sch	r->3	
u Sud	r->1	
u The	a->1	
u Wal	l->1	
u abs	o->1	
u all	a->2	s->1	t->2	v->1	
u ang	r->1	
u anm	ä->1	
u ans	e->1	
u anv	ä->1	
u att	 ->8	
u av 	d->1	e->1	
u bai	n->1	
u bar	a->2	
u bef	i->1	
u beh	a->1	ö->2	
u ber	i->1	
u bet	r->1	
u bli	r->1	v->2	
u blo	t->1	
u com	b->1	
u de 	s->1	
u def	i->1	
u des	s->1	
u det	 ->1	t->2	
u dir	e->1	
u dis	k->2	
u du 	b->1	
u där	 ->1	
u då 	i->1	
u döp	e->1	
u eft	e->1	
u ege	n->1	
u eme	l->1	
u en 	a->1	f->1	g->9	n->1	t->1	
u ett	 ->8	
u eur	o->1	
u fak	t->1	
u fat	t->1	
u fin	n->4	
u fle	x->1	
u fra	m->1	
u frå	g->1	n->1	
u får	 ->2	
u fåt	t->2	
u fög	a->1	
u för	 ->5	e->5	k->1	o->1	s->3	v->1	
u gem	e->1	
u gen	o->1	
u ger	 ->2	
u get	t->1	
u gäl	l->3	
u gå 	i->2	t->1	
u gån	g->1	
u gör	a->3	
u har	 ->18	,->1	
u hot	a->1	
u här	 ->1	
u hål	l->1	
u hår	d->2	
u hög	r->4	
u hör	 ->1	
u i T	u->1	
u i p	r->1	
u i s	a->1	
u i v	a->1	
u ige	n->1	
u inb	j->1	
u ind	i->1	
u ing	e->2	
u inl	e->1	
u inn	e->3	
u ino	m->1	
u ins	p->1	
u int	e->40	
u iso	l->1	
u kan	 ->6	d->1	
u kom	m->51	
u kon	k->1	
u led	a->2	
u lig	g->1	
u lys	s->1	
u läg	g->1	
u län	g->1	
u läs	e->1	
u lät	t->1	
u med	 ->20	,->2	d->1	
u men	 ->1	
u mer	 ->9	.->2	
u mig	 ->1	
u min	d->2	
u mor	d->1	
u mär	k->1	
u mås	t->10	
u num	m->1	
u när	 ->8	
u nåt	t->1	
u och	 ->6	
u ock	s->8	
u off	i->1	
u oft	a->2	
u oms	ä->1	
u par	l->1	
u pla	n->1	
u por	t->1	
u pri	o->1	
u prö	v->1	
u pun	k->1	
u på 	a->1	e->1	
u på.	D->1	
u påg	å->2	
u red	a->2	
u res	o->1	
u rul	l->1	
u råd	a->1	e->1	
u rös	t->1	
u sa 	a->1	
u sad	e->2	
u sam	m->2	t->1	
u ser	 ->1	
u ses	 ->1	
u sif	f->1	
u sin	 ->1	
u ska	l->4	
u ske	r->1	
u sku	l->1	
u skö	r->1	
u slå	 ->1	
u smi	d->1	
u som	 ->2	
u spe	c->1	
u sta	r->1	
u str	ä->1	
u stä	d->1	m->1	n->1	
u stå	r->3	
u stö	d->2	r->4	
u svå	r->1	
u säg	e->1	
u sät	t->1	
u så 	a->1	l->1	
u tag	i->2	
u tal	a->1	m->83	
u tar	 ->2	
u til	l->5	
u tyd	l->2	
u tyv	ä->1	
u und	e->1	
u upp	 ->1	s->1	t->1	
u utt	r->1	
u vad	 ->1	
u vem	 ->1	
u ver	k->2	
u vid	 ->1	t->1	
u vik	t->2	
u vil	l->2	
u vis	s->1	
u vän	t->1	
u äld	r->1	
u än 	f->1	
u änd	r->1	å->1	
u änt	l->5	
u är 	a->1	d->6	e->2	f->2	h->2	i->2	m->1	n->1	o->1	p->1	r->1	s->2	u->1	
u är,	 ->1	
u åte	r->2	
u", d	v->1	
u, La	n->1	
u, an	a->1	
u, ef	t->2	
u, en	 ->1	
u, ha	r->1	
u, i 	j->1	
u, me	n->2	
u, oc	h->2	
u, pr	e->1	
u, si	n->1	
u, so	m->2	
u, un	d->1	
u, åt	t->1	
u, öv	e->1	
u-län	d->1	
u..Ta	c->1	
u.Det	 ->1	
u.Ett	 ->1	
u.Jag	 ->1	
u.Kom	m->1	
u.Kon	s->1	
u.Låt	 ->1	
u.Vi 	a->1	g->1	
u: gö	r->1	
u; i 	d->1	
u?Jag	 ->1	
uMed 	h->1	
ua no	n->2	
uades	 ->1	
ual D	e->1	
ual h	a->1	
ual s	o->1	v->1	
ual v	a->1	
ual ä	r->1	
ual" 	o->1	
ual, 	o->1	
ualis	e->2	
ualit	e->1	
uanze	s->1	
uari 	1->4	2->5	e->1	f->1	i->3	m->1	n->1	o->3	
uari!	H->1	
uari,	 ->10	
uari.	H->1	V->1	
uatem	a->1	
uatio	n->129	
ubba 	a->1	
ubbar	 ->1	
ubbas	 ->1	
ubbel	 ->1	s->2	t->2	v->1	
ubbla	 ->10	s->1	
ubetä	n->1	
ubikm	e->2	
ubjek	t->1	
ublan	d->1	
ublic	 ->1	e->4	i->1	
ublik	 ->2	a->6	e->12	
ublin	 ->4	.->1	k->2	
ubrik	e->2	
ubsid	a->1	i->22	
ubsta	n->4	
ubven	t->12	
uc se	r->1	
ucces	s->5	
ucent	 ->2	a->6	e->14	
ucera	 ->4	d->1	r->2	s->2	t->3	
uceri	n->1	
uchne	r->12	
ucka 	i->1	
ucka"	,->1	
ucka,	 ->1	
uckit	 ->1	
uckne	s->1	
uckor	 ->2	
uctor	i->1	
ud 7 	p->1	
ud Ba	r->2	
ud el	l->1	
ud fa	t->1	
ud fö	r->4	
ud me	d->2	
ud mo	t->7	
ud oc	h->4	
ud re	s->1	
ud ta	g->9	
ud vi	 ->1	
ud är	 ->1	
ud, a	m->1	
ud, e	t->1	
ud, h	u->1	
ud, s	o->1	
ud.De	t->2	
ud.Va	d->1	
uda a	l->1	
uda b	e->2	å->1	
uda d	e->1	
uda e	n->2	t->1	
uda i	n->1	
uda k	o->1	
uda m	ö->1	
uda n	å->1	
uda o	s->1	
uda p	h->1	
uda u	t->1	
udakt	ö->2	
udan 	f->1	
udand	e->4	
udang	e->1	
udans	v->4	
udape	s->1	
udars	 ->1	
udas,	 ->1	
udas.	T->1	
udda 	k->1	u->1	
uddel	 ->1	e->2	
uddhi	s->1	
uddig	h->1	t->1	
ude M	a->1	
uden 	t->1	
udent	e->1	s->1	
uder 	a->1	e->1	f->1	g->1	i->1	l->1	m->1	o->1	r->2	v->1	
uder,	 ->1	
udera	 ->1	r->3	t->3	
udet 	M->1	h->2	i->1	m->3	s->1	u->1	v->2	
udet,	 ->1	
udet.	D->1	
udet?	N->1	
udeut	r->1	
udfrå	g->4	
udför	s->1	
udget	 ->9	,->4	.->6	a->3	b->1	e->16	f->11	k->17	m->1	p->14	s->4	u->10	å->10	ö->1	
udice	r->1	
udie 	o->1	
udieb	e->1	
udiep	r->1	
udier	 ->4	,->1	.->1	
udika	t->3	
udisk	a->1	
udit 	F->1	
udlig	t->1	
udlin	j->2	
udmål	e->1	s->1	
udna 	m->1	s->1	
udnin	g->1	
udord	e->1	
udre 	o->1	
udre,	 ->1	
udrek	o->1	
udrol	l->2	
udron	 ->1	
uds s	k->2	
udsak	 ->6	l->10	
udsfö	r->3	
udsin	f->2	r->1	
udska	p->10	
udsma	n->10	
udspr	i->1	
udsta	d->2	
udstä	d->2	
udsyf	t->1	
udupp	g->1	
ue ka	n->1	
ue, s	o->1	
ue, v	a->1	
ueced	o->1	
ueira	 ->1	
uela 	e->1	
uell 	e->1	f->1	i->1	l->1	o->3	r->1	u->1	
uell.	A->1	D->1	S->1	Ä->1	
uella	 ->36	,->1	.->1	
uellt	 ->14	,->1	.->1	
uen, 	S->1	
uer h	a->1	
uer s	a->1	
uer t	a->1	
uer, 	n->1	
uera 	d->1	e->3	o->1	
uerad	e->1	
uerar	 ->1	
uerat	s->1	
uerli	g->2	
uernt	u->1	
ues D	e->3	
ues e	t->1	
ues".	K->1	
uesa 	o->1	
uff n	o->1	
uffar	e->1	
ufman	n->1	
uft g	e->1	
uft.V	i->1	
uftbu	r->1	
uftet	 ->1	
uftig	 ->3	a->2	t->6	
uftom	r->1	
uföra	 ->1	
uga, 	f->1	
ugal 	K->1	b->1	k->1	o->9	p->1	t->1	ä->1	
ugal,	 ->4	
ugals	 ->7	
ugare	 ->1	
ugen 	s->1	
ugen.	H->1	
uger 	i->1	
ugg p	å->3	
ugga 	o->1	
uggan	 ->1	
uggbo	x->1	
uggen	"->1	
uggli	n->1	
ugisi	s->70	
uglig	a->5	h->1	
ugn o	c->1	
ugna 	m->1	n->1	
ugnad	e->1	
ugnan	d->1	
ugnas	.->1	
ugo g	r->1	
ugo å	r->1	
ugofe	m->1	
ugond	e->1	
ugor,	 ->1	
ugosl	a->1	
ugues	a->1	
uhame	l->1	
uhe o	c->1	
uhe, 	L->1	
uhne,	 ->1	
uierd	o->1	
uigou	 ->1	
uiner	a->1	
uins 	r->1	
uiola	 ->1	
uisen	b->3	
uisit	i->1	
uita 	o->1	
uiz s	o->1	
uk al	-->1	
uk av	 ->1	
uk me	l->1	
uk oc	h->5	
uk på	 ->1	
uk so	m->1	
uk!An	d->1	
uk, d	e->3	
uk, e	x->1	
uk, i	 ->1	
uk, m	e->1	
uk, t	i->1	r->1	
uk, v	i->1	
uk.Ja	g->1	
uka P	V->1	
uka, 	s->1	
ukade	 ->1	s->1	
ukar 	d->1	e->1	o->1	
ukar:	 ->1	
ukare	 ->5	,->1	n->1	s->1	
ukarn	a->5	
ukas 	ö->1	
ukas.	H->1	
ukasu	s->3	
ukdom	 ->1	
uken.	D->1	
uket 	(->2	-->1	a->1	f->3	i->2	k->1	o->2	s->1	
uket,	 ->2	
uket.	D->1	
uket;	 ->2	
ukets	 ->1	
ukför	s->1	
ukhus	 ->1	,->2	.->1	e->2	l->1	
ukits	 ->1	
uknin	g->3	
uksek	o->1	
uksfo	n->1	
uksfr	å->1	
ukslo	b->1	
uksom	r->2	
ukspo	l->6	
ukspr	i->1	o->2	
uksre	f->1	g->1	
uksse	k->5	
ukssy	n->1	
ukt a	v->2	
ukt h	a->1	
ukt p	å->1	
ukt s	k->1	o->2	
ukt, 	u->1	
ukt.H	e->1	
uktan	 ->1	s->6	
uktar	 ->2	,->1	.->1	
uktat	 ->1	
uktba	r->2	
ukten	 ->6	.->1	
ukter	 ->5	,->1	.->2	n->2	
uktig	a->1	
uktin	n->1	
uktio	n->39	
uktiv	 ->1	a->10	i->4	t->6	
uktor	i->6	
ukts 	l->1	o->1	
uktur	 ->15	,->4	.->3	b->1	e->51	f->58	m->1	n->1	p->12	r->1	s->3	u->2	å->1	
uktör	e->3	
ukvår	d->3	
ul fö	r->1	
ul oc	h->1	
ul om	 ->1	
ul so	m->1	
ul.Vi	 ->1	
ula o	m->1	
ula ö	v->1	
ula.J	a->1	
ulada	k->1	
ulans	 ->2	e->2	å->1	
ulari	s->1	
ulary	 ->1	
ulati	o->10	v->2	
ulato	r->2	
ulda 	d->1	
uldan	d->1	
uldbe	l->1	
ulden	 ->2	
ulder	 ->1	
ulen 	ä->1	
uler 	f->1	o->1	ä->1	
ulera	 ->28	"->1	,->1	d->4	r->13	s->4	t->4	
uleri	n->6	
ulf-M	a->2	
ulfer	i->1	
ulfkr	i->1	
ulgar	i->1	
uli 1	9->4	
uli 2	0->2	
uli f	ö->1	
uli u	n->1	
uli, 	m->1	o->1	
ulism	.->1	
uliss	e->1	
ulist	i->2	s->1	
ulkla	p->1	
ull a	p->1	v->1	
ull b	e->2	o->1	
ull e	u->1	
ull f	å->1	ö->1	
ull g	e->2	å->2	
ull h	a->1	ä->2	
ull i	n->2	
ull n	y->1	
ull o	m->1	
ull p	r->1	
ull r	e->1	o->1	
ull s	k->2	t->1	
ull v	o->1	
ull ä	r->1	
ull ö	p->1	
ull, 	j->1	n->1	s->1	
ull.D	e->3	
ull.K	o->1	
ull.O	r->1	
ull.V	i->1	
ulla 	a->3	f->2	i->2	k->1	l->1	o->1	s->7	u->1	v->1	
ulla,	 ->1	
ulla.	D->1	V->1	
ullar	 ->3	.->1	e->1	n->1	
ullas	t->1	
ullbo	r->3	
ulle 	E->3	K->1	a->7	b->20	d->40	e->8	f->24	g->16	h->21	i->24	j->44	k->65	l->5	m->4	n->3	o->9	p->4	r->5	s->28	t->13	u->14	v->120	ä->2	å->2	ö->2	
ulle,	 ->2	
ullfö	l->3	r->1	
ullgj	o->1	
ullgå	v->1	
ullgö	r->1	
ullhe	t->1	
ullit	e->1	
ullka	s->1	
ullko	m->5	
ullo 	g->1	i->1	o->1	r->1	å->1	
ullst	o->3	ä->41	
ullt 	a->2	b->3	d->3	e->1	f->3	g->1	i->3	k->2	m->3	o->5	p->1	s->1	t->1	u->11	
ullt,	 ->1	
ullt.	D->1	H->1	
ullvä	r->2	
ullän	d->2	
ulor 	o->1	
ulos 	f->1	o->4	
uls f	ö->1	
uls t	i->1	
ulser	 ->4	
ulska	 ->1	
ult d	r->1	
ult k	o->1	
ultat	 ->31	,->6	.->10	:->1	?->2	e->44	i->3	l->1	t->7	ö->6	
ultba	s->1	
ulten	 ->7	!->2	,->1	.->3	b->4	s->3	
ulter	 ->1	a->8	
ulthe	n->6	
ultie	t->3	
ultil	a->1	
ultim	a->1	
ultin	a->5	
ultra	l->1	p->1	
ultur	 ->41	,->11	-->1	.->3	?->1	a->8	e->64	f->1	h->1	o->1	p->8	s->5	u->1	
ulz e	n->1	
ulz s	a->2	
uläge	t->1	
ulära	 ->2	
ulärt	 ->1	
um - 	o->1	
um at	t->56	
um av	 ->2	g->1	
um bl	i->1	
um då	 ->1	
um eg	e->1	
um en	 ->1	
um fi	n->1	
um fr	a->1	
um fö	r->9	
um ha	d->1	r->1	
um hä	r->1	
um i 	B->1	G->1	e->1	m->13	p->1	
um in	f->3	t->2	
um me	d->2	
um mi	n->1	
um må	s->1	
um oc	h->9	
um om	 ->3	
um på	 ->4	
um sk	j->1	u->1	
um so	m->6	
um un	d->1	
um ut	a->1	
um vä	g->1	
um yt	t->1	
um än	 ->1	
um är	 ->3	,->1	
um ås	a->1	
um åt	g->1	
um!De	t->1	
um!Me	n->1	
um, b	ö->1	
um, d	e->1	å->1	
um, k	a->1	r->1	
um, m	e->1	
um, o	c->3	
um, p	å->1	
um, u	t->1	
um, v	i->1	
um. D	ä->1	
um.At	t->1	
um.Av	 ->1	
um.De	n->1	t->3	
um.He	r->1	
um.I 	d->1	
um.Lå	t->1	
um.Me	n->1	
um.OM	R->1	
um.Pr	o->1	
um.Rå	d->1	
um.So	m->1	
um.Vi	 ->2	
um.Än	d->1	
uman 	r->1	
umani	s->3	t->2	
umar 	P->1	
umati	s->1	
umbar	 ->1	
umbär	l->4	
ument	 ->78	,->9	.->7	a->3	e->60	f->6	k->1	o->1	p->2	r->1	s->5	t->1	v->2	
umera	 ->6	
umet 	a->2	b->1	f->2	
umet.	D->1	
umgän	g->1	
umhet	 ->2	,->1	
umlen	,->1	
umma 	h->1	p->3	s->1	
ummad	e->1	
umman	 ->2	
ummat	 ->1	
ummel	s->6	
ummer	 ->1	,->1	
ummip	a->1	
ummor	 ->7	.->1	
ump a	t->2	
ump s	j->1	
ump.D	e->1	
umpan	d->1	
umpas	 ->2	
umper	a->2	
umpni	n->3	
umra 	i->1	
umt a	t->1	
umtan	k->1	
umtio	n->2	
umula	t->1	
umule	r->1	
umäni	e->1	
umör 	s->1	v->1	
un sa	d->1	
un.De	n->1	
una p	e->1	
una ä	r->1	
unala	 ->2	
unalp	a->1	
unans	 ->1	
unc d	å->1	
uncht	i->1	
uncil	 ->1	
und (	k->1	r->1	
und L	T->1	
und a	t->2	v->79	
und e	l->1	
und f	i->1	ö->16	
und i	 ->2	n->1	
und o	c->1	
und s	e->6	k->1	
und t	i->1	
und u	p->1	
und v	e->1	i->1	
und ä	r->2	
und, 	m->1	o->1	
und.D	e->1	
und.N	i->1	
und.P	å->1	
und? 	H->1	
unda 	-->1	a->3	b->1	d->2	e->1	f->5	h->1	i->1	n->1	o->1	s->2	
unda,	 ->1	
unda.	B->1	K->1	
undad	 ->5	e->3	
undam	e->1	
undan	 ->7	,->1	b->2	d->3	f->1	h->1	m->1	r->6	t->36	
undar	 ->3	e->1	
undas	 ->6	
undat	 ->5	
undbu	l->1	
unde 	a->3	b->3	d->1	f->2	g->1	h->1	k->3	m->1	p->1	s->5	u->1	v->5	ö->4	
unden	 ->34	,->2	.->6	
under	 ->313	,->2	.->1	a->12	b->3	g->4	h->5	k->4	l->33	m->3	n->2	o->4	r->3	s->90	t->17	u->1	v->1	
undet	 ->10	,->3	s->1	
undfö	r->4	
undgä	n->2	
undgå	t->1	
undi 	r->1	s->1	
undi:	 ->1	
undit	 ->3	
undku	r->1	
undli	g->16	
undlä	g->74	
undna	 ->4	
undor	s->1	
undpe	l->1	
undpr	i->1	
undra	 ->5	d->8	n->2	r->9	t->9	
undre	s->2	
undri	n->1	
undsa	t->1	
undsj	u->1	
undsk	a->1	
undsl	ä->2	
undsr	e->5	
undst	e->1	
undte	s->1	
undva	g->1	l->24	t->1	
undvi	k->39	
undär	r->1	
uner 	k->1	o->1	s->4	ä->1	
unera	d->1	
unern	a->2	
uners	 ->1	
ung a	r->1	
ung b	y->1	
ung m	a->1	
ung o	c->2	l->1	
ung p	o->1	r->1	
ung u	p->1	
ung. 	S->1	
ung.I	 ->1	
ung.O	c->1	
unga 	f->1	k->2	m->2	o->1	
unga,	 ->2	
ungan	d->1	
ungar	i->15	
ungdo	m->14	
ungef	ä->8	
ungel	n->2	
ungen	 ->5	
unger	a->54	
unget	 ->1	,->1	
ungfr	u->1	
ungli	g->13	
ungme	t->6	
ungna	 ->6	
ungro	d->1	
ungsl	a->1	
ungt 	h->1	
ungt,	 ->1	
unhas	 ->1	
uni 1	9->6	
uni 2	0->2	
uni f	ö->2	
uni i	 ->1	
uni v	a->1	
unice	r->2	
unika	 ->1	t->16	
unikt	 ->1	
unila	t->2	
union	 ->13	,->5	.->6	e->406	s->7	
unism	 ->1	,->1	
unist	e->1	
unite	t->1	
unive	r->4	
unka 	a->1	b->1	n->1	
unka.	Å->1	
unker	 ->1	,->1	s->1	
unkit	 ->2	
unkla	t->1	
unkna	 ->1	d->1	r->1	t->1	
unkt 	(->2	-->2	1->3	2->3	4->2	5->1	6->1	7->1	D->1	a->4	b->1	d->4	e->2	f->6	g->3	h->4	i->16	k->2	m->4	n->2	o->6	p->29	r->1	s->20	t->2	u->1	v->2	ä->8	
unkt,	 ->14	
unkt.	 ->1	A->1	D->5	I->1	M->3	N->2	P->1	T->2	V->3	
unkt:	 ->2	
unkt?	E->1	
unkte	n->88	r->85	
unkti	o->32	
unkts	 ->1	p->1	
unktu	r->1	
unna 	a->9	b->18	d->6	e->1	f->33	g->26	h->8	i->7	k->5	l->12	m->5	n->2	o->3	p->5	r->3	s->21	t->12	u->16	v->10	y->1	ä->2	å->6	
unna.	V->1	
unnan	d->2	
unnar	 ->2	
unnat	 ->43	
unnel	n->2	t->1	
unnen	 ->2	
unnet	 ->1	
unnig	 ->2	a->1	h->2	t->1	
unnit	 ->6	,->1	.->1	s->8	
unnla	r->2	
unnor	 ->1	
uno L	e->1	
unska	p->17	
unt o	c->1	m->2	
unt t	i->1	
unt.D	e->1	
unta 	i->2	
untar	 ->1	i->4	
untli	g->8	
untom	 ->1	
untor	 ->1	
untpr	a->1	
untra	 ->6	d->1	n->3	r->8	s->3	
uo so	m->1	
uo, d	ä->1	
up , 	m->1	
up de	 ->1	
up ön	s->1	
upa f	o->1	
upa m	i->1	
upa o	c->1	
upa s	y->1	
upa u	n->1	
upa, 	p->1	
upad 	a->1	
upant	e->1	
upare	 ->1	
upas 	b->1	
upast	e->2	
upat 	s->2	
upati	o->1	
upera	d->2	t->1	
upet 	-->1	i->1	p->1	
upet,	 ->2	
upgåe	n->7	
upnin	g->5	
upp (	k->2	
upp -	 ->1	
upp E	u->1	
upp T	i->1	
upp a	l->4	n->4	t->3	v->9	
upp b	e->2	i->1	å->1	
upp d	e->40	o->1	
upp e	f->3	l->1	n->10	t->6	x->1	
upp f	o->1	r->10	u->1	ö->5	
upp g	e->2	r->1	
upp h	a->4	e->1	u->1	ä->3	
upp i	 ->17	d->1	g->4	n->2	
upp k	o->6	
upp l	a->1	i->1	ä->3	
upp m	e->8	å->1	
upp n	a->1	y->1	å->3	
upp o	c->5	l->1	m->1	r->2	
upp p	o->1	r->3	å->8	
upp r	e->2	ä->3	ö->1	
upp s	a->1	i->2	k->3	o->5	t->2	ä->2	å->1	
upp t	i->11	o->1	r->1	v->1	y->2	
upp u	n->2	t->6	
upp v	a->3	i->2	ä->2	
upp ä	n->2	r->7	
upp, 	E->1	a->1	d->1	e->4	f->1	h->2	j->1	m->2	n->1	o->1	r->1	s->3	v->1	
upp.A	h->1	
upp.D	e->4	
upp.F	a->1	
upp.J	a->7	
upp.M	e->1	
upp.P	å->1	
upp.V	i->2	
upp.Ä	n->1	v->1	
upp?H	u->1	
uppba	c->1	
uppbr	i->3	
uppby	g->20	
uppbä	r->1	
uppbå	d->1	
uppda	t->2	
uppde	l->3	
uppdr	a->22	
uppeh	å->13	
uppen	 ->44	,->3	.->3	b->35	s->13	
upper	 ->24	,->4	.->4	a->1	i->2	n->21	s->1	
uppfa	n->1	t->51	
uppfy	l->54	
uppfö	d->1	l->9	r->13	
uppgi	c->3	f->74	
uppgr	a->1	
uppgå	 ->1	n->2	r->5	
uppgö	r->2	
upphe	t->1	
uppho	v->13	
upphä	v->5	
upphö	j->1	r->9	
uppko	l->1	m->6	
upple	v->17	
uppli	v->1	
upply	s->4	
upplö	s->3	
uppma	n->58	
uppmj	u->2	
uppmu	n->21	
uppmä	r->53	t->2	
uppnå	 ->49	,->1	.->4	d->6	r->13	s->7	t->13	
uppor	d->1	
uppre	n->2	p->52	
uppri	k->6	
uppro	p->5	
uppru	s->1	
uppry	c->1	
upprä	c->2	k->1	t->35	
upprö	r->5	
upps 	u->1	v->3	
uppsa	m->4	t->3	
uppsk	a->23	j->4	o->2	
uppsp	å->2	
uppst	o->4	ä->3	å->32	
uppsä	g->1	t->2	
uppta	g->7	r->1	s->2	
uppti	l->1	
uppto	g->2	
upptr	ä->10	
upptä	c->11	
uppun	d->1	
uppvi	g->1	s->5	
uppvä	g->1	r->1	
upran	a->1	
upsin	n->1	
upskh	e->1	
upt b	e->2	
upt d	i->1	
upt o	r->1	
upt s	k->1	
upt v	a->1	
upt ö	v->1	
uptio	n->7	
upéry	s->1	
uqal 	f->1	ä->1	
ur - 	d->1	o->1	
ur 20	0->20	
ur EG	:->1	
ur EU	:->1	
ur Eu	r->2	
ur UC	L->1	
ur al	l->1	
ur an	s->1	v->1	
ur ar	b->1	
ur av	f->1	
ur ba	r->1	
ur be	k->1	s->3	v->1	
ur bi	l->2	
ur br	a->1	u->1	å->2	
ur bu	d->2	
ur by	x->1	
ur de	 ->8	l->1	n->15	r->2	s->5	t->15	
ur di	s->1	
ur dr	a->1	
ur dä	r->1	
ur ek	o->2	
ur en	 ->7	k->1	
ur er	 ->1	
ur et	t->5	
ur fa	t->1	
ur fo	l->1	r->1	
ur fr	a->1	
ur fö	r->11	
ur ge	n->1	
ur go	t->1	
ur gå	r->1	
ur gö	r->1	
ur ha	n->1	r->2	
ur ho	t->2	
ur hö	g->1	
ur i 	E->1	k->1	
ur in	f->1	t->3	
ur jo	r->1	
ur ka	n->2	
ur kl	o->3	
ur ko	m->9	s->1	
ur ku	l->1	
ur kä	n->1	
ur le	d->1	
ur li	g->1	t->1	
ur lä	g->2	n->1	
ur lå	n->5	
ur ma	n->17	r->1	t->1	
ur me	d->1	
ur mi	l->4	n->2	
ur my	c->1	n->1	
ur mä	n->1	
ur må	n->7	
ur ni	 ->2	,->1	
ur nu	 ->2	
ur oc	h->9	
ur of	t->1	
ur pa	r->1	s->2	
ur pe	n->1	r->1	
ur po	l->1	
ur pr	o->2	
ur på	 ->1	
ur ri	s->1	
ur sa	m->1	
ur se	r->3	
ur si	k->1	
ur sk	a->11	
ur sm	å->1	
ur sn	a->1	
ur so	m->19	
ur st	a->3	o->7	r->1	ö->1	
ur sv	a->1	å->4	
ur sä	r->1	
ur sö	d->1	
ur te	k->1	
ur ti	b->1	
ur tr	a->1	
ur tu	s->1	
ur tä	n->1	
ur un	d->1	i->2	
ur up	p->1	
ur ur	v->1	
ur ut	a->1	b->1	f->1	v->1	
ur ve	r->1	
ur vi	 ->21	k->6	l->3	
ur vä	l->1	x->1	
ur vå	r->1	
ur är	 ->6	
ur, (	B->1	
ur, G	a->1	
ur, a	n->1	t->1	v->1	
ur, f	ö->1	
ur, h	ö->1	
ur, l	i->1	
ur, m	e->2	i->1	
ur, o	c->2	m->1	
ur, s	i->1	
ur, t	r->2	
ur, u	n->3	
ur, å	t->1	
ur- o	c->4	
ur.De	 ->1	t->2	
ur.Dä	r->1	
ur.Fo	l->1	
ur.He	r->1	
ur.Ko	m->1	
ur.Ni	 ->1	
ur.Om	 ->1	
ur.Rå	d->1	
ur.Ty	v->1	
ur.Vi	 ->3	
ur?Me	n->1	
ura f	ö->3	
ura o	c->1	
ura s	o->1	å->1	
ura, 	d->1	s->1	
ura.D	e->1	
urakt	i->1	
urali	s->1	
uran 	H->1	a->1	h->1	
uran.	D->1	
uran?	O->1	
urani	u->2	
urans	l->1	
uranv	a->4	
urar 	o->1	
urarb	e->1	
urarn	a->1	
urart	e->1	
urarv	 ->1	,->2	.->1	e->1	
uras 	a->1	
urat 	F->1	
urato	m->4	
urban	i->1	
urbes	t->1	
urd i	v->1	
urell	 ->10	a->22	t->8	
uren 	b->2	d->2	e->2	f->3	h->2	i->6	k->2	o->8	p->1	s->3	t->2	u->1	ä->3	
uren,	 ->5	
uren.	D->2	R->1	T->1	
uren?	I->1	
urens	 ->8	
urer 	a->1	i->1	k->1	o->3	p->1	s->4	å->1	
urer,	 ->4	
urer.	D->1	E->1	K->1	V->1	
urera	 ->1	d->4	t->1	
ureri	n->10	
urern	a->6	
urers	 ->1	
ures 	e->1	
uret 	h->1	o->1	
urfod	e->4	
urfon	d->58	
urfor	m->1	
urför	t->2	
urg f	i->1	
urg i	 ->1	
urg m	e->2	
urg u	t->1	
urg ö	p->1	
urg, 	B->1	I->1	f->1	j->1	
urg.D	e->1	
urg.J	a->1	
urg.L	e->1	
urg.V	i->1	
urgar	e->1	
urgh.	V->1	
urhis	t->1	
urhol	k->4	
uri.B	å->1	
uridi	s->30	
urie-	s->1	
urien	.->1	
uris 	h->1	l->1	o->1	ä->1	
uris.	J->1	
urisd	i->5	
urism	 ->9	,->4	.->3	e->4	
urist	e->8	i->1	s->2	
urit 	p->1	
urita	n->1	
urk-d	a->1	
urkar	,->1	n->1	
urkat	a->13	
urkie	t->35	
urkis	k->6	
urkme	n->2	
urlan	g->6	
urlig	a->3	t->99	
urliv	,->1	.->1	
urmin	n->1	
urmäs	s->1	
urna.	D->1	
urnal	i->2	
urner	i->1	
urnät	e->1	
urnöd	v->1	
uro 1	9->1	
uro b	e->1	
uro f	ö->6	
uro h	a->1	
uro i	 ->1	
uro o	c->1	
uro p	e->2	å->1	
uro t	i->1	
uro u	n->1	
uro!A	l->1	
uro, 	f->1	h->1	k->1	o->2	s->2	v->1	
uro-r	å->1	
uro.D	e->2	ä->1	
uro.H	u->1	
uro.K	n->1	
uro.N	ä->1	
uro.S	e->1	
uro.V	i->1	
uroda	c->5	
urofe	d->1	
uroju	s->6	
uromr	å->2	
uron 	e->1	o->1	s->1	
uron,	 ->1	
urons	 ->3	
uroom	r->1	
uropa	 ->141	!->2	"->1	,->36	.->60	;->1	?->3	N->1	d->2	g->1	k->1	m->1	n->1	p->166	r->1	s->46	t->1	v->3	
urope	i->712	
uropo	l->16	
uropr	o->1	
uropé	 ->1	e->9	
urosk	e->3	
urost	a->1	
urpol	i->16	
urpro	g->3	j->1	
urref	o->1	
urreg	l->1	
urren	s->278	t->2	
urrer	a->5	
urs d	u->1	
urs i	 ->1	
urs m	e->1	å->1	
urs o	c->1	
urs, 	o->1	
urs.D	e->1	
ursbr	i->1	
ursek	t->5	
ursen	 ->3	,->1	
urser	 ->26	,->3	.->7	n->16	
ursfö	r->1	
urski	l->3	
ursku	l->1	
urspr	u->19	
urspå	r->1	
urssl	ö->1	
ursti	l->1	
urstö	d->3	
ursäk	t->14	
ursän	d->1	
urt a	t->1	
urt m	o->1	
urtz 	o->1	s->1	
urtz,	 ->1	
urutg	i->1	
uruts	k->1	
urutv	e->1	
uruvi	d->15	
urval	 ->3	e->1	s->1	
urvat	t->8	
urvet	e->1	
urvis	 ->1	
uråtg	ä->1	
us 19	9->1	
us 20	 ->1	
us an	m->1	
us av	 ->1	
us be	t->3	
us en	 ->1	l->1	
us fy	r->1	
us fö	r->1	
us ha	r->1	
us ju	r->5	
us ka	n->1	
us kr	ä->1	
us oc	h->2	k->1	
us på	 ->1	
us qu	o->2	
us so	m->1	
us st	a->1	
us tj	u->1	
us tr	e->1	
us un	d->1	
us är	 ->1	
us, e	f->1	
us, f	ö->1	
us, h	e->1	
us, m	e->1	y->1	
us-be	s->1	
us.De	t->2	
us.Eu	r->1	
us.Ge	n->1	
us.He	r->1	
us.In	t->1	
us?Oc	h->1	
usa v	i->1	
usale	m->2	
usar 	i->1	å->1	
uschw	i->1	
usdim	e->1	
use",	 ->1	
useff	e->3	
usen 	E->1	b->1	d->1	o->1	t->1	
usen,	 ->1	
usend	e->3	
usent	a->10	
usera	 ->1	r->1	t->1	
uset 	-->1	a->5	i->3	p->1	
uset.	J->1	
usewi	e->1	
usför	h->1	
usgas	e->4	
usgra	d->2	
ush P	o->1	
ush, 	a->1	
ushål	l->1	
usias	m->3	
usik 	i->1	m->1	
usike	n->1	r->1	
usion	 ->1	e->4	s->3	
usiv 	r->1	
usiva	 ->1	
usive	 ->17	
usivt	 ->1	
usk.H	e->1	
uskou	r->1	
usläk	a->1	
usp",	 ->1	
uspen	s->1	
usqui	n->1	
ussa 	t->1	
ussag	 ->1	
ussar	 ->1	,->1	
ussas	 ->1	
ussel	-->1	o->1	
ussen	 ->1	
ussin	 ->1	
ussio	n->61	
ussla	 ->1	n->1	
ust a	l->1	n->1	t->1	
ust b	e->1	i->1	l->1	
ust d	e->14	ä->4	
ust e	f->1	t->1	
ust f	l->1	r->1	ö->10	
ust g	e->1	j->2	
ust h	a->12	ä->3	
ust i	 ->6	
ust l	ä->2	
ust m	e->3	
ust n	u->10	ä->4	
ust o	f->1	
ust p	r->1	å->5	
ust r	ö->1	
ust s	a->4	k->2	o->2	
ust v	a->1	i->2	
ust ö	v->1	
ust, 	d->1	
ust.D	e->1	
ust.K	o->1	
ust.V	i->1	
ust: 	m->1	
usta 	d->1	
ustaa	f->1	
ustad	 ->2	
ustbe	s->1	v->1	
ustbr	i->1	
usten	 ->9	,->4	.->4	N->1	
uster	 ->4	.->2	a->5	i->3	n->7	
ustic	e->4	
ustit	i->6	
ustli	n->2	
ustmy	n->3	
ustni	n->5	
ustom	r->2	
ustra	t->1	
ustre	g->1	r->1	
ustri	 ->11	,->3	-->1	e->8	f->4	l->2	n->80	p->2	s->3	
ustva	k->1	
usul 	o->1	s->1	
usul.	V->1	
usule	r->3	
usí ä	r->1	
usöve	r->1	
ut - 	o->1	
ut 10	 ->1	
ut 88	/->2	
ut 94	/->1	
ut To	t->1	
ut ac	c->1	
ut am	e->1	
ut an	s->2	
ut at	t->8	
ut av	 ->3	
ut be	h->2	k->1	r->1	
ut bo	r->1	
ut bö	r->2	
ut de	m->1	n->5	t->1	
ut di	s->1	
ut en	 ->5	
ut et	t->2	
ut ex	p->1	
ut fa	t->1	
ut fo	k->1	
ut fr	a->1	å->8	
ut fö	r->9	
ut ge	n->1	
ut go	d->1	
ut ha	m->1	n->2	r->3	
ut hö	g->1	
ut i 	P->1	d->1	f->2	k->3	r->1	s->1	v->1	
ut in	o->2	t->8	
ut ka	n->2	
ut ko	m->1	n->1	
ut ku	n->1	
ut la	d->1	
ut ly	c->1	
ut lä	n->1	
ut lå	t->1	
ut me	d->4	
ut mi	g->1	n->1	
ut mo	t->2	
ut my	c->2	
ut mö	j->1	
ut na	m->1	
ut nr	 ->1	
ut nä	r->1	
ut nå	g->1	
ut nö	d->10	
ut oc	h->10	k->1	
ut om	 ->19	f->1	
ut os	s->1	
ut pe	n->2	
ut pl	ö->1	
ut po	l->1	
ut pr	e->1	o->1	
ut på	 ->22	.->1	m->1	
ut re	g->1	n->1	s->1	
ut se	 ->1	
ut si	g->1	n->1	
ut sk	u->1	
ut so	m->14	
ut st	o->1	ö->1	
ut sy	f->1	
ut sä	g->1	
ut så	 ->2	
ut ta	 ->1	
ut ti	d->1	l->3	
ut un	d->2	
ut up	p->1	
ut ut	a->1	g->1	t->1	
ut va	r->1	
ut vi	d->1	l->1	
ut än	 ->1	
ut är	 ->3	
ut ås	t->1	
ut öv	e->5	
ut, a	l->1	t->3	
ut, b	l->1	
ut, e	f->1	
ut, f	a->1	ö->1	
ut, h	a->2	o->1	u->1	
ut, i	 ->2	
ut, m	e->4	
ut, n	ä->1	
ut, o	c->4	m->1	
ut, s	a->1	o->2	å->1	
ut, t	i->2	
ut, u	t->2	
ut, v	i->1	
ut, å	t->1	
ut. D	e->2	
ut.(P	a->1	
ut.)F	r->1	
ut.De	t->7	
ut.Då	 ->2	
ut.Fi	n->1	
ut.Fr	å->1	
ut.Fö	r->2	
ut.Gr	e->1	
ut.In	t->1	
ut.Ja	g->5	
ut.Kr	a->1	
ut.Na	t->2	
ut.Oc	h->1	
ut.Sk	a->1	
ut.St	ö->1	
ut.Tv	å->1	
ut.Va	d->1	
ut.Vi	 ->1	
ut.Äv	e->1	
ut: f	r->1	
ut; d	e->1	
ut?. 	(->1	
ut?Et	t->1	
uta a	r->1	t->1	
uta d	e->4	
uta e	n->1	t->1	
uta f	ö->2	
uta g	e->1	r->1	
uta i	 ->1	h->1	
uta k	r->1	
uta l	ä->1	
uta m	e->5	i->1	y->1	
uta o	m->11	s->1	
uta p	r->1	
uta r	e->2	
uta s	i->6	o->1	
uta u	n->1	p->5	
uta v	e->1	i->1	
uta Ö	s->2	
uta, 	e->1	h->1	m->1	u->2	
utabe	l->2	
utabl	a->1	
utad,	 ->1	
utad.	(->1	F->1	H->1	O->14	R->1	
utade	 ->6	s->5	
utafr	å->10	
utal.	H->1	
utala	 ->1	
utan 	I->1	a->65	b->6	d->32	e->14	f->7	g->3	h->8	i->6	j->1	k->10	m->8	n->10	o->36	p->9	r->5	s->17	t->34	u->2	v->5	ä->10	ö->3	
utan,	 ->4	
utan.	M->1	
utand	e->27	
utanf	ö->32	
utanv	ä->1	
utapo	l->1	
utar 	A->1	a->2	e->1	m->1	n->1	o->2	
utar.	D->1	
utarb	e->31	
utarm	a->10	
utas 	c->1	f->1	h->1	i->1	m->2	o->1	p->2	u->2	
utasp	e->2	
utat 	a->4	d->2	e->2	o->1	s->1	v->1	
utats	 ->2	.->1	
utaun	i->3	
utbas	u->1	
utbes	t->1	
utbet	a->7	
utbil	d->60	
utbre	d->4	
utbud	 ->3	s->1	
utbyg	g->3	
utbyt	a->1	e->16	
utdel	a->1	
ute e	f->1	
ute p	å->1	
ute t	i->1	
ute u	p->1	
uteau	 ->1	,->2	
utelä	m->3	
uten 	P->1	a->1	d->2	e->1	f->1	i->1	o->2	p->1	s->1	t->2	v->1	ä->1	
uten,	 ->2	
uten.	F->1	J->1	O->1	
utens	 ->1	
uter 	b->1	d->1	f->1	i->2	j->2	m->4	n->1	s->2	t->1	u->1	ö->1	
uter,	 ->1	
uter.	J->4	T->1	V->1	
utera	 ->23	.->3	d->9	r->22	s->10	t->11	
uterr	e->2	
utesl	u->17	ö->2	
utest	ä->4	
utet 	a->28	f->5	h->1	i->1	k->1	m->1	o->6	p->2	s->2	t->1	u->1	v->2	ä->1	
utet,	 ->2	
utet.	F->1	
utet?	Ä->1	
utets	 ->1	
utfal	l->1	
utfas	n->3	
utfla	g->1	
utfly	t->1	
utfor	m->39	s->1	
utfrå	g->7	
utfär	d->12	
utfäs	t->1	
utför	 ->7	a->17	d->3	l->3	s->3	t->13	
utgav	s->1	
utgic	k->1	
utgif	t->14	
utgil	t->8	
utgiv	i->1	n->1	
utgjo	r->4	
utgå 	e->1	f->2	t->1	
utgån	g->16	
utgår	 ->8	
utgåv	o->1	
utgör	 ->45	,->1	.->1	a->10	s->2	
uthan	t->1	
uther	a->1	
uthär	d->4	
utier	 ->1	
utifr	å->16	
utik 	o->1	
utine	n->1	r->6	
utinm	ä->1	
ution	 ->43	,->11	.->13	e->177	s->16	
utiqu	e->1	
utit 	e->1	m->1	s->2	
utits	 ->7	
utjäm	n->5	
utkan	t->1	
utkas	t->15	
utkom	.->1	m->1	s->1	
utkon	k->1	
utkrä	v->3	
utlan	d->5	
utlig	 ->1	a->8	e->63	
utlov	a->3	
utläg	g->1	
utläm	n->2	
utlän	d->3	n->1	
utlåt	a->2	
utlös	a->1	t->1	
utman	a->1	i->19	
utmyn	n->1	
utmär	k->32	
utna 	a->1	d->1	h->1	i->1	m->1	o->2	t->2	v->1	
utna,	 ->3	
utna.	 ->1	D->1	E->1	U->1	
utnin	g->41	
utnyt	t->41	
utnäm	n->4	
uto/O	i->1	
utom 	P->1	a->9	b->8	d->4	e->2	f->5	g->3	h->3	i->2	k->8	m->7	n->2	o->1	p->3	r->3	s->4	t->3	v->5	ä->5	
utom,	 ->2	
utoma	t->8	
utome	u->3	
utomo	r->7	
utoms	t->2	
utopi	l->1	
utor 	t->1	
utpek	a->1	
utper	i->1	
utplå	n->2	
utpre	s->1	
utprä	g->1	
utpun	k->1	
utral	i->1	t->1	
utre 	p->1	
utred	a->3	d->1	n->4	
utres	 ->1	u->3	
utrik	e->19	
utrop	a->2	
utrot	a->2	n->2	
utrou	x->1	
utrus	t->4	
utrym	m->11	
uträt	t->2	
uts k	r->1	
uts s	t->1	
uts u	p->4	
uts-b	e->1	
utsam	 ->2	h->6	t->6	
utsar	 ->1	
utsat	 ->1	s->41	t->8	
utsce	n->1	
utsch	e->1	
utse 	d->1	e->2	m->1	o->2	v->1	
utse.	E->1	
utsed	d->1	
utsee	n->1	
utser	 ->1	
utses	 ->2	.->1	
utset	t->3	
utsfa	t->11	
utsfö	r->1	
utsig	a->1	
utsik	t->1	
utsko	t->157	
utsla	g->15	
utslä	p->9	
utspr	o->4	
utsrä	t->1	
utsta	t->11	
utstr	ä->28	
utstä	l->2	
utstå	t->1	
utstö	t->1	
utsug	a->1	
utsäg	a->1	e->1	
utsät	t->61	
utsåg	s->3	
utta 	r->1	ö->1	
uttal	a->98	
utte 	O->1	
utten	 ->1	
uttig	a->1	
uttit	 ->1	
uttjä	n->24	
uttna	 ->1	.->1	
uttol	k->1	
utton	 ->1	a->1	d->1	
uttor	k->1	
uttry	c->72	
utträ	d->1	
uttöm	d->1	m->3	t->1	
utval	d->1	
utvap	e->1	
utvar	a->2	
utvec	k->237	
utver	k->3	s->1	
utvid	g->106	
utvis	a->1	
utvär	d->32	
utyp,	 ->1	
utänd	a->5	
utåt"	,->1	
utöka	 ->6	d->1	n->1	s->2	t->1	
utökn	i->1	
utöva	 ->7	n->1	r->3	s->4	
utöve	r->14	
utövn	i->1	
uum o	c->1	
uumta	n->1	
uva i	 ->1	
uvara	n->46	
uvele	n->1	r->1	
uverg	n->1	
uvern	ö->1	
uverä	n->17	
uvida	 ->15	
uvriè	r->1	
uvud 	t->9	
uvuda	k->2	n->5	
uvudd	e->3	
uvude	t->1	
uvudf	r->4	ö->1	
uvudl	i->2	
uvudm	å->2	
uvudr	e->1	o->2	
uvuds	a->16	t->4	y->1	
uvudu	p->1	
ux, n	o->1	ä->1	
ux-af	f->1	
uxemb	u->6	
uxhav	e->1	
uxit 	u->1	
uxna 	e->1	
uxna.	H->1	
uyu i	 ->1	
uyu s	a->1	
v "pa	r->1	
v "re	s->1	
v "ri	k->1	
v (KO	M->1	
v - d	e->1	
v - i	n->1	
v - o	c->3	
v - p	å->1	
v - s	a->1	o->1	
v - u	t->1	
v 14 	m->1	
v 19 	d->1	
v 199	9->2	
v 200	0->1	
v 40 	p->1	
v 410	 ->1	
v 5 0	0->1	
v 540	 ->1	
v 8 4	6->1	
v 93/	7->1	
v 94/	5->2	
v 96/	3->3	7->2	
v Ahe	r->2	
v Ame	r->1	
v Ams	t->1	
v Ara	b->1	
v BNI	 ->1	
v BNP	 ->4	,->1	
v BSE	-->1	
v Bar	e->1	n->1	
v Ber	e->2	g->4	n->2	
v Bou	r->1	
v Bro	k->2	
v Can	d->1	
v Da 	C->1	
v Dav	i->1	
v Dem	i->1	
v Dim	i->2	
v Dub	l->1	
v Düh	r->1	
v EG-	d->1	
v EU 	a->1	o->1	s->1	
v EU,	 ->1	
v EU-	b->1	g->1	k->1	l->1	
v EU.	D->1	V->1	
v EU:	s->7	
v Enl	i->1	
v Eri	k->1	
v Eur	o->70	
v Exx	o->2	
v FN:	s->1	
v FPÖ	 ->1	:->1	
v Flo	r->1	
v För	e->7	i->1	
v Gaz	a->1	
v Gen	e->2	
v Gra	c->1	ç->1	
v Gro	s->1	
v Hai	d->1	
v Hen	r->1	
v Hit	l->1	
v Isr	a->2	
v Jac	o->1	
v Jer	u->1	
v Jon	c->2	
v Kin	n->3	
v Koc	h->3	
v Kos	o->7	
v Kul	t->1	
v Lan	g->3	
v Lib	a->1	
v Löö	w->1	
v Mar	i->2	
v McN	a->1	
v Mor	g->1	
v OLA	F->3	
v Osm	a->1	
v Oz 	d->1	
v Pal	a->1	
v Pat	t->1	
v Por	t->1	
v Pét	a->1	
v Rap	k->1	
v Rii	s->1	
v Sam	m->1	
v Sch	e->3	r->3	
v Tac	i->1	
v Ter	r->1	
v The	a->3	
v Thy	s->1	
v Tib	e->1	
v Tot	a->1	
v UNM	I->1	
v Van	 ->1	
v Var	e->1	
v Väs	t->1	
v Wal	e->1	
v Wie	l->1	
v Wye	-->1	
v acc	e->1	
v adm	i->1	
v adv	o->1	
v age	r->1	
v alb	a->1	
v ald	r->1	
v alk	o->1	
v all	 ->2	a->12	e->1	m->4	t->11	v->3	
v anb	u->1	
v and	a->2	r->3	
v anl	e->1	ä->1	
v anm	ä->1	
v ano	n->1	
v ans	e->1	j->1	k->1	l->1	t->1	v->11	
v ant	a->3	
v anv	ä->2	
v apr	i->2	
v arb	e->20	
v art	e->1	i->19	
v asy	l->1	
v att	 ->69	i->1	
v av 	"->1	a->2	d->1	e->4	f->1	p->1	s->3	v->1	ö->1	
v av,	 ->1	
v av.	O->1	
v avf	a->1	
v avg	ö->4	
v avp	r->1	
v avs	l->1	p->1	
v avt	a->2	
v avv	e->2	
v bar	b->1	n->1	
v bas	e->1	
v bed	r->1	
v bef	i->2	o->4	
v beg	r->1	
v beh	a->2	o->1	ö->3	
v bek	v->1	
v bes	l->9	t->6	ö->1	
v bet	r->1	y->2	ä->6	
v bev	i->2	
v bid	r->3	
v bil	a->4	d->1	e->1	i->1	t->1	v->3	
v bio	p->1	
v bla	n->2	
v bly	 ->1	
v blå	 ->1	
v bol	a->1	
v bom	b->1	u->1	
v bre	v->1	
v bri	s->4	
v bro	t->4	
v bru	t->1	
v bud	g->8	
v byg	g->2	
v båd	e->2	
v böc	k->1	
v bör	d->2	
v cen	t->2	
v cir	k->2	
v civ	i->4	
v com	m->1	
v dag	.->1	e->3	o->1	
v dat	a->1	
v de 	C->2	a->7	b->9	d->1	e->11	f->27	g->5	h->4	i->6	k->2	l->2	m->15	n->13	o->4	p->11	r->7	s->19	t->7	u->1	v->6	ä->1	å->4	ö->1	
v deb	a->3	
v def	i->1	
v del	a->2	t->1	
v dem	 ->16	,->1	.->5	:->1	o->4	
v den	 ->149	,->1	.->1	n->32	
v der	a->6	
v des	s->45	
v det	 ->83	,->2	.->2	t->41	
v dip	l->1	
v dir	e->21	
v dis	c->1	k->5	
v div	e->1	
v dju	n->1	p->1	
v dok	u->1	
v dom	a->5	i->1	s->5	
v dri	v->1	
v där	 ->1	f->1	
v eff	e->2	
v eft	e->3	
v ege	n->2	
v eko	l->2	n->10	
v en 	a->8	b->4	d->4	e->5	f->4	g->2	h->2	i->1	k->5	l->2	m->10	n->2	o->5	p->12	r->10	s->14	t->3	u->3	å->1	ö->2	
v enb	a->1	
v ene	r->9	
v enh	e->1	
v eni	g->1	
v eno	r->1	
v ent	r->2	
v er 	a->1	b->1	h->2	k->1	s->2	t->1	u->1	
v er,	 ->2	
v er:	 ->1	
v era	 ->3	
v erf	a->1	
v ert	 ->2	
v etn	i->1	
v ett	 ->51	
v eur	o->7	
v eve	n->1	
v exa	k->1	m->5	
v exp	e->1	
v ext	e->1	
v fak	t->3	
v fal	l->2	s->1	
v far	l->31	t->8	
v fat	t->4	
v fin	a->3	
v fis	k->3	
v fjo	r->2	
v fle	r->7	x->2	
v flo	t->1	
v fly	k->6	
v fol	k->1	
v fon	d->1	
v for	d->4	s->2	
v fra	m->1	
v fre	d->1	
v fri	a->3	h->6	s->1	v->1	
v frä	m->5	
v frå	g->7	n->11	
v ful	l->2	
v fun	g->1	
v fus	i->2	
v fys	i->1	
v fäd	e->1	
v få 	i->1	
v fån	g->1	
v får	 ->3	
v föl	j->2	
v för	 ->13	a->1	d->12	e->28	f->1	h->7	l->3	n->13	o->2	r->5	s->24	t->3	u->4	v->4	ä->2	å->1	
v gam	l->3	
v gem	e->28	
v gen	e->2	o->1	
v geo	g->1	
v gif	t->1	
v gig	a->1	
v giv	a->1	
v glo	b->1	
v god	a->1	k->1	
v gra	d->1	n->1	
v gro	v->1	
v gru	n->3	
v grä	n->4	
v grö	n->1	
v gör	 ->1	
v ha 	b->1	
v han	 ->1	d->3	s->1	
v har	 ->7	m->1	
v hat	 ->1	i->1	
v hav	e->3	s->1	
v hel	a->6	
v hem	l->1	
v hie	r->1	
v hig	h->1	
v his	t->3	
v hjä	l->1	
v hon	o->1	
v hun	d->1	
v hur	 ->5	u->2	
v hän	v->1	
v här	.->1	
v hög	 ->1	s->1	
v hör	 ->1	
v i K	o->1	
v i d	a->1	e->7	
v i e	g->1	
v i s	a->1	n->1	v->1	y->1	
v i v	i->1	
v ibe	r->1	
v ick	e->3	
v ide	a->1	
v idé	e->1	
v imp	o->4	u->1	
v in 	i->1	
v ind	u->1	
v ine	f->1	
v inf	o->3	r->1	
v ini	t->2	
v inn	e->2	o->1	
v ino	m->2	
v inr	e->2	
v ins	t->4	y->1	
v int	e->10	o->1	r->2	
v inv	a->2	e->1	
v jor	d->5	
v jur	i->1	
v jus	t->3	
v jäm	s->2	
v kam	m->2	
v kan	 ->1	a->2	d->1	
v kap	i->1	
v kar	a->1	t->2	
v kat	a->3	
v kla	r->2	s->2	
v knu	t->1	
v koa	l->2	
v kol	d->3	l->1	
v kom	m->61	
v kon	c->2	f->4	k->31	s->2	t->4	
v kor	t->2	
v kos	t->7	
v kri	g->1	m->1	s->1	t->1	
v krä	n->1	
v kul	t->4	
v kus	t->1	
v kva	l->1	r->1	
v kvi	n->4	
v kvo	t->1	
v kär	n->8	
v lag	 ->1	.->1	s->10	
v lan	d->8	
v las	t->1	
v led	a->8	e->1	n->1	
v leg	i->1	
v lej	d->1	
v lib	e->2	
v lic	e->1	
v lik	n->2	
v lis	t->3	
v liv	 ->1	s->7	
v loj	a->2	
v lok	a->3	
v läg	e->1	
v läm	n->1	
v län	d->1	g->1	
v lät	t->1	
v lån	g->1	
v lös	n->1	
v löv	s->1	
v mak	t->2	
v man	 ->1	d->1	
v mar	g->1	k->6	s->3	
v mat	e->4	
v med	 ->8	b->5	e->2	l->12	
v men	i->1	
v mer	 ->1	i->1	v->1	
v mig	 ->2	
v mil	j->14	
v min	 ->7	a->7	d->2	o->1	s->1	
v mis	s->3	
v mit	t->3	
v mod	e->2	
v mon	o->1	
v mot	 ->1	i->1	s->1	
v myc	k->3	
v män	n->7	
v mål	 ->2	s->1	
v mån	g->4	
v mås	t->1	
v möj	l->1	
v nat	i->9	u->4	
v naz	i->1	
v ni 	l->1	
v nor	d->1	
v ny 	i->1	v->1	
v nya	 ->6	
v nyb	i->1	
v nyh	e->1	
v nyl	i->1	
v nyn	a->1	
v nys	s->1	
v när	 ->1	
v näs	t->1	
v någ	o->6	
v nöd	v->2	
v oac	c->1	
v oan	s->1	
v oav	s->1	
v obe	r->2	s->1	
v obl	i->1	
v och	 ->25	
v ock	s->4	
v off	e->3	r->1	
v ofr	e->1	
v okl	a->1	
v oli	k->8	
v olj	a->1	e->2	
v oly	c->3	
v om 	a->1	d->1	e->2	f->2	g->1	h->3	l->2	s->3	t->2	u->5	v->2	ä->1	
v omb	u->1	
v ome	d->1	
v omf	å->1	
v omk	r->1	
v omr	ö->2	
v oms	t->2	
v ond	o->1	
v opi	n->1	
v ord	a->1	f->6	
v ori	k->1	
v ork	a->1	
v ors	a->2	
v oss	 ->10	,->1	.->1	
v otr	y->1	
v otv	e->1	
v oun	d->1	
v ova	n->1	
v pak	t->1	
v pal	e->1	
v par	l->18	t->2	
v pen	g->6	n->1	
v per	s->5	
v pio	n->1	
v pol	i->9	
v pre	s->1	
v pri	n->4	o->2	s->2	
v pro	b->3	c->1	d->4	g->11	j->4	t->5	
v på 	8->1	a->4	b->3	d->7	e->5	f->1	h->1	i->2	m->2	n->1	r->1	s->3	
v påv	e->2	
v ram	a->2	
v rap	p->3	
v ras	i->1	
v ref	o->3	
v reg	e->9	i->4	l->4	
v rek	o->1	
v ren	 ->1	
v rep	u->1	
v res	o->2	p->2	u->4	
v ret	r->1	
v rev	i->1	
v rik	t->5	
v ris	k->3	
v rol	l->2	
v rys	k->1	
v räd	s->1	
v räk	e->4	n->1	
v rät	t->6	
v råd	e->12	
v rös	t->1	
v sak	 ->1	
v sam	a->2	f->2	h->3	m->5	o->1	t->1	v->1	
v sce	n->1	
v se 	t->1	
v sed	a->1	
v seg	e->1	
v sek	r->1	t->1	
v sen	a->1	
v ser	b->1	
v ses	s->2	
v sex	u->1	
v sid	a->1	
v sig	 ->3	
v sin	 ->3	a->10	
v sis	t->1	
v sit	t->2	u->5	
v sju	k->1	
v sjä	l->1	
v sjö	v->1	
v ska	d->1	l->4	n->1	p->1	t->3	
v ske	p->1	
v sko	g->4	
v skr	o->3	
v sku	l->1	
v skä	l->3	
v skö	r->1	
v slu	t->2	
v små	 ->2	
v sna	b->1	
v soc	i->7	
v sol	i->1	
v som	 ->37	m->1	
v spe	c->1	
v spl	i->1	
v sta	b->5	r->1	t->18	
v sti	c->1	m->1	
v sto	r->14	
v str	a->3	u->13	
v sty	r->1	
v stä	d->1	
v stå	l->2	n->1	
v stö	d->11	r->8	t->1	
v sub	s->3	
v suc	c->1	
v sva	r->1	
v svä	l->1	
v syf	t->2	
v syn	s->1	
v sys	s->16	t->5	
v säg	e->1	
v säk	e->9	
v sär	s->5	
v så 	a->2	s->3	u->1	
v såd	a->8	
v sås	o->1	
v ta 	a->1	
v tal	a->1	m->1	r->1	
v tek	n->4	
v tel	e->1	
v ter	r->3	
v tid	i->1	s->1	
v til	l->36	
v tim	m->2	
v tjä	n->28	
v tot	a->2	
v tra	d->2	n->5	
v tre	 ->2	d->1	
v try	c->1	
v trä	 ->1	d->1	
v tun	g->4	n->1	
v tur	i->1	
v tvu	n->1	
v två	 ->1	
v tyd	l->1	
v typ	 ->1	
v tän	k->1	
v und	a->3	e->5	
v ung	a->2	
v uni	o->20	
v upp	 ->1	g->2	m->3	
v uta	n->1	r->5	
v utb	i->2	
v utf	a->1	ä->1	
v utg	i->3	
v utn	y->1	
v utr	i->1	u->1	
v uts	k->7	
v utt	j->3	
v utv	e->6	i->5	
v vad	 ->11	?->1	
v van	 ->3	
v vap	e->1	
v var	f->1	i->1	j->4	
v vat	t->1	
v ved	e->1	
v ver	k->2	t->1	
v vet	 ->1	e->5	
v vi 	h->1	
v vic	e->4	
v vid	 ->1	
v vik	t->3	
v vil	k->5	l->2	
v vis	s->9	
v vit	b->1	
v von	 ->4	
v väg	a->1	
v väl	 ->1	f->1	j->1	
v vän	d->1	s->1	
v vär	d->3	l->4	s->1	
v väx	e->1	t->5	
v vår	 ->4	a->15	d->1	t->4	
v ytt	e->4	r->1	
v Öst	e->2	
v äld	r->1	
v ämn	e->1	
v än 	d->1	
v änd	r->4	
v änn	u->1	
v är 	a->1	d->3	f->1	g->1	n->1	s->1	v->1	
v åld	e->1	
v år 	2->5	e->1	
v åre	t->1	
v årh	u->1	
v åsi	k->1	
v åte	r->4	
v åtg	ä->12	
v öbo	 ->1	
v öde	m->1	
v öka	d->3	r->1	
v öpp	e->4	
v öst	e->2	
v öve	r->4	
v", d	ä->1	
v, 95	/->1	
v, an	v->1	
v, at	t->2	
v, ba	r->1	
v, de	 ->1	l->1	t->1	
v, dv	s->1	
v, dä	r->1	
v, ef	t->1	
v, en	 ->1	k->1	
v, fr	a->1	
v, ha	r->1	
v, he	r->2	
v, hy	s->1	
v, in	t->1	
v, ja	g->1	
v, li	k->1	
v, me	n->4	
v, mi	n->1	
v, nä	m->1	
v, nå	g->1	
v, oc	h->7	
v, om	 ->1	
v, so	m->4	
v, st	ö->1	
v, sä	r->1	
v, så	 ->2	
v, ti	l->1	
v, tr	o->1	
v, un	d->1	
v, är	 ->2	
v. De	 ->1	
v. Me	n->1	
v. Va	r->1	
v. Vi	 ->1	
v. me	n->1	
v."De	t->1	
v.(Sa	m->1	
v., ä	v->1	
v.. (	E->2	
v..He	r->1	
v.?An	s->1	
v.Att	 ->1	
v.Av 	d->1	
v.Avs	l->1	
v.Bar	a->1	
v.Bla	n->1	
v.De 	1->1	n->1	p->1	
v.Den	 ->1	
v.Det	 ->5	t->2	
v.Där	f->1	
v.Då 	s->1	
v.Eff	e->1	
v.En 	a->1	v->1	
v.Eri	k->1	
v.Fru	 ->1	
v.För	 ->4	
v.Her	r->1	
v.I d	a->1	
v.I v	a->1	
v.Ing	e->1	
v.Jag	 ->2	
v.Kom	m->1	
v.Låt	 ->1	
v.Men	 ->3	
v.OLA	F->1	
v.Om 	e->1	
v.Rik	t->1	
v.Råd	e->1	
v.Sve	p->1	
v.Sås	o->1	
v.Upp	r->1	
v.Vi 	d->1	ä->1	
v.Vis	s->1	
v.Ytt	e->1	
v: Fö	r->1	
v: vå	g->1	
v; an	t->1	
v?För	 ->1	
v?Nej	,->1	
v?Vil	k->1	
va 40	 ->1	
va Eu	r->2	
va an	s->4	t->1	
va ar	b->1	
va at	t->7	
va av	 ->1	s->3	t->1	
va ba	s->1	
va be	f->1	s->2	t->2	
va bi	e->2	l->1	
va bj	u->1	
va bo	r->2	
va br	i->1	
va bä	r->1	
va ce	n->1	
va da	g->1	
va de	 ->1	b->1	m->6	n->3	s->1	t->6	
va dr	a->1	
va du	b->2	
va dä	r->1	
va ef	f->4	t->3	
va en	 ->16	e->1	
va et	t->2	
va eu	r->1	
va ex	a->1	
va fa	k->1	n->1	t->1	
va fi	n->1	
va fl	e->1	
va fu	n->1	
va fö	l->3	r->7	
va ga	m->1	
va gä	c->1	
va gö	r->3	
va ha	n->1	r->2	
va hu	r->2	
va hö	g->1	
va i 	K->1	S->1	d->1	f->1	h->1	k->1	m->1	s->2	
va id	é->1	
va ig	e->1	
va im	p->1	
va in	d->1	f->1	s->1	
va ju	r->1	
va ka	n->1	p->2	r->1	
va kl	a->2	
va ko	m->3	n->3	s->1	
va kr	a->1	i->2	
va ku	n->1	
va kä	n->1	r->3	
va la	g->1	
va le	v->1	
va li	k->1	s->1	
va lö	s->1	
va me	d->3	r->1	
va mi	n->1	
va mo	t->1	
va må	l->1	s->1	
va ni	v->1	
va nå	g->4	
va oc	h->13	
va of	f->1	
va om	 ->1	
va or	d->2	g->1	
va pa	r->2	
va po	l->4	
va pr	i->1	o->1	
va pu	n->1	
va på	 ->4	m->1	t->1	
va ra	m->1	
va re	a->1	f->2	g->2	s->1	
va ri	k->1	
va ro	l->1	
va ru	t->1	
va rä	t->1	
va rå	d->1	
va sa	m->3	
va se	k->1	
va si	d->1	n->2	
va sj	ä->1	
va sk	a->1	r->1	
va sl	u->1	
va so	m->2	
va st	a->1	o->1	å->1	
va sv	å->1	
va sy	f->1	n->1	s->1	
va te	a->1	n->1	
va ti	d->3	l->11	
va tr	a->1	
va tv	å->1	
va un	i->1	
va up	p->2	
va ur	s->1	
va ut	 ->1	t->1	v->1	
va ve	r->29	
va vä	g->2	
va vå	r->2	
va är	 ->2	
va år	 ->1	,->1	
va ås	i->1	
va åt	g->5	
va ök	a->2	
va öv	e->1	
va, d	å->1	
va, f	ö->1	
va, i	n->1	
va, s	k->1	å->2	
va, u	t->2	
va, ä	r->1	
va.Al	l->1	
va.De	t->1	
va.He	r->1	
va.Lå	t->1	
va.Nä	r->1	
va.Om	 ->1	
va.Va	d->1	
va.Vå	r->1	
va?Ne	j->1	
vacke	r->2	
vackl	a->1	
vackr	a->6	
vad B	N->1	
vad E	u->1	
vad G	u->1	
vad K	u->2	
vad S	y->1	
vad a	l->1	
vad b	e->14	
vad d	a->1	e->28	o->1	
vad e	n->2	t->1	
vad f	ö->3	
vad g	e->1	r->1	ä->45	
vad h	a->3	ä->1	
vad i	d->1	
vad j	a->7	
vad k	a->1	o->7	
vad m	a->8	e->1	
vad n	a->1	i->4	
vad o	c->1	m->1	r->1	
vad p	r->1	
vad r	i->1	å->1	
vad s	o->55	t->3	y->2	
vad t	j->1	
vad v	a->1	e->4	i->18	o->1	å->3	
vad ä	r->5	v->1	
vad?D	ä->1	
vade 	i->2	j->1	m->3	p->1	s->2	
vade.	S->1	
vades	 ->2	
vag i	n->1	
vag p	o->1	
vag s	t->1	
vaga 	H->1	d->4	j->1	o->1	r->2	s->1	
vaga,	 ->2	
vagad	e->3	
vagar	 ->4	e->2	
vagas	 ->3	,->1	.->1	t->2	
vagat	s->2	
vaghe	t->12	
vagne	n->2	
vagni	n->1	
vagt.	J->1	
vaka 	-->1	E->1	d->1	f->1	g->1	i->1	o->2	v->1	ö->1	
vaka.	L->1	
vakar	 ->4	e->1	
vakas	 ->2	
vakat	 ->1	
vakie	n->1	
vakni	n->14	
vaksa	m->9	
vakt 	o->1	
vakta	n->4	r->2	
vakte	r->1	
vakuu	m->2	
val a	t->1	v->21	
val d	e->1	
val e	n->1	
val f	ö->1	
val g	ö->1	
val i	 ->1	n->1	
val l	ä->1	
val m	ö->1	
val s	k->1	o->1	
val u	n->1	
val ä	n->1	
val å	t->1	
val, 	o->3	
val.D	e->1	
val.I	n->1	
val.M	e->1	
val.S	t->1	
val.V	i->1	
val; 	a->1	
valar	 ->1	.->2	
valba	r->1	
vald 	f->4	k->1	p->2	r->1	
vald.	J->1	
valda	 ->13	,->1	?->1	g->1	
valde	 ->2	l->3	s->3	
valdi	s->1	
valen	 ->5	,->1	
vales	e->1	
valet	 ->6	
valfr	a->3	i->2	
valif	i->15	
valit	a->6	e->30	
valkr	e->4	
vallf	ä->1	
vallp	o->1	
valre	s->1	
valsk	o->1	
valt 	a->3	d->1	u->1	
valt,	 ->1	
valta	 ->1	k->1	r->1	
valti	d->1	
valtn	i->47	
valts	 ->3	.->1	
valut	a->23	
van D	a->2	
van G	o->1	
van H	u->20	
van V	e->1	
van a	t->3	
van d	e->9	
van e	f->3	
van m	o->1	
van o	c->1	
van, 	f->1	
van.D	å->1	
van.T	y->1	
vana 	a->1	v->1	
vance	r->1	
vanda	n->1	
vande	 ->21	,->1	.->2	;->1	n->7	t->4	
vandl	a->7	i->2	
vandr	a->11	i->7	
vanhe	d->2	
vanif	r->1	
vanli	g->12	
vannä	m->2	
vanor	.->1	
vanos	 ->1	!->1	
vanpå	 ->1	
vans 	a->1	f->2	l->1	
vans,	 ->4	
vanse	n->1	
vansi	n->1	
vansk	a->2	l->1	
vanst	å->1	
vansv	ä->1	
vant 	f->2	g->1	s->1	
vanta	 ->6	
vanti	f->4	t->4	
vapen	 ->13	,->3	.->4	?->1	h->1	i->1	s->1	t->1	u->1	
vapne	n->2	
var -	 ->2	
var 1	,->1	5->1	9->3	
var 9	7->1	
var K	u->1	
var W	a->1	
var a	k->1	l->2	n->1	t->15	v->6	
var b	a->3	e->2	l->3	r->3	ä->1	å->1	ö->1	
var d	a->1	e->30	o->1	ä->4	å->1	
var e	f->5	l->1	m->1	n->18	r->1	t->8	x->2	
var f	a->2	l->1	r->2	ö->35	
var g	e->3	i->1	ä->1	
var h	a->1	e->2	o->3	ä->1	ö->1	
var i	 ->11	n->15	
var j	a->4	
var k	a->2	l->1	o->2	v->1	
var l	i->2	y->1	ä->2	ö->1	
var m	a->2	e->7	y->6	å->2	ö->1	
var n	a->2	e->1	i->2	ä->3	å->1	ö->2	
var o	a->1	c->11	e->1	k->1	s->1	
var p	r->1	å->24	
var r	e->1	i->1	ä->2	å->1	
var s	a->1	e->1	i->2	j->2	o->11	t->2	ä->2	å->6	
var t	a->1	i->1	u->1	v->4	y->1	
var u	p->2	t->1	
var v	e->1	i->7	ä->3	
var ä	n->2	r->5	
var ö	v->4	
var, 	a->2	d->3	f->3	h->1	i->1	k->1	l->3	m->1	o->9	s->2	v->2	ä->1	å->1	
var. 	M->1	
var.D	e->14	
var.E	r->1	
var.F	ö->1	
var.G	e->2	ö->1	
var.I	 ->2	
var.J	a->5	
var.M	e->4	
var.N	å->1	
var.O	m->1	
var.P	å->1	
var.R	e->1	
var.S	e->2	o->1	
var.V	i->5	
var; 	o->1	
var?I	 ->1	
vara 	"->1	1->1	B->1	E->2	a->21	b->14	c->2	d->23	e->59	f->33	g->7	h->9	i->11	j->2	k->17	l->12	m->42	n->18	o->13	p->8	r->8	s->34	t->19	u->8	v->14	y->1	ä->3	ö->5	
vara"	.->1	
vara,	 ->2	
vara.	D->1	J->2	M->1	
vara:	 ->1	
varad	 ->1	e->10	
varak	t->4	
varan	.->1	d->120	n->1	
varar	 ->32	,->1	e->2	
varas	 ->2	
varat	 ->3	s->3	
varav	 ->4	
varda	g->4	
varde	r->1	
vare 	a->2	d->3	e->1	f->8	h->1	i->2	k->4	l->1	m->1	o->2	p->2	r->1	s->17	t->1	ä->2	
vare"	 ->1	,->1	
vare,	 ->5	
vare.	D->2	U->1	V->2	Ä->2	
varef	t->1	
varen	 ->5	,->2	d->2	s->2	
vares	 ->1	
varet	 ->54	,->2	.->16	
varfö	r->39	
varga	r->1	
varhä	n->1	
varhå	l->2	
vari 	e->1	
varie	r->2	
varig	 ->18	,->3	a->29	e->1	h->5	t->6	
varit	 ->71	
varje	 ->84	
varke	n->14	
varko	n->1	
varli	g->62	
varlä	n->1	
varma	 ->3	
varmt	 ->12	
varna	 ->9	"->1	,->4	.->2	d->1	g->1	r->3	s->2	
varni	n->7	
varo 	-->1	i->1	n->1	v->1	
varo,	 ->1	
varon	 ->2	,->1	
varor	,->1	.->1	
varpa	r->1	
varr 	i->1	
vars 	a->1	b->2	e->2	f->5	g->2	h->2	l->1	m->1	n->2	p->1	r->2	s->2	t->1	u->2	ä->1	å->1	
vars.	D->1	
varsa	m->1	v->1	
varsb	e->2	u->1	
varsf	r->47	u->4	ö->4	
varsk	u->1	ä->3	
varsl	a->1	
varsm	a->1	e->1	i->1	
varso	m->6	r->1	
varsp	o->5	
varst	a->2	i->1	å->7	
vart 	d->1	i->1	o->1	r->1	
varta	 ->2	n->3	
varte	n->1	
varv,	 ->1	
varve	n->1	
varvi	d->3	
varvs	i->1	s->2	
vas a	n->1	t->1	v->6	
vas e	n->1	t->2	
vas f	ö->1	
vas h	a->1	
vas i	 ->3	
vas m	e->2	
vas o	c->3	m->1	
vas s	ä->1	
vas, 	s->1	v->1	
vas.C	e->1	
vas.G	e->1	
vas.H	e->1	
vas.I	 ->1	
vas.M	i->1	
vas.V	i->1	
vaste	 ->1	
vat -	 ->1	
vat E	u->1	
vat a	t->2	
vat b	e->1	
vat d	e->1	i->1	
vat e	f->1	
vat f	i->1	
vat o	c->1	
vat r	ä->1	
vat t	r->1	
vat u	t->1	
vat.J	a->1	
vat.Å	 ->1	
vata 	a->1	f->5	i->1	k->1	m->1	o->4	s->4	å->1	
vatek	o->1	
vatio	n->8	
vatis	e->2	
vativ	 ->1	a->8	
vats 	b->1	i->2	p->1	
vats,	 ->1	
vats.	Ä->1	
vatte	n->33	
vattn	a->6	e->8	i->2	
vatör	e->1	
vavta	l->7	
vbest	ä->3	
vbetä	n->1	
vbiog	r->1	
vbord	s->1	
vbrin	g->1	
vbrot	t->4	
vbrut	e->2	
vbryt	e->3	
vbröt	 ->4	s->2	
vbära	n->1	
vda a	t->6	
vda d	e->1	
vdade	 ->3	
vdar 	a->7	b->1	d->1	i->1	
vdar,	 ->1	
vdar.	J->1	
vdat 	a->2	b->1	d->1	
vdat.	T->1	
vde d	e->1	
vde e	n->1	
vde f	a->1	
vde g	o->1	ö->1	
vde, 	f->1	
vdeln	i->8	
vdes 	e->2	
vdvun	n->1	
ve (C	5->2	
ve 19	5->1	
ve Eu	r->1	
ve al	l->1	
ve an	s->1	
ve be	f->2	s->1	
ve bu	d->1	
ve de	n->4	
ve en	e->1	
ve et	t->2	
ve fo	l->1	
ve ka	n->1	
ve ko	m->2	n->1	
ve la	g->1	n->1	
ve my	n->2	
ve må	s->1	
ve pa	r->3	
ve re	a->1	
ve ru	l->1	
ve rä	t->1	
ve sj	u->1	
ve ti	d->1	
ve tr	e->1	
ve är	 ->1	
ve, a	t->1	
ve, å	t->1	
ve- p	r->1	
ve-pr	o->2	
veNäs	t->1	
vebrö	d->1	
vec l	'->1	
vecka	 ->6	.->1	n->17	
veckl	a->73	i->175	
vecko	r->17	
veder	b->11	g->1	t->1	
vek h	o->1	
vek o	s->1	
veka 	a->1	f->1	r->1	
vekad	e->1	
vekan	 ->14	,->1	
vekar	 ->3	
vekat	 ->2	
vekhe	t->4	
veklö	s->1	
vekon	v->1	
veksa	m->5	
vel a	l->1	n->1	t->5	
vel g	a->1	e->1	ö->1	
vel l	e->1	
vel n	y->1	
vel o	m->6	
vel p	å->1	
vel s	t->1	
vel t	i->2	
vel u	n->1	
vel v	a->1	
vel ä	r->1	v->1	
vel, 	a->1	j->1	
velak	t->3	
velat	 ->7	
velen	"->1	
veler	.->1	
velse	 ->5	r->1	
velsu	t->3	
vem b	e->1	
vem f	a->1	
vem i	 ->1	
vem s	k->2	o->10	t->1	
vem ä	r->1	
vembe	r->11	
vems 	a->1	
ven -	 ->1	
ven 7	9->1	
ven E	U->2	u->2	
ven G	r->1	
ven R	a->1	e->1	
ven a	c->1	n->4	r->2	t->5	v->5	
ven b	e->1	r->1	y->1	ö->1	
ven d	e->18	o->1	ä->3	
ven e	f->1	k->1	l->1	n->6	t->2	v->1	
ven f	a->1	i->3	r->7	å->1	ö->17	
ven g	e->2	
ven h	e->1	ä->5	ö->1	
ven i	 ->42	h->1	n->8	
ven j	a->13	
ven k	a->1	o->6	r->2	u->2	
ven l	o->1	ä->3	
ven m	e->11	i->4	y->1	å->3	
ven n	i->1	ä->6	å->1	ö->1	
ven o	c->7	m->80	s->1	
ven p	a->2	r->1	å->14	
ven r	e->2	å->1	
ven s	k->6	m->1	o->2	p->1	t->2	
ven t	a->4	i->5	r->1	v->1	ä->1	
ven u	n->3	p->2	t->2	
ven v	a->2	i->3	ä->1	
ven y	t->1	
ven ä	g->1	n->2	r->2	
ven ö	p->1	v->2	
ven, 	A->1	C->1	n->1	s->1	
ven.D	e->2	
ven.K	r->1	
ven.N	ä->1	
ven.S	a->1	ä->1	
ven.T	o->2	
ven.V	i->1	
ven: 	i->1	
venem	a->1	
vener	a->2	
venhe	t->4	
vens 	a->3	e->1	m->1	
vens.	D->1	
vense	n->3	r->38	
vensk	 ->1	a->2	
vent 	b->2	g->1	o->3	r->1	s->2	u->1	
vent,	 ->2	
venta	 ->4	r->1	
vente	r->1	
venti	l->2	o->40	
ventu	e->21	
venty	r->9	
vep a	t->1	
vepes	k->1	
vepsk	ä->1	
vepte	 ->1	
ver -	 ->2	
ver 1	0->1	
ver 2	0->1	
ver 3	2->1	5->1	
ver 4	 ->1	
ver 5	 ->1	
ver 7	 ->1	
ver 8	0->2	
ver 9	0->1	
ver B	N->1	
ver E	U->1	u->4	
ver H	i->1	
ver O	r->1	
ver a	l->3	n->2	r->2	t->42	v->9	
ver b	e->3	
ver d	a->1	e->46	ä->1	
ver e	k->1	l->1	n->25	t->13	
ver f	r->3	å->1	ö->10	
ver g	a->1	e->2	o->1	r->7	ö->3	
ver h	a->7	e->12	o->1	u->17	ä->1	
ver i	 ->5	n->6	
ver j	a->3	u->1	ä->1	
ver k	a->1	l->1	n->1	o->6	u->1	
ver l	i->1	u->1	ä->1	å->1	
ver m	a->3	e->4	i->3	o->1	y->1	å->2	ö->1	
ver n	a->2	i->1	u->1	y->2	å->3	
ver o	b->1	c->7	m->1	r->3	
ver p	a->1	e->1	r->1	å->4	
ver r	e->6	i->1	ä->1	å->1	
ver s	a->1	e->1	i->4	j->1	k->2	o->2	p->1	t->9	y->1	
ver t	i->4	r->2	v->1	
ver u	n->7	p->1	t->3	
ver v	a->4	e->3	i->22	ä->1	å->2	
ver y	t->1	
ver Ö	s->1	
ver ä	n->1	r->3	
ver å	t->1	
ver, 	k->2	m->1	o->1	s->2	ä->2	
ver. 	F->1	
ver.D	e->2	
ver.H	e->1	
ver.J	a->1	
ver.K	o->2	
ver.M	a->1	
ver.O	r->1	
ver.S	a->1	o->1	
ver.T	i->1	
ver.V	a->1	i->1	
vera 	d->3	f->1	s->1	t->1	
verad	e->10	
veral	l->9	
veran	d->4	t->3	
verar	 ->7	
veras	,->1	.->1	
verat	 ->1	s->1	
verba	l->1	
verbe	l->3	m->1	
verbl	i->1	
verbr	i->1	y->3	
verce	n->1	
verdr	i->14	
veren	s->71	
verer	a->5	
veret	,->1	
verfa	l->3	
verfi	s->1	
verfl	y->2	ö->1	
verfö	l->2	r->14	
verge	 ->2	n->4	r->7	s->2	
vergi	v->2	
vergn	e->1	
vergr	i->14	
vergå	 ->1	n->11	r->3	
verha	n->1	
verhe	a->1	
verhä	n->1	
verhö	g->2	
veri 	-->1	i->1	ä->2	ö->1	
veri,	 ->1	
verie	r->1	t->1	
verif	i->1	
verig	e->7	
verin	g->6	s->1	
verk 	-->1	a->1	b->1	f->3	g->1	i->8	k->1	m->2	o->1	p->1	s->4	u->1	ä->2	
verk,	 ->3	
verk.	B->1	D->1	S->1	V->1	
verk?	R->1	
verka	 ->40	,->1	d->2	n->21	r->121	s->9	t->9	
verke	n->6	t->40	
verkl	a->6	i->205	
verkn	i->15	
verks	a->51	t->19	
verkt	y->8	
verla	g->1	
verle	v->5	
verlä	g->6	m->15	
verlå	t->8	
vermo	d->1	r->1	
verna	t->3	
verni	t->1	
vernö	r->1	
veror	d->1	
verpr	i->1	
verra	s->1	
verre	g->2	
verrö	s->1	
vers,	 ->1	
versa	l->1	t->1	
verse	 ->2	l->3	n->1	r->1	
versi	e->2	f->2	k->18	o->13	
versk	r->17	å->6	
verst	a->4	i->5	
versv	ä->7	
versy	n->1	
versä	t->11	
verta	 ->1	g->3	l->1	r->1	
verti	k->3	
verto	g->1	n->1	
vertr	a->1	ä->6	
verty	g->38	
vertä	n->1	
verva	k->25	
vervi	n->8	
vervu	n->1	
vervä	g->35	l->3	
very,	 ->1	
verän	 ->2	a->3	i->12	
ves h	a->1	
ves o	c->1	
veste	r->15	
vesto	r->3	
vet "	O->1	
vet -	 ->2	
vet E	q->8	
vet L	e->1	
vet S	j->1	
vet a	l->4	t->50	v->23	
vet b	e->1	y->1	ä->1	
vet f	r->5	ö->7	
vet g	e->3	ä->1	ö->1	
vet h	a->7	e->1	o->1	u->1	ö->1	
vet i	 ->4	g->1	n->14	
vet j	a->3	
vet k	a->1	o->2	v->1	
vet m	e->3	y->3	
vet n	a->1	i->3	å->1	
vet o	c->9	m->12	
vet p	o->1	å->10	
vet r	e->1	i->1	
vet s	k->4	o->4	t->1	ä->1	å->3	
vet t	i->1	r->1	
vet u	p->3	t->4	
vet v	a->3	i->7	
vet ä	n->1	r->11	
vet" 	o->1	
vet, 	a->1	d->3	e->2	h->1	i->1	j->1	k->1	m->1	n->2	o->7	s->1	t->1	v->4	ä->2	
vet. 	K->1	
vet.D	e->7	
vet.E	f->1	t->1	
vet.F	r->1	ö->2	
vet.H	ä->1	
vet.I	 ->1	
vet.J	a->4	
vet.M	e->1	i->1	
vet.N	ä->1	
vet.R	e->1	
vet.S	å->1	
vet.T	i->1	
vet.V	i->1	
veta 	-->1	a->9	d->1	f->2	h->1	m->1	o->5	v->7	
veta,	 ->1	
vetan	d->4	
veten	 ->14	h->1	s->70	
veter	a->8	i->3	l->1	
vetet	 ->8	
vetna	 ->17	
vets 	a->1	d->1	i->1	m->1	o->2	p->1	r->1	s->1	t->3	
vetss	k->1	
vette	-->1	
vetti	g->3	
vettv	i->1	
vetvi	s->27	
vetyd	i->7	
veuro	p->1	
vfall	 ->5	,->1	.->5	e->8	s->6	
vfolk	n->1	
vförd	 ->1	
vförm	å->1	
vförs	 ->1	l->3	
vfört	r->1	s->1	
vgase	r->1	
vgav 	s->1	
vge e	n->3	
vger 	e->2	i->1	j->1	v->1	
vges 	p->1	
vgett	 ->1	
vgick	,->2	.->2	
vgift	 ->1	e->3	
vgivi	t->1	
vgjor	d->1	t->3	
vgrän	s->4	
vgå.S	o->1	
vgåen	d->1	
vgång	 ->2	e->1	
vgår 	f->1	
vgått	 ->1	
vgör 	h->1	
vgöra	 ->4	n->51	s->2	
vgörs	 ->3	
vhet 	i->1	
vhjäl	p->3	
vhjär	t->1	
vhänd	e->1	
vhäng	i->1	
vhåll	a->1	
vi - 	d->1	j->1	r->1	
vi 19	9->1	
vi 55	 ->1	
vi Eu	r->2	
vi In	t->1	
vi Li	b->1	
vi Pr	o->1	
vi a)	 ->1	
vi ab	s->3	
vi ac	c->1	
vi ag	e->2	
vi al	d->1	l->36	
vi an	a->2	l->1	s->16	t->1	v->10	
vi ar	b->6	
vi at	t->41	
vi av	g->2	s->2	v->3	
vi ba	r->5	
vi be	d->3	f->9	h->26	k->4	n->1	r->5	t->5	v->1	
vi bi	b->1	d->2	
vi bl	a->1	e->1	i->4	
vi bo	k->1	r->9	
vi br	u->1	å->1	
vi by	g->1	
vi bö	r->27	
vi da	g->1	
vi de	 ->1	l->2	m->1	n->8	s->3	t->11	
vi di	r->1	s->14	
vi do	c->1	
vi dr	a->1	
vi dä	r->6	
vi då	 ->6	
vi ef	f->1	t->4	
vi eg	e->3	
vi ek	o->1	
vi em	e->5	
vi en	 ->10	a->1	h->1	i->1	l->1	
vi er	f->1	k->2	
vi et	t->9	
vi eu	r->2	
vi ev	e->1	
vi ex	p->1	
vi fa	k->6	r->2	s->3	t->3	
vi fi	c->1	n->1	
vi fo	k->1	r->12	
vi fr	a->3	å->3	
vi fu	l->2	n->1	
vi få	 ->3	r->10	t->5	
vi fö	l->1	r->40	
vi ga	n->1	
vi ge	 ->3	n->6	r->6	
vi gi	c->1	
vi gj	o->4	
vi gl	a->1	ä->2	ö->1	
vi go	d->4	
vi gr	a->1	u->1	
vi gä	r->2	
vi gö	r->19	
vi ha	 ->4	d->6	f->2	n->2	r->121	
vi he	l->7	
vi hi	t->5	
vi hj	ä->1	
vi ho	p->4	
vi hä	n->1	r->12	v->1	
vi hå	l->7	
vi hö	l->1	r->1	
vi i 	E->3	I->1	M->1	P->1	a->1	d->22	e->3	f->1	g->1	j->1	k->2	m->7	o->1	s->8	v->3	
vi ia	k->1	
vi ib	l->2	
vi ig	å->1	
vi in	b->1	f->3	g->3	h->1	l->4	n->1	o->2	r->2	s->8	t->108	v->1	
vi ju	 ->3	s->8	
vi ka	l->1	n->64	
vi kl	a->2	
vi kn	y->1	
vi ko	m->35	n->6	
vi kr	y->1	ä->3	
vi ku	n->7	
vi kv	a->1	
vi kä	n->2	
vi la	g->3	
vi li	b->1	d->1	k->1	t->4	
vi lo	v->1	
vi ly	c->3	s->2	
vi lä	g->7	m->1	r->1	
vi lå	t->2	
vi me	d->18	n->2	
vi mi	n->1	s->2	
vi mo	d->1	t->2	
vi my	c->1	
vi må	n->1	s->62	
vi na	t->4	
vi nu	 ->21	
vi ny	l->2	
vi nä	r->6	
vi nå	 ->1	g->1	
vi ob	j->1	
vi oc	h->2	k->29	
vi of	f->1	t->1	
vi om	 ->1	
vi os	s->9	
vi pl	a->1	ö->1	
vi pr	o->1	
vi på	 ->11	b->1	
vi re	a->1	d->8	s->4	
vi ri	k->1	m->1	
vi ro	p->1	
vi ru	s->2	
vi rä	k->2	
vi rå	d->1	
vi rö	s->7	
vi sa	d->1	k->1	m->4	
vi se	 ->11	n->1	r->5	
vi sj	u->1	ä->3	
vi sk	a->54	i->2	r->1	u->10	y->1	
vi sl	i->2	ö->1	
vi sn	a->8	
vi so	c->3	l->1	m->12	
vi sp	e->2	
vi st	y->1	ä->10	å->5	ö->8	
vi sv	å->1	
vi sy	m->1	s->1	
vi sä	g->3	k->1	r->2	
vi så	 ->2	g->1	l->1	
vi t.	e->1	
vi ta	 ->2	c->2	g->2	l->11	r->7	
vi te	m->1	
vi ti	d->2	l->12	t->1	
vi to	l->1	
vi tr	e->1	o->6	ä->1	
vi tv	ä->1	
vi ty	c->4	d->1	v->2	
vi tä	n->4	
vi un	d->7	
vi up	p->17	
vi ur	 ->1	
vi ut	a->3	f->1	s->1	t->3	v->5	
vi va	r->9	
vi ve	l->1	m->1	r->8	t->12	
vi vi	d->3	l->28	s->3	
vi vä	l->2	n->4	
vi vå	r->3	
vi yt	t->1	
vi äg	n->4	
vi än	 ->1	d->4	n->5	
vi är	 ->28	
vi äv	e->5	
vi ål	ä->1	
vi år	 ->1	
vi ås	t->1	
vi åt	e->3	m->1	
vi ön	s->5	
vi öv	e->3	
vi, g	i->1	
vi, j	a->2	u->1	
vi, k	a->1	
vi, l	i->1	
vi, m	e->1	
vi, n	ä->1	
vi, s	e->1	o->4	
vi, t	r->1	
vi, ä	n->1	v->1	
vi.Vi	 ->1	
vi?.H	e->1	
via B	r->1	
via E	u->1	
via R	o->1	
via a	l->1	
via b	i->1	
via d	e->1	
via e	n->1	
via k	o->1	
via o	m->1	
via s	t->1	
via t	y->1	
via u	n->1	
viano	 ->1	
vic i	 ->1	
vice 	o->11	t->2	
vice.	A->1	J->1	O->1	S->1	
vicek	o->1	v->1	
vicen	,->1	
vicks	i->3	
vid 1	2->1	
vid 7	0->1	
vid B	y->3	
vid E	G->3	u->3	
vid G	e->1	
vid H	a->1	
vid K	y->1	
vid L	a->1	
vid M	e->1	
vid P	a->1	
vid a	)->1	l->2	n->6	r->1	t->3	v->1	
vid b	e->5	r->1	ö->1	
vid d	a->1	e->32	o->2	
vid e	f->1	n->5	t->8	v->1	
vid f	a->2	l->6	r->4	ö->9	
vid g	o->1	r->2	
vid h	a->4	j->1	ö->1	
vid i	n->1	
vid j	o->1	ä->1	
vid k	o->5	u->2	ä->1	
vid l	i->1	
vid m	a->1	i->1	å->1	ö->2	
vid n	a->1	u->1	y->1	ä->1	å->1	
vid o	f->1	m->6	r->1	
vid p	a->2	l->2	r->2	u->2	å->1	
vid r	e->4	ä->1	
vid s	a->3	i->6	j->1	k->2	l->1	t->3	ä->1	
vid t	e->1	i->4	o->2	r->4	v->1	
vid u	p->3	t->11	
vid v	a->4	i->3	å->1	
vid å	r->2	
vid ö	v->2	
vid, 	a->2	
vid.H	a->1	
vid.J	a->1	
vida 	G->1	a->1	b->1	d->10	i->2	k->2	m->1	n->2	u->1	
vidar	e->37	
vidd 	b->1	h->1	o->1	
vidd.	J->1	
vidde	n->1	
vider	 ->2	.->1	a->7	i->11	s->1	
vidga	 ->14	?->1	d->5	r->3	s->13	t->2	
vidgn	i->71	
vidhå	l->4	
vidhö	l->1	
vidla	g->1	
vidma	k->1	
vidst	r->1	
vidta	 ->33	g->6	l->1	r->8	s->14	
vidto	g->2	
vidua	l->1	
vidue	l->7	
vienn	e->1	
viens	 ->1	
vier 	D->1	
vifta	r->1	
vig v	a->1	
vigla	n->1	
vigt 	b->1	
vigt,	 ->1	
vigt.	D->1	
vigva	t->1	
vigör	 ->1	
vika 	a->7	d->5	e->3	f->1	i->2	m->1	n->2	o->1	s->2	t->1	v->2	
vikan	d->4	
vikas	 ->2	.->2	
vikel	s->5	
viken	 ->2	
viker	 ->6	
viket	 ->1	
vikit	 ->1	
vikli	g->4	
vikna	.->1	
vikt 	a->1	f->1	l->2	m->1	o->1	p->1	s->1	v->7	
vikt,	 ->2	
vikt.	O->1	R->1	
vikt;	 ->1	
vikte	n->12	
vikti	g->328	
viktn	i->3	
vikts	f->1	m->1	
vil e	l->2	
vil s	o->1	ä->2	
vil- 	o->1	
vila 	s->3	
vilar	 ->3	
vilbe	f->2	
vilda	 ->1	
vileg	e->2	i->4	
vilfö	r->2	
vilig	i->1	
vilis	a->1	e->1	
vilja	 ->181	,->2	.->2	d->3	n->18	r->6	s->7	t->8	
vilje	m->1	s->1	
vilka	 ->88	s->2	
vilke	n->49	t->178	
vill 	-->1	I->1	M->1	a->29	b->38	d->23	e->8	f->31	g->28	h->27	i->19	j->98	k->9	l->6	m->6	n->7	o->27	p->10	r->4	s->57	t->36	u->15	v->33	ä->11	å->2	ö->2	
vill,	 ->8	
vill.	J->1	V->1	
ville	 ->10	
villi	g->19	n->1	
villk	o->63	
villo	r->1	
vilrä	t->1	
vilse	 ->1	l->2	
vilsk	y->2	
vilt 	s->1	
vilt,	 ->1	
vin E	u->1	
vin o	c->1	
vind 	o->1	
vindf	ä->4	
vinga	 ->6	d->5	n->5	r->5	s->10	t->1	
vinis	t->1	
vinke	l->11	
vinkl	a->1	
vinna	 ->18	,->1	.->1	s->9	
vinne	r->18	
vinni	n->49	
vinnl	i->2	
vinno	p->2	r->59	
vinns	 ->1	.->1	
vins 	l->1	å->1	
vinse	r->1	
vinst	 ->3	e->6	i->1	m->1	s->1	
virke	s->3	
virra	d->2	n->1	t->1	
virri	n->8	
virrv	a->1	
vis -	 ->3	
vis A	l->1	
vis G	o->1	
vis a	l->3	n->4	t->12	v->4	
vis b	a->2	e->4	r->2	å->1	
vis d	e->8	ä->1	
vis e	l->1	n->4	t->1	x->1	
vis f	i->2	o->1	r->3	u->1	y->1	å->2	ö->4	
vis g	e->2	o->3	r->1	ä->1	å->2	
vis h	a->7	e->1	j->1	o->1	ä->1	ö->1	
vis i	 ->5	l->1	n->16	
vis k	a->2	e->1	o->3	
vis l	e->1	i->1	o->1	
vis m	e->4	i->3	y->1	å->3	
vis n	ä->1	
vis o	a->1	c->16	m->5	r->1	t->1	
vis p	e->2	r->1	å->8	
vis r	e->1	o->1	ä->1	
vis s	a->2	e->1	j->1	k->10	m->1	o->3	t->3	v->1	ä->2	å->3	
vis t	a->1	e->1	i->1	
vis u	n->2	t->3	
vis v	i->8	ä->2	
vis ä	n->1	r->13	v->4	
vis å	s->1	t->1	
vis ö	v->3	
vis) 	f->1	
vis, 	E->1	a->2	d->2	e->1	k->1	m->2	n->1	o->2	p->1	s->2	t->1	v->1	
vis. 	M->1	
vis.D	a->1	å->1	
vis.E	f->1	
vis.H	u->1	
vis.J	a->1	
vis.M	e->1	
vis.S	e->1	
vis.Ä	n->1	
visa 	(->1	R->1	a->7	b->2	d->3	e->2	f->2	g->1	h->2	i->7	k->1	l->1	m->1	o->3	p->4	s->9	t->10	u->1	v->4	ä->3	
visa,	 ->8	
visa.	.->1	B->1	D->4	E->1	F->1	J->1	K->1	R->1	S->1	U->1	Å->1	
visa?	P->1	
visad	e->19	
visan	 ->4	.->1	d->2	s->1	
visar	 ->66	,->2	.->1	e->2	
visas	 ->9	,->1	
visat	 ->32	,->1	.->2	s->3	
visav	i->1	
visba	r->1	
visbe	s->9	
visbö	r->7	
visdo	m->1	
visen	 ->3	
viser	a->6	i->3	
viset	 ->7	.->1	
visfi	s->3	
vishe	t->3	
visio	n->24	
visk 	d->1	
viska	d->1	
viskv	o->2	
vism 	ö->1	
visni	n->14	
visor	.->2	i->2	n->1	
viss 	b->1	f->4	h->1	i->1	m->7	o->4	p->2	r->1	s->2	t->5	u->2	v->1	å->3	ö->1	
vissa	 ->127	.->1	d->2	
visse	r->11	
vissh	e->4	
visso	 ->5	,->1	
visst	 ->6	e->4	
vist 	E->3	P->1	a->3	f->3	o->2	s->2	v->1	
vist,	 ->1	
vista	s->3	t->1	
viste	f->1	l->1	n->1	r->4	
visua	l->1	
visue	l->1	
visum	 ->1	
vit a	l->1	t->1	
vit b	i->1	å->1	
vit d	e->1	
vit e	n->5	t->3	
vit f	r->1	ö->1	
vit g	o->1	
vit h	ö->1	
vit i	n->1	
vit l	e->1	i->1	o->1	
vit m	y->1	
vit o	c->1	
vit s	e->1	i->1	j->1	p->1	y->1	å->2	
vit t	a->1	i->1	
vit u	n->3	t->3	
vit v	a->1	
vit.F	ö->1	
vitbo	k->50	
vitet	 ->11	,->5	.->7	e->14	s->2	
vits 	a->3	f->1	i->3	m->1	s->1	
vits,	 ->1	
vitt 	i->1	v->1	
vittn	a->3	e->2	
vivel	 ->25	,->2	a->3	s->3	
vivla	 ->1	.->1	d->1	r->5	t->2	
vjas 	i->1	
vjett	i->1	
vju m	e->1	
vju s	o->1	
vjuad	e->1	
vkart	a->1	
vklar	 ->2	a->2	t->17	
vkons	t->1	
vkost	n->1	
vkraf	t->3	
vkräv	a->1	
vkunn	a->1	
vla d	e->1	
vla f	ö->1	
vla s	o->1	
vla v	i->1	
vla ä	r->1	
vla" 	s->1	v->1	
vla.V	i->1	
vlade	 ->4	
vlagt	 ->1	
vlan"	.->1	
vlar 	i->3	p->1	s->1	v->1	
vlat 	p->1	v->1	
vledd	a->2	
vlig 	m->1	s->1	
vlig.	O->1	
vliga	 ->3	
vlige	n->1	
vligh	e->1	
vligt	 ->2	
vling	 ->1	
vlist	a->2	
vliva	s->1	
vlopp	e->1	
vlägg	a->1	
vlägs	e->4	n->5	
vlåde	f->1	
vmatt	n->1	
vmilj	o->1	
vna a	v->1	
vna b	e->1	i->2	
vna c	e->1	
vna f	ö->2	
vna i	 ->1	
vna ä	n->1	
vnad 	a->1	b->1	k->1	s->1	
vnad,	 ->2	
vnad.	H->1	
vnad?	V->1	
vnade	n->1	r->1	
vnads	n->1	s->3	v->2	
vning	 ->14	,->2	.->4	a->8	e->2	s->6	
vo (K	O->2	
vo Tr	a->1	
vo at	t->1	
vo bä	r->1	
vo fr	å->1	
vo fö	r->2	
vo ha	r->1	
vo in	t->1	
vo ka	n->1	
vo kä	m->1	
vo me	d->1	
vo oc	h->6	k->1	
vo ti	l->1	
vo ut	a->1	
vo va	r->1	
vo är	 ->3	
vo, e	l->1	t->1	
vo, h	e->1	
vo, i	 ->1	
vo, m	e->1	o->1	
vo, o	c->3	
vo, s	o->1	
vo, v	i->1	
vo.- 	(->1	
vo.Av	s->1	
vo.De	t->2	
vo.Eu	r->1	
vo.Fö	r->1	
vo.He	r->1	
vo.Ko	m->1	
vo.Lå	t->1	
vo.Me	n->1	
vo.Oc	h->1	
vo.Vi	 ->1	
vo? D	e->1	
vo?Hu	r->1	
voNäs	t->1	
voffe	n->1	
vokat	 ->2	.->1	e->2	
vokon	f->1	
vokri	g->1	
volun	t->4	
volut	i->1	
volve	r->9	
volym	 ->2	e->2	
von B	o->1	
von E	i->1	
von W	o->16	
vor t	i->1	
vor.L	i->1	
vorda	 ->2	
vore 	b->2	d->5	e->6	f->3	h->1	i->2	l->1	m->2	o->3	p->1	t->1	v->1	ö->1	
vorit	l->1	
vos a	l->1	
vos d	e->1	
vos e	x->1	
vos l	e->1	
vos m	i->1	
vos s	e->1	
vos y	t->1	
vot p	å->1	
vot s	k->1	
vot v	i->1	
vot ä	r->1	
vot!D	e->1	
vot, 	v->1	
voten	 ->2	.->1	
voter	 ->1	.->1	i->5	n->3	
votum	 ->1	
voår 	f->1	
vplåg	e->1	
vpric	k->1	
vrade	s->1	
vrak 	m->1	s->2	ö->1	
vrak,	 ->1	
vrak.	D->2	
vrak?	N->1	
vrake	t->2	
vrand	e->1	
vrapp	o->1	
vrar,	 ->1	
vras,	 ->1	
vredg	a->1	
vregl	e->2	
vrida	 ->1	
vride	n->1	r->5	
vridn	i->7	
vrig 	i->1	
vriga	 ->31	,->1	.->1	
vrigt	 ->30	,->2	
vrik 	e->1	
vrièr	e->1	
vrund	a->1	
vräkt	s->1	
vräng	a->1	d->1	
vrätt	 ->1	,->1	.->1	a->1	e->1	
vs av	 ->6	
vs be	s->1	
vs de	t->13	
vs dr	a->1	
vs ef	t->1	
vs eg	e->1	
vs en	 ->14	e->1	l->1	
vs et	t->2	
vs fr	a->1	
vs fö	r->9	
vs ge	n->1	
vs ha	n->1	r->2	
vs i 	a->2	d->5	e->1	h->1	v->1	
vs in	g->2	t->1	
vs kr	a->1	
vs me	l->1	r->2	
vs my	c->1	
vs nå	g->1	
vs oc	h->2	k->1	
vs om	f->1	
vs pr	e->1	
vs på	 ->1	
vs ra	m->1	
vs sk	a->1	
vs so	m->4	
vs sp	e->1	
vs st	a->1	
vs sä	k->1	
vs så	 ->1	l->1	
vs up	p->1	
vs ut	 ->1	a->1	
vs ve	r->2	
vs vi	d->2	
vs är	 ->1	
vs öv	e->1	
vs, f	r->1	ö->1	
vs, m	e->4	
vs, o	c->2	
vs, s	å->2	
vs. 1	1->2	
vs. E	q->1	
vs. W	a->1	
vs. a	r->1	t->10	
vs. d	e->4	
vs. e	n->1	r->1	t->1	
vs. f	o->1	ö->2	
vs. g	r->1	
vs. h	o->1	u->1	
vs. i	 ->1	d->1	n->3	
vs. j	a->1	
vs. m	a->2	e->1	i->1	
vs. n	ä->1	
vs. o	m->2	
vs. p	å->1	
vs. s	p->1	
vs. v	a->1	i->1	
vs.Al	l->1	
vs.De	 ->1	t->2	
vs.Et	t->2	
vs.Fr	å->1	
vs.I 	k->1	
vs.Re	s->1	
vs.Sa	n->1	
vs.Sl	u->1	
vs.Vi	 ->1	
vs?Ti	l->1	
vsakn	a->4	
vsarb	e->3	
vsatt	 ->2	a->1	e->1	
vscyk	e->3	
vsdug	l->2	
vse f	o->1	
vsedd	 ->2	a->1	
vseen	d->47	
vser 	E->1	a->5	b->1	d->1	e->1	h->1	m->1	n->2	r->1	v->1	
vses 	g->1	
vsett	 ->13	,->1	
vsevä	r->14	
vsfor	s->1	
vsför	o->1	
vsida	n->1	
vside	s->1	
vsikt	 ->25	e->7	l->4	s->2	
vsind	u->1	
vskaf	f->19	
vsked	.->1	a->4	
vskil	j->1	
vskog	a->1	
vskon	t->2	
vskra	f->1	
vskrä	c->2	
vskva	l->5	
vsky 	f->1	
vskyv	ä->1	
vslag	,->1	.->1	
vslog	 ->2	
vslut	a->52	n->22	
vslän	d->1	g->1	
vslå 	e->1	m->1	
vslår	 ->1	
vslöj	a->6	
vsman	 ->1	n->1	
vsmed	e->88	
vsmil	j->5	
vsmän	 ->1	n->2	
vsnit	t->4	
vsomr	å->1	
vspeg	l->5	
vsstö	d->2	
vsta 	f->1	
vstam	p->1	
vstes	t->1	
vstod	 ->2	
vstym	p->1	
vstyr	a->4	e->2	
vstän	d->8	g->3	
vstå 	f->7	
vståe	n->1	
vstån	d->11	
vstår	 ->5	
vståt	t->2	
vsupp	e->1	
vsvat	t->1	
vsvil	l->1	
vsäga	n->1	
vsäke	r->1	
vsätt	a->3	n->1	
vt - 	d->1	
vt an	s->1	
vt ar	b->3	
vt at	t->7	
vt be	s->3	
vt bl	y->1	
vt de	 ->1	l->1	t->1	
vt di	r->1	
vt el	e->1	
vt en	 ->2	
vt et	t->1	
vt fr	ä->1	
vt fu	n->1	
vt fö	r->6	
vt ha	r->2	
vt hö	g->1	
vt i 	K->1	e->1	f->2	
vt in	f->4	t->1	
vt ka	n->3	
vt ko	m->1	
vt me	d->2	
vt mo	t->1	
vt my	c->1	
vt nå	g->1	
vt oc	h->12	
vt om	 ->3	f->1	
vt ot	i->1	
vt pr	o->2	
vt på	 ->4	
vt re	g->1	s->1	
vt rä	t->2	
vt sa	m->2	
vt se	 ->1	d->1	
vt si	n->1	
vt sk	u->1	y->1	
vt sn	a->1	
vt so	m->2	
vt sp	r->1	
vt st	e->1	r->1	ä->1	ö->2	
vt sv	a->2	
vt sä	k->2	t->13	
vt ta	l->1	
vt ti	l->6	
vt ut	n->1	p->1	
vt ve	r->1	
vt yt	t->1	
vt är	 ->1	
vt ål	ä->2	
vt år	 ->1	,->1	
vt ök	a->1	
vt, d	e->1	ä->1	
vt, i	n->1	
vt, m	e->1	
vt, o	c->1	
vt, p	r->1	
vt, r	ä->1	
vt. D	e->1	
vt.De	t->2	
vt.En	 ->1	
vt.In	t->1	
vt.Pa	r->1	
vt.Äv	e->1	
vtal 	-->1	b->1	d->1	e->1	f->2	i->5	m->12	o->6	r->1	s->15	u->2	v->1	ä->3	
vtal"	 ->1	
vtal,	 ->2	
vtal.	D->1	E->1	F->1	J->1	K->1	
vtal:	 ->1	
vtale	n->6	t->22	
vtals	l->1	
vtar.	V->1	
vtids	b->1	
vtimm	e->2	
vtrup	p->1	
vts d	ä->1	
vts ä	r->1	
vts.E	f->1	
vtvin	g->1	
vud t	a->9	
vudak	t->2	
vudan	g->1	s->4	
vudde	l->3	
vudet	 ->1	
vudfr	å->4	
vudfö	r->1	
vudli	n->2	
vudmå	l->2	
vudre	k->1	
vudro	l->2	
vudsa	k->16	
vudst	a->2	ä->2	
vudsy	f->1	
vudup	p->1	
vulen	 ->1	
vulsk	a->1	
vunds	j->1	
vunge	n->5	
vungn	a->6	
vunna	 ->2	
vunne	n->1	t->1	
vunni	t->7	
vuxit	 ->1	
vuxna	 ->1	.->1	
vvakt	a->6	
vveck	l->8	
vverk	n->2	
vvika	n->4	
vvike	l->1	r->3	
vvisa	 ->2	d->3	n->1	r->3	s->1	t->3	
vvisn	i->2	
vvägd	 ->2	
vvägn	i->1	
vvägs	 ->2	
vvärd	 ->1	a->1	
vyttr	i->1	
väcka	 ->4	n->6	
väcke	r->5	
väcks	 ->1	
väckt	 ->2	e->4	s->1	
väder	 ->1	s->1	
vädja	 ->2	n->1	r->6	
vädre	t->1	
väg [	K->1	
väg a	n->1	t->6	v->1	
väg b	o->1	
väg e	l->6	
väg f	ä->1	ö->1	
väg g	e->2	
väg h	i->1	ä->1	
väg i	 ->1	n->1	
väg k	u->1	
väg m	e->1	o->1	
väg o	c->2	
väg s	i->1	
väg t	r->1	
väg ä	r->1	
väg å	s->1	
väg, 	e->1	f->1	g->1	j->6	o->1	p->1	s->4	v->1	
väg.A	l->1	
väg.B	i->1	
väg.D	e->1	
väg.E	f->1	
väg.J	a->1	
väg.M	e->1	i->1	
väg.O	a->1	
väg.V	a->1	
vägNä	s->1	
väga 	a->4	b->1	d->4	e->2	f->1	h->2	l->1	o->3	s->1	
väga,	 ->1	
väga.	D->1	
vägag	å->6	
vägan	d->8	
vägar	 ->7	,->6	.->5	n->2	
vägby	g->1	
vägd 	g->1	l->1	
vägda	 ->1	
vägen	 ->13	,->2	.->1	:->1	
väger	 ->10	
väggi	g->3	
vägle	d->5	
vägmä	r->1	
vägna	r->16	
vägni	n->1	
vägra	 ->4	d->4	n->5	r->4	s->1	t->4	
vägrö	j->1	
vägs 	g->1	i->1	
vägsk	ä->2	
vägsn	ä->2	
vägso	m->1	
vägt 	d->1	f->1	
väkar	e->1	
väkta	r->2	
väl S	h->1	
väl a	l->1	t->4	v->4	
väl b	e->3	
väl d	e->5	
väl e	k->1	n->2	
väl f	r->1	u->1	ö->5	
väl g	e->2	
väl h	a->3	u->1	
väl i	 ->6	n->5	
väl k	a->2	u->1	v->1	ä->1	
väl l	ä->1	
väl m	a->1	e->6	o->1	y->1	
väl o	c->1	f->1	
väl p	å->3	
väl r	e->3	
väl s	i->1	o->7	t->2	
väl t	i->3	
väl u	n->1	p->1	r->3	t->5	
väl v	a->1	e->1	i->1	å->1	
väl ä	n->2	r->1	
väl å	t->1	
väl ö	v->1	
väl, 	m->1	o->1	
väl.J	a->1	
väl.M	i->1	
väl.S	a->1	
välbe	s->1	
väldi	g->23	
välfu	n->1	
välfä	r->8	
välgr	u->2	
välgö	r->1	
välja	 ->6	r->11	
välje	r->5	
välkl	i->1	
välko	m->50	
välkä	n->3	
väll 	u->1	ä->1	
väll,	 ->2	
väll.	J->1	O->1	
väll?	K->1	
välla	r->1	
välle	n->2	r->1	
välme	n->2	
välmå	e->2	
välsi	g->1	
välst	r->1	å->6	
vält 	o->1	
välta	l->2	
välts	i->1	
välut	b->1	v->2	
välva	n->1	
välvn	i->3	
vämli	g->15	
vämma	d->2	s->1	
vämni	n->4	
vämt 	a->1	
vän o	c->1	
vänd 	b->3	e->1	
vända	 ->49	.->1	m->1	n->2	r->5	s->16	
vändb	a->9	
vände	 ->3	r->32	s->6	
vändi	g->125	
vändn	i->63	
vändp	u->5	
vänds	 ->20	
vänli	g->15	
vänne	r->3	
vänsk	a->1	
vänst	e->14	r->1	
vänt 	d->1	e->1	f->1	l->1	m->1	s->3	
vänta	 ->15	.->1	d->1	n->5	r->39	s->2	t->5	
väntn	i->7	
vänts	 ->5	
väpna	d->2	
värd 	a->3	b->1	d->1	e->2	f->1	m->2	s->1	u->1	
värd.	D->1	
värda	 ->17	,->2	.->1	
värde	 ->6	,->1	.->4	f->7	g->3	l->1	n->18	r->62	s->2	t->4	
värdi	g->27	
väret	 ->1	
värld	 ->1	,->2	.->1	e->37	s->14	
värli	g->6	
värna	 ->2	r->1	
värpo	l->2	
värr 	a->1	b->3	d->3	f->3	g->1	h->6	i->4	k->3	o->2	s->4	ä->5	å->1	
värr,	 ->2	
värr.	V->1	
värra	 ->1	s->2	t->1	
värre	 ->5	,->1	
värs 	m->1	
värst	 ->1	a->7	
värt 	a->11	e->2	f->1	k->1	m->2	s->1	
värt,	 ->3	
värt.	O->1	S->1	V->1	
värto	m->17	
värva	 ->3	d->1	
värvs	a->3	
väsen	 ->2	,->2	d->6	t->26	
västk	u->1	
västr	a->2	
västv	ä->1	
vätsk	a->1	
vätt 	o->1	
vätt,	 ->2	
vätt.	V->1	
vätta	t->1	
väva 	d->1	t->1	
vävna	d->4	
vävt 	s->1	
växa 	u->1	
växa.	H->1	M->1	
växan	d->6	
växel	k->1	v->2	
växer	 ->6	,->1	
växla	n->1	r->1	
växli	n->2	
växt 	a->1	o->4	s->1	ä->1	
växt,	 ->2	
växt.	K->1	O->1	
växtb	r->1	
växte	n->8	r->2	
växth	u->7	
växts	k->3	
vå - 	o->1	
vå ak	t->1	
vå al	t->1	
vå as	p->2	
vå av	 ->8	t->1	
vå be	s->1	t->1	
vå bo	l->1	
vå da	g->1	
vå de	l->1	
vå dä	r->1	
vå el	l->2	
vå et	a->1	
vå eu	r->2	
vå ex	e->2	
vå fa	k->1	l->2	
vå fi	n->1	
vå fl	y->1	
vå fo	k->1	
vå fr	å->4	
vå fö	r->18	
vå ge	n->2	
vå gr	a->1	
vå gå	n->1	
vå ha	r->1	v->1	
vå hu	v->1	
vå i 	d->1	e->1	k->1	
vå in	n->1	s->2	
vå ir	l->1	
vå jo	r->1	
vå ko	l->1	n->1	
vå kr	a->1	
vå kä	r->1	
vå la	g->1	
vå li	k->1	
vå me	d->3	
vå mi	l->2	n->2	
vå my	c->1	
vå må	n->2	s->1	
vå mö	j->1	
vå ne	d->1	
vå ny	c->1	
vå nä	r->1	
vå oc	h->5	
vå of	t->1	
vå ol	i->1	
vå om	 ->1	
vå or	g->1	
vå pe	r->1	
vå pr	i->2	o->1	
vå pu	n->8	
vå på	 ->2	
vå re	g->1	
vå rö	d->1	
vå sa	k->3	
vå se	n->2	
vå sk	ä->2	
vå sm	å->1	
vå so	m->8	
vå st	e->1	o->1	r->1	
vå sä	t->1	
vå så	 ->1	
vå ti	d->1	l->1	m->3	
vå tr	e->2	
vå ty	s->1	
vå un	g->1	
vå up	p->2	
vå ut	a->1	g->1	r->1	
vå ve	c->1	
vå vi	k->5	s->1	
vå yt	t->1	
vå än	 ->1	d->1	
vå är	 ->1	
vå år	 ->5	,->1	s->1	
vå ås	i->1	
vå, a	l->1	
vå, b	ö->2	
vå, d	ä->1	
vå, f	r->1	ö->1	
vå, g	e->1	
vå, m	e->1	
vå, o	c->2	
vå, r	i->1	ö->1	
vå, v	å->1	
vå.At	t->1	
vå.Bi	s->1	
vå.Br	i->1	
vå.De	t->6	
vå.Dä	r->1	
vå.Fö	r->1	
vå.Ge	n->1	
vå.He	r->2	
vå.Ja	g->3	
vå.Jä	m->1	
vå.Me	n->1	
vå.Nä	r->1	
vå.På	 ->1	
vå.Vi	 ->1	
vå: d	e->2	
vå; d	e->1	
vå?Se	r->1	
vådli	g->1	
våer 	g->1	i->3	o->1	s->1	
våer,	 ->2	
våer.	D->2	K->1	M->1	
våer:	 ->1	
våern	a->1	
våg a	v->2	
vågar	 ->5	
vågat	,->1	
vågen	 ->1	
våger	p->1	
våglä	n->1	
vågru	p->3	
våhun	d->1	
våld 	i->1	o->1	
vålde	t->2	
vålds	a->3	h->2	u->1	
våldt	a->2	
vålla	r->1	
vån -	 ->1	
vån f	ö->1	
vån i	 ->2	
vån m	e->1	
vån p	å->3	
vån.D	e->3	
vån.H	ä->1	
våna 	m->1	
vånad	 ->2	e->1	
vånan	d->1	
vånar	e->6	n->5	
vånas	 ->1	
vång 	o->1	
vångr	e->1	
vångs	a->2	f->1	s->1	t->1	
vånin	g->2	
vår a	d->1	t->1	
vår b	a->1	e->6	i->1	u->1	
vår d	e->11	i->1	
vår e	g->1	n->1	r->1	
vår f	a->1	r->5	ö->7	
vår g	e->3	r->12	
vår i	n->4	
vår k	a->3	o->4	u->1	
vår l	a->2	i->2	o->2	
vår m	e->4	i->4	o->1	å->1	
vår n	y->1	
vår o	r->2	
vår p	e->1	l->3	o->4	r->1	
vår r	e->5	o->2	ä->2	ö->1	
vår s	a->2	i->2	k->2	l->1	o->3	p->1	t->6	v->1	
vår t	a->1	i->1	r->1	v->1	
vår u	n->2	p->6	t->1	
vår v	i->3	ä->2	
vår å	s->3	t->1	
vår ö	n->1	
vår, 	E->1	
våra 	a->12	b->4	d->5	e->9	f->16	g->7	h->3	i->5	k->13	l->11	m->17	n->2	o->2	p->9	r->15	s->14	t->6	u->1	v->4	ä->4	å->6	ö->4	
våra,	 ->1	
vårar	 ->1	e->4	
vårbe	d->1	g->1	
vård 	o->2	
vård)	,->1	
vård,	 ->1	
vårds	-->1	l->2	m->1	
våret	 ->2	
vårig	h->31	
vårlö	s->2	
vårss	k->2	
vårt 	E->2	a->33	b->3	d->4	e->10	f->13	g->3	h->1	i->2	k->4	l->4	m->4	n->2	o->3	p->11	r->2	s->14	t->2	u->11	v->3	y->1	
vårt,	 ->2	
våröv	e->1	
vö, f	ö->1	
vö.De	t->1	
vön s	o->1	
vördn	a->1	
w Yor	k->1	
w för	 ->1	
w til	l->1	
w, so	m->1	
w-how	 ->1	
w.Med	 ->1	
wagen	!->1	
wald,	 ->1	
wales	a->1	
wan i	n->1	
warzw	a->1	
we.Eu	r->1	
we.Vi	 ->1	
webbp	l->1	
weiz,	 ->1	
wells	k->1	
wer k	o->1	
wer, 	e->1	s->1	
wies 	v->1	
will 	f->1	
wis h	a->1	
wis n	ä->1	
witts	b->1	
witz.	 ->1	
wn av	 ->1	
wn är	 ->1	
wn, m	e->1	
wobod	a->3	
wood 	o->1	
woodf	i->1	
woods	 ->1	
worst	 ->1	
x all	v->1	
x ant	e->4	
x av 	p->1	
x avs	l->1	
x eft	e->1	
x eur	o->1	
x fle	r->1	
x inn	a->1	
x min	u->1	
x mån	a->10	
x och	 ->1	
x pla	t->1	
x pos	t->1	
x sad	e->1	
x til	l->1	
x tun	c->1	
x öve	r->1	
x!Jag	 ->1	
x, ja	g->1	
x, no	r->1	
x, nä	m->1	
x, sj	u->1	
x, so	m->1	
x-aff	ä->1	
x-fre	e->3	
x. Eu	r->1	
x. Fr	a->1	
x. Ne	d->1	
x. US	A->1	
x. at	t->1	
x. av	 ->1	
x. de	n->1	t->1	
x. et	t->1	
x. in	o->1	
x. ku	n->1	
x. kä	n->1	
x. mi	t->2	
x. nä	r->1	t->1	
x. ol	j->1	
x. på	 ->1	
x. ut	f->1	
x. va	r->1	
x.De 	b->1	
x.Jag	 ->1	
xa et	t->1	
xa ut	 ->2	
xa, t	i->1	
xa.Hä	r->1	
xa.Me	d->1	
xakt 	d->4	h->2	l->1	m->1	o->1	v->1	
xakt,	 ->1	
xakta	 ->6	
xakth	e->1	
xal s	i->2	
xala 	s->1	
xalt 	n->1	o->1	
xamen	 ->3	,->1	s->2	
xamin	a->1	e->9	
xan?V	e->1	
xande	 ->6	r->2	
xas d	a->5	
xas g	u->1	
xas i	 ->1	
xat u	p->1	
xbelo	p->1	
xcept	i->6	
xelku	r->1	
xelry	c->1	
xelve	r->2	
xembu	r->6	
xempe	l->110	
xempl	a->2	e->6	
xen s	k->1	
xer d	i->1	
xer f	r->1	
xer o	c->2	
xer s	a->1	i->1	
xer, 	v->1	
xerin	g->1	
xfick	o->1	
xhave	n->1	
xibel	 ->3	,->1	.->1	t->6	
xibil	i->10	
xibla	 ->3	.->1	r->2	
xid i	 ->1	
xid o	c->3	
xidut	s->1	
xiko,	 ->1	
xilre	g->1	
xilti	b->1	
ximal	 ->1	a->2	t->3	
ximer	a->2	
ximiå	l->1	
xin o	c->1	
xinkr	i->1	
xis a	t->1	
xis i	n->1	
xis s	o->1	t->1	
xis ä	r->1	
xis.D	e->1	
xis.F	ö->1	
xisen	 ->1	
xiska	 ->1	
xisme	n->1	
xiste	n->6	r->13	
xit u	p->1	
xklus	i->3	
xland	e->1	
xlar 	s->1	
xlar.	F->1	
xling	 ->1	a->1	
xmåna	d->1	
xna e	l->1	
xna.H	e->1	
xning	e->1	
xon V	a->3	
xor.D	e->1	
xpand	e->5	
xpans	i->1	
xpedi	t->1	
xpert	e->20	g->3	i->3	k->17	r->2	u->1	
xplic	i->1	
xplos	i->2	
xpone	n->1	r->1	
xport	 ->1	e->3	
xt av	 ->1	s->1	
xt få	r->1	
xt i 	m->1	
xt ko	m->1	
xt li	g->1	
xt oc	h->6	
xt om	 ->1	
xt sk	a->1	
xt so	m->5	
xt är	 ->1	
xt, i	n->1	
xt, o	m->1	
xt, s	o->3	å->1	
xt, ä	r->1	
xt.Ko	n->1	
xt.Me	n->1	
xt.Oc	h->1	
xtbra	n->1	
xten 	-->1	e->1	f->1	g->1	i->6	k->1	o->1	r->1	s->2	t->1	ä->1	
xten"	.->2	
xten,	 ->4	
xten.	D->1	F->1	
xter 	f->1	o->1	ä->1	
xter,	 ->2	
xter.	L->1	N->1	P->1	
xtern	a->11	
xthus	e->3	g->4	
xton.	V->1	
xtra 	E->1	f->1	r->1	s->2	
xtran	d->1	
xtrao	r->1	
xtrem	a->2	h->14	i->10	t->4	
xtsky	d->3	
xuell	 ->1	.->1	t->1	
xupér	y->1	
xvärt	 ->1	
xxon 	V->3	
y - s	a->1	
y Can	y->3	
y Eur	o->1	
y For	d->1	
y bil	.->1	
y den	 ->1	
y det	 ->2	t->1	
y end	 ->1	
y enl	i->1	
y eur	o->1	
y fas	c->1	
y for	m->1	
y för	 ->4	o->2	
y gra	n->1	
y han	 ->1	
y har	 ->1	
y här	 ->1	
y i h	ö->1	
y inf	o->1	
y ing	e->1	
y ins	t->1	
y kem	i->1	
y kom	m->3	
y kul	a->2	t->1	
y kva	l->1	
y lag	s->1	
y led	a->1	
y liv	s->1	
y myn	d->1	
y nat	u->1	
y när	 ->1	
y och	 ->3	
y olj	a->1	
y per	i->1	s->1	
y på 	d->1	s->1	
y rös	t->2	
y sek	t->1	
y sit	u->1	
y som	 ->1	
y spe	c->1	
y sto	r->1	
y syn	v->1	
y sys	s->1	
y typ	 ->1	
y und	e->1	
y upp	m->1	
y var	 ->1	
y vet	e->1	
y vi 	h->1	k->2	v->1	
y vig	ö->1	
y vit	b->1	
y är 	r->1	
y åte	r->1	
y! Ge	n->1	
y, Ha	v->1	
y, Jo	n->1	
y, at	t->1	
y, de	r->1	
y, ha	r->1	
y, ka	d->1	
y, kv	i->1	
y, so	m->1	
y, st	r->1	
y-pro	t->1	
y.And	r->1	
y.De 	b->1	
y.Vi 	h->1	k->1	
yDe f	ö->1	
ya "l	ä->1	
ya 81	 ->1	
ya EU	-->1	
ya Eu	r->2	
ya Ze	e->2	
ya ar	b->7	t->2	
ya at	t->1	
ya av	t->2	
ya be	f->2	s->4	
ya bi	l->6	
ya bu	d->1	
ya by	r->1	
ya de	l->1	m->1	
ya di	r->2	
ya do	m->1	
ya eu	r->1	
ya ex	t->1	
ya fe	m->1	
ya fr	a->1	i->1	å->1	
ya fö	d->1	r->5	
ya ge	m->2	
ya gr	u->1	
ya im	p->1	
ya in	i->2	s->1	
ya jo	b->1	
ya kl	i->1	
ya ko	a->1	m->14	n->1	
ya la	g->1	
ya le	d->1	
ya li	v->1	
ya lä	n->4	
ya ma	r->1	
ya me	d->8	
ya mi	t->1	
ya mo	d->1	
ya my	n->2	
ya må	l->1	
ya mö	j->3	
ya no	r->1	
ya nä	t->1	
ya ob	e->1	
ya oc	h->2	
ya om	r->1	s->1	
ya or	d->1	
ya pa	r->1	
ya pe	n->1	r->2	
ya pr	e->1	i->1	o->7	
ya ra	m->1	
ya re	g->10	s->1	
ya ri	k->2	
ya ru	n->1	
ya rä	t->2	
ya si	t->1	
ya sp	ö->1	
ya sy	s->4	
ya sä	t->1	
ya te	k->4	
ya ti	l->1	
ya tj	ä->2	
ya ty	s->1	
ya up	p->1	
ya ut	m->1	v->1	
ya ve	r->2	
ya vi	t->1	
ya vå	l->1	
ya än	d->2	
ya år	e->1	
ya åt	g->5	
ya, u	t->1	
ya; k	o->1	
yaber	g->1	
yabuk	t->2	
yagol	f->4	
yal U	l->1	
yande	t->1	
yanna	k->2	
yanse	r->1	
yanst	ä->2	
yar l	i->1	
yarbe	t->1	
yas o	c->1	
yaste	 ->1	
yavta	l->1	
ybar 	e->4	
ybar,	 ->1	
ybara	 ->34	
ybetä	n->2	
ybila	r->1	
ybils	k->1	p->1	
yck a	n->1	v->6	
yck e	f->1	
yck f	r->1	ö->9	
yck i	 ->2	
yck k	a->1	
yck m	o->1	
yck p	å->1	
yck s	o->1	
yck, 	i->1	m->1	
yck.D	e->1	
ycka 	a->2	d->2	e->1	i->2	m->9	o->2	p->1	s->6	t->2	v->7	ä->1	
ycka,	 ->2	
ycka.	B->1	
ycka?	"->1	
yckad	e->13	
yckan	 ->5	d->9	
yckas	 ->22	,->3	.->1	
yckat	s->20	
yckbä	r->1	
ycke 	f->1	i->1	s->2	t->2	u->1	
ycke.	F->1	H->1	V->1	
yckel	f->3	n->3	p->1	r->1	
ycken	 ->3	
ycker	 ->66	:->1	
ycket	 ->439	!->1	,->20	.->3	?->1	
yckla	n->2	
yckle	r->4	
yckli	g->28	
yckni	n->5	
yckor	 ->13	,->1	.->1	n->1	
yckos	a->1	
ycks 	a->1	d->1	e->1	i->1	m->2	o->1	t->1	v->2	ö->1	
ycksb	å->1	
ycksd	r->3	
ycksf	a->2	
ycksr	i->2	
ycksö	d->1	
yckt 	e->1	k->1	n->1	s->1	
yckte	 ->14	s->2	
yckts	 ->1	
yckön	s->5	
yclin	g->1	
yd ge	n->1	
yd i 	h->1	
yd so	m->1	
yd ti	l->1	
yd.Sa	v->1	
yda m	i->1	
yda u	n->2	
ydafr	i->2	
ydana	n->1	
ydand	e->17	
ydd a	v->4	
ydd b	a->1	
ydd e	l->1	
ydd f	ö->13	
ydd i	 ->1	n->1	
ydd m	o->2	å->1	
ydd o	c->3	
ydd s	a->2	o->1	t->1	
ydd v	i->2	
ydd ö	v->1	
ydd),	 ->1	
ydd, 	d->1	e->1	v->1	
ydd.D	e->2	
ydd.J	a->1	
ydd.N	a->1	
ydd.R	e->1	
ydd.V	i->1	
ydda 	a->1	c->1	d->5	f->2	g->3	l->1	m->5	p->1	s->4	u->1	v->1	
yddad	e->2	
yddan	d->1	
yddar	 ->1	e->1	
yddas	.->2	
ydde 	"->1	a->1	
yddes	 ->1	
yddet	 ->16	,->2	
yddsm	e->4	
yddsn	i->6	
yddso	m->1	r->1	
yddsp	r->1	
yddss	t->1	ä->1	
yddst	u->1	
ydel 	o->1	
ydels	e->75	
yder 	E->1	a->9	d->1	e->1	i->3	l->1	o->1	p->5	u->3	
yder,	 ->1	
yder:	 ->1	
ydeur	o->1	
ydig 	e->1	
ydiga	 ->3	
ydigh	e->4	
ydigt	 ->2	,->1	
ydkor	e->1	
ydkus	t->1	
ydlig	 ->13	,->1	:->1	a->29	e->3	g->4	h->1	t->73	
ydost	a->1	e->1	
yds i	 ->1	
ydväs	t->1	
ydöst	r->1	
ye Pl	a->1	
ye or	d->1	
ye-av	t->2	
yed i	s->2	
yelse	 ->3	n->2	o->1	
yens 	d->1	
yer h	a->1	
yer n	u->1	
yer.O	m->1	
yern,	 ->1	
yetab	l->1	
yfall	 ->1	
yfasc	i->1	
yft f	r->2	
yfta 	b->1	f->3	p->1	
yftad	e->3	
yftan	 ->2	
yftar	 ->30	
yftas	 ->3	
yfte 	a->9	m->1	o->1	s->1	v->1	ä->2	
yfte.	D->1	
yften	 ->4	,->1	a->1	
yfter	 ->2	
yftet	 ->22	
yftor	,->1	n->2	
yförs	l->1	
yförv	ä->1	
yg de	 ->1	
yg fr	a->1	
yg få	r->1	
yg fö	r->3	
yg i 	E->1	t->1	v->2	
yg me	d->3	
yg nä	r->1	
yg ob	e->1	
yg oc	h->1	
yg om	 ->1	
yg so	m->14	
yg så	v->1	
yg un	d->2	
yg ut	a->1	
yg), 	t->1	
yg, d	e->1	
yg, h	a->1	
yg, s	o->1	
yg, u	t->1	
yg.En	l->1	
yg.Fö	r->1	
yg.Va	r->1	
yg.Vi	s->1	
yg; m	i->1	
yg?Dä	r->1	
yga a	t->2	
yga d	e->1	
yga g	e->1	
yga i	g->1	
yga m	e->1	
yga o	c->1	
yga s	i->2	
yga v	i->1	
yga y	t->1	
ygad 	m->1	o->15	
ygade	 ->5	
ygand	e->6	
ygar 	m->1	
ygbla	d->1	
ygd i	 ->1	
ygd o	m->1	
ygd.D	e->2	
ygden	 ->13	,->3	.->7	s->8	
ygdsb	e->1	
ygdsk	o->1	
ygdso	m->4	
ygdsr	e->2	
ygdst	u->1	
ygdsu	t->1	
ygell	ö->1	
ygels	e->4	
ygen 	a->1	e->1	v->1	
ygen,	 ->3	
ygens	 ->7	
yger 	a->1	
yget 	h->1	m->1	s->3	u->1	v->1	
ygets	 ->1	
ygga 	a->2	b->1	d->2	e->3	h->1	i->1	n->1	o->3	r->1	s->2	u->15	v->4	
yggad	e->1	
yggan	d->23	
yggas	 ->3	
yggd 	i->1	p->1	
yggde	 ->1	s->1	
ygge 	s->1	
yggel	s->1	
yggen	 ->3	
ygger	 ->7	
ygget	 ->2	s->2	
ygghe	t->6	
yggna	d->19	
yggor	 ->1	
yggra	d->1	
yggs 	p->1	u->1	
yggst	e->1	
yggt 	i->1	p->1	s->1	u->1	
yggts	 ->1	
ygien	,->1	.->1	
ygkra	s->1	
ygnin	g->1	
ygpla	n->1	t->3	
ygrup	p->2	
ygsam	 ->2	m->2	
ygsbe	s->1	
ygsin	s->1	
ygssk	r->7	
ygsst	å->1	
ygssä	k->1	
ygsta	n->1	
ygsäg	a->1	
ygt 4	0->1	
ygt e	t->1	
ygt t	v->1	
ygtra	n->2	
yhet 	a->1	
yhet.	 ->1	M->1	
yhete	n->1	r->8	
yhets	r->1	
yhun 	s->1	
yhöga	 ->1	
yiste	n->1	r->1	
yk.He	r->1	
yka -	 ->1	
yka P	o->1	
yka a	t->11	
yka d	e->5	
yka e	t->1	
yka f	y->1	
yka m	i->1	
yka s	a->1	
yka u	p->2	
yka v	ä->1	
yka, 	n->1	t->1	
ykas 	a->1	f->2	ä->1	
ykel 	f->1	
ykel,	 ->1	
ykel.	T->1	
yker 	d->2	o->1	u->3	ä->1	
yklar	 ->3	n->1	
ykolo	g->1	
yks o	c->1	
yks v	i->1	
ykta 	d->1	
yktad	 ->1	
yktba	r->1	
ykte 	i->1	o->1	s->2	
ykte,	 ->1	
ykte.	M->1	
ykten	 ->3	
ykter	 ->1	t->2	
yktin	g->13	
yktra	 ->1	
yl ge	n->1	
yl oc	h->3	
yl, f	ö->1	
yl, r	ä->1	
yl- o	c->1	
yl.De	t->1	
yl.Ja	g->1	
yl.Vi	 ->1	
yla.H	e->1	
ylan 	ä->1	
ylbes	l->1	
yldig	 ->3	a->10	e->1	h->15	
ylför	f->2	
ylibe	r->1	
yliga	 ->1	
ylige	n->30	
ylika	 ->2	
ylikt	 ->1	
ylla 	A->1	d->3	e->2	f->1	g->1	h->2	i->1	k->3	s->8	v->3	
ylla.	V->1	
yllan	d->3	
yllas	 ->9	,->1	
yllde	s->1	
yller	 ->21	
yllni	n->1	
yllra	n->1	
ylls 	m->1	o->1	p->1	
ylls.	U->1	
yllt 	s->1	
yllt,	 ->2	
yllts	 ->1	
ylrät	t->2	
ylsök	a->6	
ym at	t->1	
ym me	d->1	
ym om	 ->1	
ym so	m->1	
ym.De	n->1	
yma B	r->1	
ymask	i->1	
ymbol	 ->2	i->7	
ymd t	i->1	
ymden	 ->1	
ymen 	p->1	
ymer 	i->1	
ymite	t->1	
ymma 	e->1	
ymme 	f->6	o->1	s->1	å->2	
ymme,	 ->1	
ymmer	 ->4	.->1	s->1	
ympad	 ->1	
ympat	i->8	
ympic	 ->1	
ympis	k->1	
ympni	n->2	
ympto	m->1	
ymrad	 ->5	e->2	
ymrar	 ->2	
ymrat	 ->1	
yms i	 ->1	
ymt a	t->1	
ymts 	a->1	
yn - 	t->1	
yn at	t->1	
yn av	 ->1	
yn ge	s->1	
yn ha	r->1	
yn i 	a->1	v->1	
yn ly	c->1	
yn oc	h->5	
yn på	 ->4	
yn ti	l->65	
yn va	r->1	
yn än	 ->1	
yn äv	e->1	
yn ål	ä->1	
yn, m	e->1	
yn, o	c->1	
yn.At	t->1	
yn.Et	t->1	
yn.Si	s->1	
yn.Sl	u->1	
yn; d	e->1	
yna h	u->1	
ynami	k->1	s->4	
ynand	e->1	
ynas 	a->1	
ynas.	D->1	J->1	
ynazi	s->6	
ynd a	t->1	
ynd f	ö->1	
ynd g	e->1	
ynd ä	r->1	
ynda 	a->2	k->1	p->1	s->1	
yndab	o->2	
yndan	d->1	
yndar	 ->2	s->1	
yndas	 ->1	.->2	
ynder	 ->1	
yndig	a->2	h->162	
yndro	m->1	
yndsa	m->4	
ynen 	i->2	m->1	p->1	t->1	
ynen.	D->1	
ynerg	i->2	
ynes 	b->1	
yngan	d->1	
yngd 	b->1	n->1	
yngdp	u->4	
ynger	 ->1	
yngre	 ->1	
yngst	.->1	a->2	
ynlig	 ->1	,->1	.->1	a->4	t->1	
ynn, 	d->1	
ynna 	d->1	s->3	u->1	å->2	
ynnad	e->6	
ynnar	 ->5	
ynne 	f->1	
ynne!	 ->1	
ynner	h->46	l->6	
ynnes	 ->2	
ynnsa	m->3	
ynony	m->1	
ynpun	k->29	
yns s	ä->1	
ynsta	g->2	
ynsät	t->4	
ynt n	å->1	
ynt v	å->1	
ynt, 	d->1	
yntes	.->1	
ynvin	k->12	
yo sk	u->1	
yola 	d->2	
yon 1	9->1	
yon s	a->1	
yon, 	O->1	
yosta	d->1	
yoto 	k->1	o->1	
yoto-	p->1	
yoto.	V->1	
yotop	r->2	
yotos	 ->1	
yp Ca	d->1	
yp av	 ->18	
yp få	t->1	
yp, d	e->1	
yp, l	i->1	
yp.De	t->1	
yp.Ef	t->1	
ypen 	a->12	
yper 	a->3	
ypern	 ->1	a->1	
ypfal	l->1	
ypgod	k->1	
yphål	 ->1	:->1	e->1	
yplan	t->1	
ypote	s->1	t->1	
yppas	 ->1	
ypper	l->1	
yps.M	e->1	
ypten	 ->1	,->1	
yptog	a->2	
yr al	l->1	
yr er	 ->1	
yr fr	å->1	
yr hi	s->1	
yr ja	g->1	
yr.Ef	t->1	
yra a	r->1	
yra d	e->3	
yra e	k->1	
yra f	e->1	ö->2	
yra g	e->1	
yra h	e->1	
yra i	n->1	
yra k	ä->2	
yra l	ä->1	
yra m	a->1	å->3	
yra n	y->1	
yra o	m->1	r->1	
yra p	a->1	e->2	u->3	
yra r	o->1	
yra s	a->1	y->1	ä->1	
yra u	n->1	
yra ä	n->2	r->1	
yra å	r->1	t->1	
yra, 	h->1	
yra: 	r->1	
yrami	d->1	
yrand	e->4	
yrar 	d->1	i->2	p->1	t->1	
yrare	 ->1	.->1	
yras 	a->1	
yras.	I->1	
yrd a	v->1	
yre s	o->1	
yre, 	e->1	
yregi	m->1	
yreko	n->3	
yrels	e->7	
yren,	 ->1	
yret 	i->1	
yrets	 ->2	
yrien	 ->13	,->4	.->3	f->1	s->1	
yrier	 ->1	n->5	
yrigh	t->1	
yrisk	a->3	e->1	
yrka 	b->1	f->1	i->1	k->1	m->1	o->2	p->1	
yrka,	 ->1	
yrka.	H->1	
yrkan	 ->4	s->1	
yrkar	 ->1	
yrkef	ö->1	
yrken	 ->3	
yrkep	o->1	
yrkes	a->1	e->1	k->2	l->2	m->1	u->7	v->1	
yrkog	å->1	
yrkor	 ->1	,->1	
yrne 	o->1	
yrne,	 ->1	
yrnin	g->7	
yrs a	v->2	
yrt o	c->1	
yrt. 	I->1	
yrtio	 ->3	s->1	
yrå s	o->1	
yrå ä	r->1	
yråer	,->1	
yråkr	a->30	
yrån 	f->3	
ys - 	o->1	
ys av	 ->16	
ys be	t->3	
ys de	 ->1	
ys fa	l->1	
ys fl	y->1	
ys fö	r->1	
ys ge	n->1	
ys i 	d->1	
ys ja	g->1	
ys oc	h->2	
ys or	d->1	
ys so	m->1	
ys vi	 ->1	
ys, a	l->1	
ys, d	ä->1	
ys, u	t->1	
ys, v	i->1	
ys-de	-->1	
ys.De	n->2	
ys.Fr	u->1	
ys.Ge	n->1	
ys.Hä	r->1	
ys?De	n->1	
ys?I 	s->1	
ysa f	r->1	
ysa m	i->1	
ysa o	m->2	
ysa s	k->1	
ysa u	p->2	r->1	
ysa v	å->1	
ysa ä	n->1	
ysand	e->4	
ysato	r->2	
ysen 	a->3	g->1	m->1	
yser 	b->1	i->2	j->1	s->1	v->2	
yser.	K->1	
ysera	 ->10	r->1	s->3	t->1	
ysisk	 ->2	a->6	t->1	
ysk e	n->1	
yska 	E->1	b->3	d->2	f->3	k->1	l->1	o->3	p->1	r->2	s->2	v->2	
yska,	 ->1	
yskap	a->1	
yskla	n->22	
yskt 	o->1	ö->1	
ysnin	g->5	
yss a	t->1	
yss b	e->1	
yss e	l->1	
yss g	j->1	
yss n	ä->1	
yss o	c->1	m->1	r->1	
yss s	a->2	
yss, 	a->1	i->1	
yss.S	l->1	
yssa 	p->1	
yssar	n->1	
yssel	 ->9	!->1	,->4	-->2	.->1	b->1	f->1	s->103	
yssen	 ->2	,->1	s->2	
yssla	d->1	n->4	r->5	
yssna	 ->9	,->1	d->4	r->5	t->9	
yssni	n->1	
yst f	ö->1	
yst m	i->3	å->1	
ystem	 ->75	,->9	.->11	:->1	a->10	e->81	ä->3	
yster	f->1	i->1	
ystra	 ->1	
yta a	n->1	
yta b	e->1	
yta d	e->3	
yta e	r->1	
yta h	e->1	
yta k	o->1	
yta m	o->4	
yta s	a->1	
yta.I	n->1	
ytand	e->13	
ytas 	s->1	
yte a	v->3	
yte f	ö->2	
yte k	o->1	
yte m	e->2	o->1	
yte s	a->1	
yte, 	r->1	
ytels	e->3	
yter 	e->1	m->2	t->4	v->1	
yteri	n->1	
ytet 	a->2	m->3	p->1	
ytisk	t->1	
ytlig	h->1	t->1	
ytnin	g->3	
yts t	i->1	
ytt I	N->1	
ytt a	r->1	
ytt b	o->1	y->1	
ytt e	n->1	
ytt f	ö->3	
ytt g	e->1	
ytt i	 ->2	n->1	
ytt k	a->1	o->1	
ytt l	y->1	
ytt m	i->2	
ytt o	b->1	m->1	
ytt p	a->2	l->1	o->1	r->1	
ytt s	k->2	o->3	p->1	t->2	y->2	ä->1	
ytt t	a->1	
ytt u	n->1	
ytt v	i->1	
ytt å	r->2	
ytt ö	n->1	v->1	
ytt, 	f->1	m->1	s->1	
ytt.D	e->2	
ytt.J	a->2	
ytta 	a->11	e->1	f->4	o->2	s->1	t->1	
ytta,	 ->1	
ytta.	B->1	F->1	N->1	P->1	
yttan	 ->1	
yttar	 ->3	
yttas	 ->1	
yttat	 ->1	
ytter	d->1	i->2	l->53	o->1	s->33	v->1	
yttig	 ->6	a->4	t->3	
yttja	 ->18	d->4	n->9	r->3	s->6	t->1	
yttni	n->4	
ytto-	a->1	
yttoa	n->1	
yttra	 ->4	n->32	r->1	t->2	
yttre	 ->3	
yttri	n->1	
ytts 	u->1	
yu i 	T->1	
yu sa	m->1	
yvald	a->1	
yveri	e->1	
yverk	s->1	
yvärd	a->1	
yvärr	 ->36	,->2	.->1	
ywood	f->1	
yxfic	k->1	
yårsa	f->1	
z Fis	c->3	
z Flo	r->2	
z Gon	z->1	
z ang	å->1	
z bet	ä->1	
z dyk	e->1	
z ell	e->1	
z en 	g->1	
z ett	 ->1	
z frå	g->1	
z får	 ->1	
z för	 ->1	o->1	
z had	e->1	
z i B	r->1	
z och	 ->7	
z ock	s->1	
z om 	a->1	
z sad	e->2	
z som	 ->2	
z tog	 ->2	
z)(Ta	l->1	
z).He	r->1	
z, Gi	n->1	
z, La	n->3	
z, be	s->1	
z, in	o->1	
z, på	m->1	
z, ta	l->1	
z, ut	r->1	
z-kat	a->3	
z. Eu	r->1	
zFru 	t->1	
za oc	h->1	
za, d	e->1	
za.De	t->1	
za.Si	t->1	
zakst	a->1	
zarem	s->2	
zbeki	s->2	
zbetä	n->1	
zen.J	a->1	
zes-C	a->1	
zidak	i->2	
zigen	a->3	s->1	
zio-P	l->4	
zism 	e->1	o->1	
zism.	D->1	
zisme	n->5	
zist 	o->1	
zist!	T->1	
zista	n->5	
ziste	r->2	
zistf	l->1	
zisti	s->3	
zjiki	s->5	
zmann	,->1	-->1	
zon 3	4->1	
zon V	I->2	
zon o	c->1	
zonen	 ->1	
zoner	.->1	n->1	
zonin	d->1	
zorer	n->2	
zquie	r->1	
zuela	 ->1	
zwald	,->1	
zález	 ->1	
º C. 	D->1	
Ämnar	 ->1	
Än en	 ->3	
Ända 	s->1	
Ändra	s->1	
Ändri	n->13	
Ändå 	a->1	k->3	s->1	
Ännu 	e->1	h->1	s->1	
Äntli	g->1	
Är Is	r->1	
Är de	n->2	t->17	
Är hy	s->1	
Är in	t->1	
Är ko	m->2	
Är rå	d->1	
Är st	a->1	
Är vi	 ->1	
Ärade	 ->6	
Även 	E->2	d->3	h->2	i->3	j->10	k->1	m->2	o->19	p->2	ä->2	
Å EDD	-->1	
Å PSE	-->1	
Å and	r->10	
Å ena	 ->2	
Å kom	m->1	
Å soc	i->1	
ÅDSKA	N->1	
ÅGORN	ä->1	
År 19	9->4	
År 20	0->1	
Året 	s->1	
Årlig	e->1	
Åtaga	n->1	
Återi	n->1	
Återu	p->2	
Återv	i->1	
Åtgär	d->5	
Île-d	e->1	
Ö (Ös	t->2	
Ö för	 ->1	
Ö häv	d->1	
Ö ino	m->1	
Ö min	i->1	
Ö och	 ->3	
Ö om 	d->1	
Ö som	 ->1	
Ö vid	 ->1	
Ö är 	e->1	
Ö) si	n->1	
Ö).Ja	g->1	
Ö-led	a->1	
Ö-med	l->1	
Ö:s a	r->1	
Ö:s d	e->1	
Ö:s f	r->1	
Ö:s s	t->1	
ÖSTNI	N->2	
ÖVP (	Ö->2	
ÖVP a	t->2	
ÖVP m	i->1	
ÖVP) 	o->1	
Ögonb	l->2	
Ökad 	k->1	
Öppen	h->1	
Öster	r->81	
Östeu	r->5	
Östty	s->2	
Över 	8->1	
Överv	ä->1	
Övrig	a->1	
ález 	o->1	
án, a	t->1	
ánche	z->1	
ão To	m->2	
ä utg	ö->1	
ä öve	r->1	
äck m	e->1	
äck o	c->1	
äck s	o->1	
äcka 	a->1	d->1	e->1	f->1	m->2	n->2	r->2	s->4	t->4	u->2	v->1	å->1	
äcka,	 ->1	
äckad	 ->1	
äckan	d->12	
äckas	!->1	
äcken	s->1	
äcker	 ->36	.->1	
äckhe	t->1	
äckla	r->1	
äckli	g->77	
äckni	n->32	
äckor	 ->1	
äcks 	a->3	n->1	s->1	u->1	
äcks.	U->1	
äcks;	 ->1	
äcksc	e->1	
äckt 	f->1	h->2	n->1	s->2	u->1	v->1	ä->1	
äckte	 ->3	s->3	
äckts	 ->2	!->1	
äckvi	d->3	
äd be	h->1	
äd fä	l->1	
äd ha	d->1	r->1	
äd up	p->1	
äd, o	c->1	
äd.De	n->1	
äda E	u->1	
äda e	f->1	
äda i	 ->6	
äda s	o->1	
äda u	p->1	r->1	
äda, 	h->1	
ädand	e->10	
ädare	 ->37	,->5	.->1	?->1	n->1	s->2	
ädarn	a->10	
ädat 	u->1	
ädd a	t->1	v->1	
ädd f	ö->3	
ädd, 	h->1	
ädda 	6->1	a->2	d->1	i->2	k->1	o->1	s->1	
äddad	e->3	
äddar	s->1	
äddat	s->1	
ädde 	A->1	i->5	v->1	
äddni	n->4	
äde -	 ->1	
äde a	t->1	
äde e	n->1	
äde f	r->1	
äde h	a->1	
äde i	 ->1	
äde k	a->1	
äde m	e->1	
äde o	c->3	
äde t	i->4	
äde.H	a->1	
äde.J	a->2	
ädeHe	r->1	
ädePr	o->1	
ädels	e->6	
äden 	i->1	v->1	ä->1	
ädena	 ->1	
äder 	-->1	a->1	d->1	e->1	h->1	i->9	j->1	m->11	o->6	s->6	t->1	u->1	v->1	
äder,	 ->3	
äder.	S->1	
ädera	r->1	
äderi	,->1	n->2	
ädern	a->7	e->1	
äders	t->1	
ädes 	o->1	
ädes,	 ->1	
ädesp	e->7	
ädesv	i->2	
ädet 	a->4	d->1	h->1	i->2	o->1	t->1	
ädet,	 ->1	
ädet.	F->1	
ädja 	m->1	o->2	s->1	t->2	
ädjan	 ->1	d->3	
ädjar	 ->6	
ädjas	 ->1	
ädje 	-->1	a->1	f->1	k->1	n->1	ö->2	
ädret	 ->1	
äds a	v->1	
äds d	ä->1	
äds i	 ->1	
äds m	e->1	
äds r	å->1	
äds å	t->2	
äds ö	v->1	
ädsla	 ->4	,->1	.->1	n->3	
äer; 	e->1	
äffa 	d->1	e->1	i->1	o->1	u->1	
äffa,	 ->2	
äffa.	M->1	
äffad	e->6	
äffan	d->41	
äffar	 ->34	,->4	.->9	:->1	?->1	
äffas	 ->1	.->1	
äffat	 ->5	.->3	s->1	
äffli	g->2	
äfta 	a->5	d->2	f->1	h->1	o->1	v->1	
äfta,	 ->1	
äftad	e->3	
äftar	 ->3	
äftas	 ->4	.->1	
äftat	 ->5	s->2	
äftel	s->1	
äftig	a->1	
äg [K	O->1	
äg an	m->1	
äg at	t->6	
äg av	 ->1	
äg bo	r->1	
äg el	l->6	
äg fä	l->1	
äg fö	r->1	
äg ge	n->2	
äg hi	t->1	
äg hä	v->1	
äg i 	s->1	
äg in	n->1	
äg ku	n->1	
äg me	n->1	
äg mi	g->1	
äg mo	t->1	
äg oc	h->2	
äg si	n->1	
äg tr	ä->1	
äg är	 ->1	
äg ås	t->1	
äg, e	f->1	
äg, f	a->1	
äg, g	u->1	
äg, j	ä->6	
äg, o	c->1	
äg, p	å->1	
äg, s	o->3	å->1	
äg, v	i->1	
äg.Al	l->1	
äg.Bi	l->1	
äg.De	t->1	
äg.Ef	t->1	
äg.Ja	g->1	
äg.Me	n->1	
äg.Mi	n->1	
äg.Oa	v->1	
äg.Va	d->1	
äg: D	e->1	
ägNäs	t->1	
äga "	i->1	
äga -	 ->1	
äga F	r->1	
äga S	a->1	v->1	
äga a	n->1	t->79	
äga b	e->1	i->1	
äga d	e->13	
äga e	f->1	l->1	n->2	r->1	t->1	
äga f	ö->5	
äga g	e->1	
äga h	e->2	u->4	
äga i	 ->3	n->2	
äga j	a->1	
äga k	o->2	
äga l	i->2	ä->1	
äga m	e->1	
äga n	e->1	ä->3	å->7	
äga o	c->2	f->1	m->5	s->1	
äga r	e->1	u->18	
äga s	e->1	k->1	o->1	
äga t	i->8	
äga v	a->1	e->1	
äga ä	n->1	r->1	
äga å	t->1	
äga, 	a->1	d->1	e->1	f->1	h->4	i->1	k->1	l->1	o->2	u->1	v->1	å->1	
äga.D	e->1	
äga.J	a->1	
äga.M	e->1	
äga: 	"->1	D->1	F->1	d->1	
ägagå	n->6	
ägand	e->13	
ägar 	(->2	e->1	f->1	o->1	s->1	ä->1	
ägar,	 ->6	
ägar.	F->2	H->1	J->1	V->1	
ägara	n->1	
ägare	 ->2	!->1	,->1	.->2	?->1	n->11	
ägarn	a->6	
ägas 	a->2	t->1	v->1	
ägas,	 ->1	
ägbyg	g->1	
ägd g	e->1	
ägd l	ö->1	
ägda 	t->1	
ägde 	"->1	
äge d	ä->1	å->1	
äge g	e->1	
äge m	e->2	
äge s	n->1	o->2	
äge ä	r->1	
äge, 	b->1	
äge.H	e->1	
äge.V	å->1	
ägels	e->8	
ägen 	f->4	m->3	o->5	t->1	ä->1	ö->1	
ägen,	 ->3	
ägen.	H->1	
ägen:	 ->1	
ägenh	e->12	
äger 	1->1	E->1	a->27	d->3	e->5	f->1	h->1	i->5	j->10	k->2	l->2	m->3	n->6	o->1	p->1	r->2	s->1	t->5	ä->1	
äger,	 ->4	
äger.	F->1	O->1	
äger:	 ->5	
ägeri	 ->5	,->5	-->1	.->1	b->4	e->17	k->1	l->1	m->1	
ägesb	e->1	
ägesr	a->2	
äget 	a->4	f->2	i->3	m->2	o->1	s->1	ä->3	
äget,	 ->1	
äget.	J->2	
ägg d	ä->1	
ägg f	r->1	
ägg g	e->1	
ägg h	a->2	
ägg i	 ->3	n->1	
ägg k	u->1	
ägg l	å->1	
ägg m	ä->1	
ägg s	o->1	
ägg t	i->4	
ägg u	n->2	p->1	t->1	
ägg v	i->1	
ägg" 	s->1	
ägg, 	e->1	
ägg.F	ö->1	
ägga 	I->1	a->7	d->2	e->4	f->46	g->1	i->2	k->2	m->1	n->3	o->2	p->1	r->1	s->5	t->7	u->4	v->2	ö->1	
ägga,	 ->1	
äggan	d->76	
äggas	 ->8	,->2	.->1	
äggen	 ->2	
ägger	 ->39	
ägget	 ->1	,->1	
äggig	t->3	
äggni	n->27	
äggs 	f->7	i->3	n->1	p->4	u->1	v->1	
äggs,	 ->1	
äggsb	u->1	
äggsf	r->1	
äggsk	r->1	
äglad	 ->1	e->3	
äglas	 ->1	
ägled	a->3	n->2	
äglig	 ->1	t->1	
ägmär	k->1	
ägna 	a->1	g->1	i->1	l->1	m->1	o->3	r->1	s->6	t->1	
ägna,	 ->2	
ägnar	 ->22	,->3	.->4	
ägnas	 ->2	
ägnat	 ->3	s->1	
ägner	.->1	
ägnin	g->2	
ägra 	d->1	e->2	l->1	
ägrad	,->1	e->3	
ägran	 ->5	
ägrar	 ->4	
ägras	 ->1	
ägrat	 ->3	s->1	
ägre 	B->1	e->1	k->1	m->1	n->2	p->1	ä->1	
ägre.	S->1	Ä->1	
ägren	s->1	
ägröj	a->1	
ägs d	e->2	
ägs e	m->1	
ägs g	e->1	
ägs h	ä->1	
ägs i	g->1	n->1	
ägsen	 ->2	
ägset	 ->4	
ägskä	l->2	
ägsna	 ->4	,->1	
ägsnä	t->2	
ägsom	r->1	
ägsta	 ->1	
ägt d	e->1	
ägt f	r->1	
ägt r	u->9	
äkare	 ->1	,->2	u->1	
äkark	o->2	
äkeme	d->1	
äkens	k->9	
äker 	p->19	r->1	
äker,	 ->1	
äker.	P->1	
äkerh	e->235	
äkerl	i->15	
äkers	t->24	
äkert	 ->24	!->1	,->2	h->1	
äkna 	d->1	i->1	m->4	u->3	
äknad	e->1	
äknar	 ->21	
äknas	 ->4	
äknat	 ->3	s->2	
äknee	x->1	
äknel	i->1	
äknin	g->14	
äkra 	a->1	e->12	g->1	h->1	i->1	k->1	m->1	o->4	p->5	s->3	ö->1	
äkrar	 ->2	e->2	
äkras	.->1	t->4	
äkrin	g->24	
äkt f	ö->7	
äkt.O	m->1	
äkta 	a->2	m->2	p->1	s->1	
äktad	e->1	
äktar	 ->1	e->3	n->1	
äkten	 ->2	s->1	
äkter	,->1	
äktet	 ->1	
äktig	a->2	
äktin	g->1	
äkts 	ö->1	
äktsa	n->3	
äktsb	a->1	
äktsf	ö->1	
äl - 	o->1	u->1	
äl 6,	 ->1	
äl Sh	e->1	
äl al	l->1	
äl at	t->6	
äl av	 ->3	v->1	
äl be	f->1	g->1	r->1	
äl bi	b->1	
äl de	n->1	t->5	
äl då	?->1	
äl ef	t->1	
äl ek	o->1	
äl en	 ->2	
äl fr	å->1	
äl fu	n->1	
äl fö	r->9	
äl ge	n->2	
äl gä	l->1	
äl ha	n->1	r->4	
äl hu	r->1	
äl hä	r->1	
äl i 	D->1	E->1	F->1	o->1	p->1	s->1	
äl in	 ->1	n->1	o->1	t->6	ö->1	
äl ka	n->2	
äl ku	n->1	
äl kv	i->1	
äl kä	n->1	
äl lä	t->1	
äl ma	r->1	
äl me	d->5	l->1	
äl mo	t->1	
äl my	c->1	
äl ni	 ->1	
äl oc	h->3	
äl of	ö->1	
äl på	 ->3	
äl re	d->2	k->1	
äl si	n->1	
äl sk	u->1	
äl so	m->12	
äl st	a->1	r->1	
äl ti	l->8	
äl un	d->1	
äl up	p->1	
äl ur	 ->3	
äl ut	a->1	f->2	t->1	v->1	
äl va	r->1	
äl ve	t->1	
äl vi	a->1	
äl vå	r->1	
äl än	d->2	
äl är	 ->3	
äl åt	e->1	
äl öv	e->1	
äl, i	n->1	
äl, k	u->1	
äl, m	e->2	
äl, o	c->1	
äl.Al	l->1	
äl.De	 ->1	
äl.Fr	u->1	
äl.Fö	r->2	
äl.Ja	g->2	
äl.Mi	n->1	
äl.Sa	m->1	
äla d	e->1	
äla v	i->1	
älan 	o->1	
älbes	t->1	
äld å	t->1	
älda 	s->1	
äldig	a->3	t->20	
äldre	 ->5	,->1	.->1	
älen 	f->1	t->2	
älen"	,->1	
älen.	H->1	
äler.	D->1	
äleri	 ->1	
älet 	a->1	m->1	s->1	t->4	ä->1	
älet,	 ->1	
älfte	n->3	
älfun	n->1	
älfär	d->8	
älgru	n->2	
älgör	a->1	
älhav	a->1	
älig 	g->1	
älja 	H->1	e->2	n->1	o->1	s->2	u->1	
äljar	b->1	e->7	n->5	
äljas	 ->1	
äljer	 ->5	
äljni	n->3	
älkli	n->1	
älkom	m->7	n->42	s->1	
älkän	d->2	t->1	
äll u	t->1	
äll ä	r->1	
äll, 	a->1	b->1	
äll.J	a->1	
äll.O	m->1	
äll?K	o->1	
älla 	P->1	a->16	b->2	d->15	e->9	f->10	h->2	i->2	k->5	l->1	m->4	n->1	o->3	p->2	r->4	s->6	t->4	u->5	v->1	å->1	
älla,	 ->1	
älla.	D->1	H->1	
älla:	F->1	
ällan	 ->2	d->52	
ällar	 ->1	e->4	n->1	
ällas	 ->17	,->2	.->1	
ällba	r->1	
älld 	a->1	b->1	p->2	t->1	
ällda	 ->11	,->4	.->6	s->2	
ällde	 ->21	s->8	
älldh	e->23	
älle 	-->1	a->17	d->1	f->4	h->1	i->2	k->1	m->1	n->1	o->3	s->2	u->1	ä->1	
älle,	 ->1	
älle.	J->1	
ällel	s->7	
ällen	 ->36	"->1	,->7	.->13	a->5	s->2	
äller	 ->401	,->3	.->1	
älles	 ->2	
ället	 ->70	,->3	.->11	:->1	s->3	
ällig	 ->6	a->7	h->24	t->19	
ällni	n->71	
ällor	 ->17	,->5	.->12	n->5	
älls 	a->2	h->1	i->5	p->2	s->2	t->2	u->3	å->1	
älls.	N->1	Y->1	
ällse	k->3	
ällsk	a->8	
ällsm	e->1	
ällso	m->1	
ällss	e->1	
ällsv	ä->1	
ällsy	n->2	
ällt 	1->1	a->2	d->1	f->2	k->1	m->1	n->1	o->2	s->1	t->1	u->1	ä->1	
ällt,	 ->1	
ällt.	V->1	
ällts	 ->8	:->1	
älmen	t->2	
älmåe	n->2	
älnin	g->12	
älp a	t->1	v->26	
älp d	e->1	
älp f	r->3	ö->3	
älp n	i->1	
älp o	c->2	
älp p	å->1	
älp s	k->1	o->1	
älp t	i->5	
älp v	i->2	
älp ö	v->1	
älp, 	d->1	m->1	
älp.D	e->1	
älp.H	ä->1	
älp.I	 ->1	
älp.J	a->1	
älp.V	i->1	
älpa 	W->1	a->1	d->5	f->2	g->1	h->1	i->1	k->2	l->1	m->8	o->3	p->1	s->2	t->7	v->1	
älpan	d->3	
älpar	e->1	
älpen	 ->4	
älper	 ->1	
älpli	g->1	
älps.	J->1	
älpt 	t->1	
älpta	.->1	
älpte	 ->1	
älpvi	l->1	
äls m	å->1	
äls t	i->1	
älsa 	k->1	o->11	p->1	s->1	t->1	
älsa,	 ->3	
älsa.	H->1	
älsan	 ->1	,->2	.->1	
älsar	 ->1	
älsig	n->1	
älska	 ->1	r->1	
älsni	n->2	
älso-	 ->1	
älsoe	f->1	
älsor	e->1	i->1	
älsos	k->1	
älsov	å->3	
älstr	u->1	
älstå	n->6	
ält a	r->1	
ält e	f->1	
ält i	n->1	
ält o	c->1	
ält p	å->1	
ält s	i->1	
ältal	i->2	
älte 	k->1	v->1	
älte,	 ->2	
älten	.->1	a->1	
ältet	 ->5	"->1	.->3	
ältni	n->1	
ältsi	t->1	
älutb	i->1	
älutv	e->2	
älv a	n->1	r->1	t->3	
älv b	e->1	i->1	
älv f	r->2	ö->3	
älv g	o->1	
älv h	a->2	ö->1	
älv i	 ->3	
älv k	o->1	
älv m	e->1	
älv o	c->3	
älv s	a->1	e->1	k->1	o->3	ä->1	
älv t	a->1	
älv u	n->1	t->1	
älv v	a->1	e->1	
älv ä	r->3	
älv, 	h->3	m->2	
älv.D	e->1	
älv.J	a->1	
älv.K	o->1	
älv.V	i->1	
älva 	E->1	a->1	b->5	d->3	f->1	h->1	i->1	k->6	l->1	m->1	o->4	r->1	s->5	t->1	u->1	v->26	ä->2	
älva,	 ->3	
älva.	D->1	L->1	N->1	O->1	V->1	
älvan	d->1	
älvbe	s->3	
älvbi	o->1	
älvbä	r->1	
älvfa	l->2	
älvfö	r->1	
älvhj	ä->1	
älvkl	a->20	
älvko	s->1	
älvni	n->3	
älvpl	å->1	
älvst	y->7	ä->8	
älvsä	k->1	
älvt 	d->1	h->2	k->1	s->1	
älvän	d->1	
ämbet	e->5	s->3	
ämd a	t->1	
ämd h	ö->1	
ämd i	n->1	
ämd o	m->1	
ämd t	i->1	
ämd v	i->1	
ämda 	a->1	m->1	o->1	r->1	v->1	å->3	
ämda,	 ->1	
ämde 	T->1	i->1	m->2	s->1	
ämdhe	t->1	
ämels	e->1	
ämför	 ->3	b->4	e->2	t->9	
ämja 	a->2	d->4	e->8	f->3	g->2	h->1	i->1	k->4	l->2	p->1	s->4	v->1	y->1	å->2	
ämja.	K->1	
ämjan	d->17	
ämjar	 ->6	
ämjas	,->1	
ämjat	 ->1	
ämka 	i->1	
ämkar	 ->1	
ämlig	a->1	e->46	h->15	
ämlik	 ->1	h->12	
ämlin	g->34	
ämma 	a->1	d->1	i->6	k->1	m->5	o->1	p->1	v->1	ö->1	
ämma,	 ->1	
ämmad	 ->1	e->2	
ämman	d->10	
ämmar	 ->1	
ämmas	 ->2	,->1	
ämmel	s->122	
ämmer	 ->37	,->1	.->1	
ämmig	a->1	h->2	t->1	
ämn s	p->1	
ämn, 	f->1	
ämn.D	e->1	
ämna 	A->1	L->1	a->4	b->1	d->9	e->5	f->4	g->1	h->3	i->5	k->1	m->1	n->1	o->1	p->1	s->6	t->4	u->3	v->2	
ämna,	 ->1	
ämnad	 ->1	e->8	
ämnan	d->3	
ämnar	 ->19	e->4	
ämnas	 ->11	,->2	
ämnat	 ->13	s->5	
ämnda	 ->7	s->1	
ämnde	 ->11	,->4	.->2	s->1	
ämne 	h->1	i->1	s->1	
ämne.	D->2	
ämne:	 ->1	
ämnen	 ->11	,->2	.->5	a->1	
ämner	 ->4	.->1	
ämnet	 ->2	.->2	
ämnin	g->17	
ämns 	a->1	e->1	f->1	h->1	i->1	m->1	o->1	u->1	
ämns.	D->1	
ämnt 	b->1	e->1	f->1	g->1	i->1	k->1	l->1	n->1	p->1	
ämnt,	 ->2	
ämnt.	D->2	
ämnts	 ->2	,->2	.->2	
ämnvi	k->1	
ämnvä	r->1	
ämpa 	-->1	a->7	b->3	d->12	e->4	f->12	g->3	i->1	k->5	m->1	n->1	o->2	p->5	r->2	s->6	t->1	u->2	å->1	
ämpad	 ->1	
ämpan	d->3	
ämpar	 ->12	.->1	
ämpas	 ->32	,->1	.->8	:->1	
ämpat	 ->3	s->5	
ämpel	 ->1	
ämpli	g->60	n->1	
ämpni	n->80	
ämra 	e->1	k->1	
ämrad	 ->2	e->2	
ämran	d->1	
ämrar	 ->1	
ämras	 ->1	.->1	
ämre 	b->1	f->2	l->1	s->1	
äms u	t->1	
ämsid	e->1	
ämst 	I->1	a->2	d->2	e->2	g->2	i->5	k->3	l->3	m->1	o->3	p->2	s->1	t->2	u->2	v->7	ö->1	
ämst.	F->1	
ämsta	 ->13	
ämstä	l->24	
ämt a	l->1	t->3	
ämt e	n->1	
ämt f	a->1	r->1	
ämt i	 ->1	
ämt o	c->1	
ämt p	o->1	
ämt s	a->1	i->2	t->1	
ämt t	i->1	
ämt ö	k->1	v->1	
ämt, 	f->1	g->1	v->1	
ämt.D	e->1	
ämta 	s->2	u->1	
ämtan	d->1	
ämtar	 ->1	
ämtas	 ->1	
ämtat	 ->1	
ämtni	n->1	
ämtsa	m->1	
ämvik	t->2	
än 1 	p->2	
än 10	 ->1	0->2	
än 16	 ->1	
än 20	 ->1	
än 21	 ->1	
än 30	 ->2	
än Eu	r->1	
än Fo	l->1	
än Wa	l->1	
än ac	c->1	
än al	l->2	
än at	t->13	
än av	 ->1	
än ba	r->2	
än de	 ->4	b->2	m->1	n->8	t->5	
än di	r->1	t->1	
än ej	 ->1	
än el	l->1	
än en	 ->29	d->1	
än et	t->4	
än fa	r->2	
än fe	d->1	m->2	
än fr	a->1	
än fö	r->7	
än ge	n->2	
än gi	l->2	
än ha	r->3	
än hi	t->1	
än i 	a->2	d->5	e->1	f->2	h->1	l->1	p->1	v->1	
än in	f->1	g->1	s->1	
än ja	g->1	
än ka	n->2	
än ko	m->1	n->3	
än li	v->1	
än lo	g->1	
än lä	m->1	n->1	
än ma	g->1	n->4	
än me	d->2	
än mi	n->5	
än my	c->1	
än må	 ->1	
än na	t->1	
än nä	r->2	
än nå	g->6	
än oc	h->13	
än om	 ->1	d->1	r->1	
än p.	g->1	
än pe	r->1	
än po	l->1	
än på	 ->3	s->1	
än ra	m->2	
än re	a->2	e->1	l->1	
än sa	n->1	
än sk	a->2	
än so	m->10	
än st	a->2	o->1	
än sä	g->1	
än så	 ->4	:->1	h->1	
än ti	l->6	o->1	
än tr	e->2	
än tv	å->2	
än ut	a->1	s->1	
än va	d->7	
än vi	 ->2	,->1	.->1	k->1	l->1	s->1	
än vä	l->2	n->1	
än vå	r->1	
än är	 ->1	,->1	.->2	
än åk	l->6	
än år	 ->2	
än, e	t->1	
än, m	e->1	
än.In	t->1	
än.Ja	g->2	
än.Ty	v->1	
än; d	e->1	
äna a	n->1	
äna n	å->1	
äna r	ä->1	
äna s	i->1	o->1	t->2	
änade	 ->1	
änar 	a->3	d->3	f->1	i->3	s->1	t->2	v->1	
änar.	.->1	H->1	
änd (	e->1	
änd b	e->3	
änd e	r->1	
änd m	e->1	i->3	
änd, 	b->1	n->1	
änd.K	o->1	
ända 	1->1	E->1	a->5	b->1	d->15	e->6	f->9	g->2	h->1	i->8	j->2	m->4	n->1	o->3	p->4	r->2	s->11	t->5	u->2	v->1	ä->4	
ända,	 ->1	
ända.	D->1	F->1	N->1	V->2	
ända?	D->1	
ändam	å->13	
ändan	 ->3	,->1	.->1	d->2	o->1	
ändar	 ->1	e->5	n->3	
ändas	 ->11	,->1	.->4	
ändat	,->1	
ändba	r->9	
ände 	E->2	d->4	e->1	f->4	i->2	j->1	k->3	m->1	n->2	p->1	s->1	t->1	u->2	å->1	
ände,	 ->1	
ände.	D->1	
ändeb	u->9	
ändel	s->27	
änder	 ->114	"->1	,->21	.->25	?->2	l->1	n->79	s->6	
ändes	 ->10	,->1	
ändet	 ->1	
ändig	 ->25	,->2	.->3	a->36	h->48	t->118	
ändli	g->5	
ändlö	s->1	
ändni	n->64	
ändpu	n->6	
ändra	 ->36	,->1	d->8	r->5	s->13	t->12	
ändri	n->293	
änds 	a->1	d->1	f->5	i->2	m->3	o->1	p->6	v->1	
ändsk	 ->5	-->1	a->19	t->1	
ändå 	A->1	a->7	b->5	d->1	e->5	f->5	g->2	h->3	i->4	k->1	l->1	o->2	s->3	t->4	u->4	v->1	ä->2	
ändå,	 ->1	
ändå.	.->1	
änför	 ->1	
äng g	e->1	
äng k	o->2	
äng o	c->1	
äng å	t->1	
äng.D	e->1	
änga 	b->1	e->1	f->1	m->3	n->1	r->2	s->3	å->1	
änga,	 ->1	
ängan	d->3	
ängar	e->6	
ängas	 ->1	.->1	t->2	
ängbr	o->1	
ängd 	a->1	b->1	f->5	i->1	o->4	s->2	y->1	ä->1	å->1	
ängda	 ->1	
ängde	 ->2	n->5	r->5	
änge 	E->1	a->2	b->1	d->4	i->2	k->2	m->1	n->1	p->3	s->10	t->1	u->1	v->4	ä->1	å->1	
ängel	s->1	
änger	 ->18	
änges	f->1	
änget	t->1	
ängig	g->1	t->1	
ängil	t->1	
ängli	g->23	
ängni	n->44	
ängre	 ->55	,->1	.->6	
ängs 	e->1	k->1	
ängsl	i->1	
ängsy	s->2	
ängt 	a->1	f->1	m->1	s->3	
ängta	r->1	
ängte	r->8	
änhet	 ->5	,->1	.->6	e->35	
änien	 ->1	
äning	.->1	
änite	t->12	
änk b	a->1	
änk p	å->1	
änk t	i->1	
änka 	a->3	d->2	e->2	h->2	m->2	o->1	p->16	s->7	ö->2	
änka,	 ->1	
änkan	d->288	
änkas	 ->2	,->1	
änkba	r->4	
änken	 ->1	
änker	 ->41	
änkli	g->5	
änkni	n->15	
änks 	o->2	t->1	
änksa	m->2	
änkt 	a->2	g->1	h->1	s->1	
änkt.	V->1	
änkta	 ->6	,->1	.->1	
änkte	 ->3	
änkts	 ->3	
änlig	 ->2	a->8	e->1	t->4	
änna 	T->1	a->7	b->1	d->5	e->2	f->2	g->2	i->3	k->5	m->3	n->1	o->5	p->6	r->5	s->10	t->2	u->1	v->5	ä->1	å->2	
änna,	 ->1	
änna.	 ->1	U->1	
ännag	a->3	e->3	i->3	
ännan	d->26	
ännas	 ->6	,->1	.->1	
änne 	å->1	
änned	o->1	
ännel	i->1	
ännen	 ->21	,->1	.->2	s->4	
änner	 ->70	,->2	.->2	
ännet	e->6	
ännin	g->10	
ännis	k->98	
änns 	d->1	m->1	o->1	
änns.	E->1	
ännu 	a->1	e->11	f->1	h->5	i->32	m->8	n->1	p->1	s->9	v->2	ä->1	
ännu.	D->1	K->2	V->1	
ännu;	 ->1	
ännyt	t->2	
äns f	ö->1	
äns p	r->1	
äns s	i->2	
äns v	i->2	
änsa 	a->2	d->2	m->1	p->1	s->3	t->2	u->1	
änsa,	 ->1	
änsad	 ->13	,->1	.->3	e->10	
änsan	d->3	
änsar	 ->5	
änsas	 ->5	
änsat	 ->5	.->3	s->1	
änsch	 ->1	?->1	
änsee	n->8	
änsen	 ->3	.->1	
änser	 ->12	,->1	.->2	?->3	n->12	
änsfr	å->2	
änska	p->1	
änskl	i->42	
änsko	n->7	
änsla	 ->13	"->1	,->1	
änsle	n->2	s->5	
änsli	g->21	
änslo	l->1	m->1	r->5	
änsni	n->12	
änsom	r->1	
änspr	o->1	
änst 	i->2	o->2	s->1	å->1	
änst,	 ->1	
änst.	J->2	
änste	e->5	f->6	l->1	m->39	n->4	p->1	r->66	s->2	
änstf	u->1	
änstg	ö->3	
änstr	a->1	
änsvä	r->1	
änsyn	 ->67	;->1	e->2	s->2	
änsöv	e->12	
änt -	 ->1	
änt a	n->2	t->3	v->3	
änt d	e->3	
änt e	n->1	t->1	x->2	
änt f	a->1	ö->1	
änt g	ä->1	
änt h	å->1	
änt i	n->3	
änt k	ä->1	
änt l	ö->1	
änt m	a->1	e->1	i->1	å->2	
änt o	m->1	
änt p	l->1	r->1	
änt s	e->3	i->2	o->1	t->1	v->1	ä->1	
änt t	a->1	i->1	v->1	
änt u	n->3	r->1	t->1	
änt, 	l->1	m->1	u->1	
änt.J	a->1	
änt.V	i->1	
änt: 	U->1	
änta 	a->2	b->4	e->2	f->22	i->1	m->2	o->1	p->4	r->1	s->1	t->3	
änta.	 ->1	D->1	
äntad	e->1	
äntan	 ->4	.->1	
äntar	 ->38	.->1	
äntas	 ->2	
äntat	 ->4	.->1	
äntli	g->20	
äntni	n->7	
änts 	a->5	e->1	f->1	i->2	m->2	p->1	v->1	
änvis	a->25	n->10	
äpade	s->1	
äpnad	e->2	
äpnin	g->1	
äpp a	v->1	
äpp k	a->1	
äpp, 	a->1	
äpp.D	e->1	
äppa 	e->1	i->3	t->3	
äppan	d->2	
äppen	 ->2	,->1	
äpper	 ->2	
äppet	 ->1	
äpphä	n->1	
äppsr	ä->1	
äppte	 ->1	s->2	
äprod	u->1	
är "k	r->1	
är - 	a->1	d->1	f->1	i->2	j->1	o->4	s->2	ö->1	
är 1,	2->1	
är 1/	3->1	
är 10	 ->1	0->1	
är 16	7->1	
är 25	 ->1	
är 29	 ->1	
är 30	 ->1	
är 50	 ->1	
är 7 	p->1	
är 80	 ->1	
är An	t->1	
är Ba	r->8	
är Bo	l->1	
är CE	N->1	
är Do	r->1	
är EU	 ->1	-->3	:->1	
är Eg	y->1	
är Eu	r->11	
är FN	.->1	
är FP	Ö->1	
är Ki	n->5	
är Lu	x->1	
är Ma	r->1	
är Mo	n->13	
är Ni	e->1	
är Pa	l->1	t->16	
är Po	m->1	r->1	
är Pr	e->1	
är Re	d->2	
är Sc	h->1	
är So	l->1	
är Vi	t->4	
är Wa	l->1	s->1	
är ab	s->10	
är ac	c->2	
är ak	t->5	
är al	l->45	
är am	b->1	
är an	a->1	d->2	g->7	l->3	m->1	n->1	o->1	s->22	t->1	v->1	
är ar	b->4	
är at	t->167	
är av	 ->21	g->7	h->1	l->1	s->10	
är ba	r->12	s->2	
är be	d->1	f->3	g->5	h->7	k->6	r->34	s->4	t->19	v->2	
är bl	a->1	i->2	
är bo	s->2	v->1	
är br	a->18	i->4	
är bu	d->1	
är by	g->1	
är bä	r->1	s->1	t->5	
är bå	d->5	
är bö	r->3	
är ce	n->2	
är ci	t->1	
är co	r->1	
är da	g->7	
är de	 ->56	,->1	b->7	f->2	l->1	m->1	n->74	r->1	s->15	t->421	
är di	r->4	s->2	
är dj	u->4	
är do	c->16	m->2	
är dr	i->1	o->1	
är dä	r->29	
är då	 ->2	l->3	
är dö	d->1	
är ef	f->3	t->1	
är eg	e->6	
är ek	o->1	
är el	l->1	
är em	e->10	o->2	
är en	 ->215	b->2	d->4	g->2	h->2	k->3	l->10	o->2	s->3	
är er	a->1	
är et	a->3	t->120	
är eu	r->1	
är ev	i->1	
är ex	c->1	e->2	p->3	
är fa	k->5	l->19	r->3	s->3	
är fe	l->6	m->1	
är fi	n->10	
är fl	e->1	i->1	o->2	
är fo	l->1	n->1	r->14	
är fr	a->5	e->3	u->1	ä->2	å->35	
är fu	l->11	
är fy	l->1	
är fä	r->1	
är få	,->1	
är fö	g->1	l->3	r->96	
är ga	n->6	r->1	
är ge	m->5	n->5	r->1	
är gi	v->2	
är gj	o->2	
är gl	a->12	ä->1	
är go	d->8	
är gr	u->7	
är gå	 ->1	n->3	r->1	
är ha	l->2	n->16	r->16	v->1	
är he	d->1	l->31	
är hi	s->1	t->1	
är hj	ä->1	
är ho	m->1	n->1	r->1	t->2	
är hu	r->5	v->1	
är hä	n->1	r->3	
är hå	l->1	r->1	
är hö	g->1	
är i 	2->1	E->6	I->1	S->1	a->5	b->1	d->20	e->2	f->5	g->3	h->1	k->9	m->1	n->1	o->1	p->14	r->2	s->8	t->2	u->1	v->2	å->1	ö->1	
är ib	l->2	
är id	e->1	é->1	
är il	l->1	
är in	 ->1	c->1	f->3	g->17	k->1	l->2	n->2	o->2	r->2	s->4	t->117	v->4	
är is	r->1	
är ja	g->51	
är ju	 ->11	,->1	r->2	s->4	
är jä	m->1	
är ka	m->1	n->9	t->3	
är kl	a->13	o->1	
är kn	a->2	u->3	
är ko	a->1	l->1	m->37	n->14	r->4	s->1	
är kr	a->1	i->1	ä->1	
är ku	l->1	
är kv	a->1	ä->1	
är kä	n->6	r->1	
är la	g->5	n->1	
är le	d->4	g->2	
är li	g->1	k->12	s->1	t->7	
är lo	g->1	k->1	
är ly	c->2	
är lä	g->1	m->9	n->1	t->5	
är lå	n->6	
är lö	j->2	s->2	
är ma	n->47	s->1	
är me	d->34	n->5	r->9	s->2	
är mi	l->2	n->8	s->1	t->4	
är mo	d->1	t->3	
är mu	n->1	
är my	c->56	
är mä	n->2	
är må	l->2	n->4	s->4	
är mö	j->21	
är na	t->18	
är ne	g->1	j->1	r->3	
är ni	 ->6	,->2	
är no	g->1	r->1	
är nu	 ->10	:->1	
är ny	 ->1	a->3	c->1	t->1	
är nä	m->1	r->10	s->2	
är nå	g->29	
är nö	d->30	j->4	
är oa	c->5	
är ob	e->4	
är oc	h->16	k->39	
är oe	n->1	r->6	t->1	
är of	f->4	t->1	u->1	ö->4	
är oj	ä->1	
är ok	l->2	
är ol	i->1	j->1	y->2	
är om	 ->5	f->2	r->5	ö->3	
är on	ö->1	
är or	d->1	o->2	s->1	ä->2	
är os	ä->1	å->1	
är ot	i->3	
är ou	m->1	n->1	t->1	
är pa	r->7	
är pe	n->1	r->2	
är pl	a->5	e->1	
är po	l->4	s->5	ä->1	
är pr	e->9	i->3	o->10	
är pu	n->2	
är på	 ->17	b->1	
är re	a->1	d->7	f->1	g->7	l->3	n->1	p->3	s->3	t->1	v->1	
är ri	k->8	m->3	n->1	
är ro	l->1	s->1	
är ru	i->1	n->1	s->1	
är rä	d->2	k->1	t->10	
är rå	d->2	
är rö	r->1	
är sa	k->2	m->6	n->8	
är se	d->1	r->2	x->1	
är si	s->1	t->4	
är sj	u->1	ä->7	ö->1	
är sk	a->4	i->2	r->2	u->2	y->6	ä->3	ö->1	
är sl	a->2	u->1	
är sn	a->3	
är so	c->1	m->16	
är sp	a->3	e->2	ä->1	
är st	a->5	o->9	r->4	å->1	ö->4	
är su	b->1	n->1	
är sv	a->1	å->10	
är sy	f->3	n->3	s->1	
är sä	k->18	m->1	n->1	r->25	t->1	
är så	 ->15	,->1	d->1	l->9	v->1	
är ta	c->1	r->1	
är te	k->2	m->1	x->2	
är ti	d->1	l->38	t->1	
är tj	ä->2	
är to	r->1	t->1	
är tr	a->1	e->1	o->2	å->1	ö->1	
är tv	i->1	å->9	
är ty	d->8	p->11	v->2	
är tä	n->3	
är un	d->4	g->2	i->4	
är up	p->23	
är ur	s->1	
är ut	a->9	e->4	i->1	o->3	p->1	r->2	s->2	t->2	v->2	
är va	d->9	k->2	r->1	t->1	
är ve	c->2	r->12	t->3	
är vi	 ->99	k->50	l->9	s->2	t->1	
är vu	n->1	
är vä	g->1	l->18	r->11	s->2	
är vå	r->10	
är yp	p->1	
är yr	k->1	
är yt	t->10	
är Ös	t->1	
är äg	n->1	
är äl	d->2	
är än	 ->1	d->6	g->1	n->4	
är är	 ->14	l->1	
är äv	e->4	
är år	e->2	
är åt	e->3	
är öd	e->1	
är ök	a->1	
är ön	s->2	
är öp	p->3	
är öv	e->29	r->1	
är! 1	9->1	
är! B	e->1	
är! C	e->1	
är! D	e->2	
är! E	f->2	t->1	
är! F	ö->1	
är! I	 ->2	
är! J	a->6	
är! L	å->2	
är! N	i->1	ä->1	
är! O	m->1	
är! T	a->1	
är! U	n->1	
är! V	i->4	
är! Ä	v->1	
är!.H	e->1	
är!De	t->1	
är!Er	i->1	
är!Ja	g->1	
är, a	l->1	n->1	t->11	
är, b	ä->3	
är, d	e->2	å->1	
är, f	r->1	å->1	ö->7	
är, h	e->5	ä->1	
är, i	 ->3	n->1	
är, j	a->3	
är, k	o->2	ä->12	
är, l	ä->1	
är, m	e->8	i->6	å->1	
är, n	a->1	i->1	ä->2	
är, o	c->5	m->3	r->1	
är, p	å->1	
är, r	ä->1	
är, s	a->1	o->2	v->1	å->1	
är, t	i->1	y->2	
är, u	n->1	p->1	
är, v	e->1	i->5	ä->3	
är, ä	r->10	
är. D	e->1	
är. N	i->1	
är. i	n->1	
är.. 	(->1	
är.De	 ->2	n->2	t->5	
är.Dä	r->1	
är.Ef	t->1	
är.En	 ->1	
är.Fö	r->4	
är.Ge	m->1	
är.He	r->1	
är.I 	e->1	
är.Ja	g->11	
är.Ko	m->1	
är.Ra	s->1	
är.So	m->2	
är.Så	l->1	
är.Va	d->1	
är.Vi	 ->7	
är.ko	m->1	
är: F	ö->1	
är: h	u->1	
är: n	u->1	
är: v	e->1	
är: Ä	r->1	
är; v	i->1	
är?De	t->1	
är?Ha	r->1	
är?Ja	g->1	
ära 5	 ->1	
ära a	n->2	t->12	
ära b	e->2	
ära d	e->2	i->1	
ära e	k->1	n->3	t->1	
ära f	a->2	r->5	ö->4	
ära h	e->3	u->1	å->1	
ära i	g->1	
ära k	o->56	r->1	u->2	
ära l	e->2	
ära m	a->1	e->3	
ära o	c->3	r->3	s->1	
ära p	a->1	e->1	l->1	
ära r	a->1	
ära s	a->5	i->4	k->1	l->1	t->2	
ära u	n->5	
ära ä	n->1	r->1	
ära å	t->1	
ära, 	o->1	s->1	
ära.N	ä->1	
ärade	 ->22	
äran 	a->5	f->3	g->1	i->1	j->1	m->1	o->5	s->1	
äran,	 ->3	
äran.	)->1	F->1	N->1	
äran?	F->1	
ärand	e->3	
ärare	 ->1	n->1	
ärart	,->1	
äras 	a->1	f->3	g->1	h->1	
ärav 	d->1	f->1	s->1	v->1	
ärbes	t->1	
ärd 2	 ->1	
ärd a	t->2	v->2	
ärd b	r->1	
ärd d	e->1	ä->1	
ärd e	k->1	l->1	n->1	
ärd f	ö->2	
ärd k	o->1	
ärd m	a->1	e->1	i->1	
ärd o	c->4	
ärd s	i->1	o->2	
ärd u	r->1	
ärd v	i->2	
ärd, 	b->1	d->1	h->1	m->1	s->1	t->2	ä->1	
ärd.D	e->3	
ärd.H	e->1	
ärd.I	 ->1	
ärd.J	a->1	
ärd; 	d->1	i->1	
ärda 	a->2	d->1	e->3	f->1	g->1	h->2	k->2	n->1	o->1	p->1	r->1	s->3	t->2	v->1	ä->1	
ärda,	 ->2	
ärda.	O->1	
ärdan	d->5	
ärdar	 ->2	
ärdas	 ->1	.->1	
ärdat	 ->2	
ärde 	a->1	d->3	f->1	m->1	o->2	p->5	r->1	s->3	u->1	
ärde,	 ->1	
ärde-	 ->1	
ärde.	D->1	G->1	J->1	T->1	
ärded	e->2	
ärdef	u->7	
ärdeg	e->3	
ärdel	ö->1	
ärden	 ->9	,->3	.->3	a->4	s->1	
ärder	 ->151	,->13	.->20	?->1	a->19	i->43	n->21	
ärdes	s->2	
ärdet	 ->4	
ärdig	 ->6	.->1	a->11	h->18	s->1	t->4	
ärdli	g->3	
ärdom	 ->6	,->1	
ärds 	r->1	
ärdsb	u->1	
ärdsl	i->1	
ärdsm	å->1	
ärdso	m->1	
ärdsp	a->2	l->3	r->1	u->1	
ärdss	k->1	t->2	
ärdsv	i->1	
äre k	o->1	
äreft	e->12	
äremo	t->19	
ären 	-->2	a->1	b->1	f->7	g->1	h->1	i->5	j->1	m->2	n->1	o->8	p->2	s->5	u->1	v->2	ä->1	
ären,	 ->6	
ären.	J->1	V->1	
ären?	V->1	
ärend	e->21	
ärens	 ->3	
ärer 	b->1	e->1	f->1	h->1	i->1	m->1	o->5	s->3	
ärer!	 ->1	
ärer,	 ->5	
ärer.	D->1	
ärern	a->14	
äret 	a->1	
ärfrå	g->1	
ärför	 ->271	,->7	.->1	:->1	
ärg, 	k->1	s->1	
ärgad	 ->1	
ärhet	 ->1	e->4	
ärhän	;->1	
äri s	e->1	
äri v	a->1	
äribl	a->6	
ärifr	å->2	
ärige	n->19	
äring	s->12	
ärjad	e->2	
ärka 	-->2	2->1	E->1	a->2	d->5	i->1	k->3	m->1	p->1	r->1	s->2	t->3	u->1	v->2	
ärka,	 ->1	
ärkan	d->2	
ärkas	 ->2	.->1	
ärkba	r->3	
ärke 	i->2	t->5	
ärkel	s->5	
ärken	 ->2	
ärker	 ->7	
ärket	,->1	
ärkil	t->1	
ärkli	g->5	
ärkni	n->19	
ärks 	b->1	g->1	o->1	
ärks.	D->1	O->1	V->1	
ärksa	m->53	
ärkt 	E->2	a->3	b->3	c->1	d->1	e->1	i->2	k->1	o->2	p->1	r->2	s->2	
ärkt.	D->1	
ärkta	 ->18	
ärkts	 ->1	
ärl o	c->1	
ärld 	s->1	
ärld,	 ->2	
ärld.	J->1	
ärlde	n->37	
ärlds	d->1	e->1	f->1	h->4	k->6	l->1	m->1	n->1	o->1	
ärled	a->1	
ärlek	e->2	
ärlig	 ->3	!->1	,->1	.->1	a->9	t->5	
ärlin	g->1	
ärma 	s->1	v->1	
ärman	d->1	
ärmar	 ->5	e->15	
ärmas	t->13	
ärmed	 ->47	,->2	
ärmel	s->1	
ärmin	i->10	
ärmni	n->5	
ärn- 	o->2	
ärna 	b->1	f->1	g->3	h->3	k->3	m->1	o->2	s->5	t->3	u->3	v->9	
ärna.	F->1	
ärnan	 ->6	
ärnar	 ->1	
ärnen	e->8	
ärnfr	å->2	
ärnin	g->4	
ärnka	t->1	
ärnkr	a->22	
ärnpr	i->2	
ärnpu	n->2	
ärnst	r->1	
ärnsä	k->3	
ärnte	k->2	n->1	
ärnva	p->8	
ärnvä	g->15	
äro t	r->1	
äroan	s->1	
ärom 	d->1	
ärosa	t->1	
ärpa 	a->1	b->1	d->1	h->1	k->1	t->1	
ärpas	 ->1	?->1	
ärper	s->1	
ärpla	n->1	
ärpni	n->1	
ärpol	i->2	
ärpta	 ->2	
ärpå 	k->1	t->1	
ärr a	l->1	
ärr b	a->1	l->1	ö->1	
ärr d	e->3	
ärr f	i->1	o->1	ö->1	
ärr g	ö->1	
ärr h	a->6	
ärr i	n->4	
ärr k	a->2	o->1	
ärr n	ä->1	
ärr o	c->1	f->1	
ärr s	a->1	e->1	t->1	ä->1	
ärr ä	n->1	r->3	v->1	
ärr å	t->1	
ärr, 	i->1	ä->1	
ärr.V	i->1	
ärra 	p->1	
ärrar	.->1	;->1	
ärras	 ->1	,->1	
ärrat	s->1	
ärre 	a->1	i->1	k->1	m->1	o->1	s->2	ä->1	
ärre,	 ->1	
ärrät	t->1	
ärrör	 ->4	
ärs f	r->1	ö->1	
ärs h	a->1	
ärs m	o->1	
ärs n	e->1	
ärs s	å->1	
ärski	l->158	
ärskt	 ->1	
ärsmä	n->1	
ärst 	j->1	
ärsta	 ->7	
ärsyn	t->1	
ärt F	P->1	
ärt a	r->1	t->11	
ärt b	i->1	
ärt e	l->1	m->1	n->3	
ärt f	r->1	
ärt g	e->1	
ärt i	n->1	
ärt k	r->1	
ärt m	e->1	y->1	
ärt o	r->2	s->1	
ärt p	å->1	
ärt s	i->1	k->1	
ärt, 	h->1	o->1	s->1	t->1	v->1	
ärt.J	a->1	
ärt.O	c->1	
ärt.S	l->1	
ärt.V	i->1	
ärta 	m->1	r->1	s->1	
ärtad	 ->1	
ärtan	s->2	
ärtar	 ->1	
ärtat	 ->10	,->1	.->2	:->1	
ärtil	l->2	
ärtli	g->7	
ärtom	 ->12	!->1	,->3	.->1	
ärtsa	m->1	
ärutö	v->1	
ärv o	c->1	
ärva 	d->1	f->1	n->1	o->1	p->1	r->1	
ärvad	e->1	
ärvar	a->42	e->1	o->4	
ärvat	 ->1	
ärvbr	i->1	
ärvhe	t->1	
ärvid	 ->5	l->1	
ärvli	g->1	
ärvsa	r->3	
ärvt 	p->2	
äs te	x->1	
äs un	d->1	
äs yt	t->1	
äsa k	o->1	
äsa o	m->1	
äsa v	a->1	
äsbar	 ->1	a->1	
äsch 	i->1	
äsche	n->1	
äsduk	a->1	
äsen 	a->1	f->1	
äsen,	 ->2	
äsend	e->6	
äsent	l->26	
äser 	b->1	d->4	k->1	
äsfrä	m->1	
äsk.H	e->1	
äskun	n->1	
äsnin	g->2	
äsong	s->1	
ässig	 ->3	a->15	t->13	
äst D	a->1	
äst a	t->1	
äst d	e->2	
äst e	n->1	t->1	
äst f	r->1	
äst g	e->1	
äst k	a->1	
äst r	e->1	
äst s	t->1	
äst t	i->1	
ästa 	b->2	d->2	e->3	f->4	g->4	k->6	l->1	m->9	n->1	o->2	p->27	r->13	s->16	t->2	u->3	v->1	å->1	
ästa.	D->1	H->1	V->2	
ästan	 ->16	.->1	d->2	
ästar	e->1	i->1	
ästba	n->4	
äste 	b->1	u->1	v->1	
ästel	s->1	
ästen	.->1	
äster	 ->8	
ästes	 ->1	
ästku	s->1	
ästma	k->1	
ästni	n->2	
ästra	 ->3	
ästs 	v->1	
ästvä	r->1	
ät dä	r->1	
ät ka	n->1	
ät mi	g->1	
ät oc	h->1	
ät os	v->1	
ät si	g->1	
ät sk	u->1	ä->1	
ät so	m->2	
ät. D	e->1	
äta d	e->1	
äta s	i->1	
äta, 	f->1	
ätare	 ->2	
ätas 	d->1	u->1	
äte.O	m->1	
äten 	f->3	m->1	
äter 	f->1	h->1	
ätet 	o->2	
äthet	e->1	
ätigt	 ->1	
ätor 	f->1	
ätska	 ->1	
ätstr	u->1	
ätt (	5->1	9->1	
ätt -	 ->2	
ätt H	a->1	
ätt a	l->1	n->3	t->51	
ätt b	e->7	o->1	ö->1	
ätt e	l->3	n->1	r->1	t->2	
ätt f	a->1	i->1	å->1	ö->15	
ätt g	e->5	r->1	ö->1	
ätt h	a->2	j->1	o->1	u->1	ä->1	å->2	
ätt i	 ->12	.->1	n->4	r->1	
ätt k	a->12	o->7	r->1	ä->1	ö->2	
ätt l	e->1	ä->1	ö->1	
ätt m	a->2	e->1	i->1	å->1	
ätt n	a->1	i->2	ä->1	
ätt o	c->22	m->1	s->1	
ätt p	l->1	o->1	å->7	
ätt r	i->6	
ätt s	a->2	e->1	i->2	k->6	o->28	t->3	ä->4	å->1	
ätt t	i->21	ä->1	
ätt u	n->5	r->1	t->2	
ätt v	a->2	e->1	i->6	ä->2	
ätt ä	n->2	r->7	v->1	
ätt å	t->2	
ätt ö	g->1	v->1	
ätt, 	a->2	b->1	d->1	e->4	f->1	g->1	h->4	i->1	k->1	m->3	n->1	o->7	p->1	s->5	t->1	v->2	ä->1	
ätt. 	D->2	
ätt.A	l->2	
ätt.B	e->1	
ätt.D	e->12	ä->1	
ätt.E	n->2	r->1	
ätt.F	ö->2	
ätt.H	e->6	
ätt.I	 ->1	
ätt.J	a->7	
ätt.K	o->2	
ätt.L	å->1	
ätt.M	a->1	e->3	i->1	
ätt.N	a->1	ä->1	
ätt.S	l->1	o->1	t->1	y->1	
ätt.V	i->5	
ätt.Ä	v->1	
ätt: 	"->1	j->1	
ätt?A	n->1	
ätt?D	e->1	
ätt?O	m->1	
ätt?S	k->1	
ätta 	E->1	a->19	b->1	d->22	e->31	f->11	g->2	h->1	i->8	k->1	l->2	m->16	n->3	o->5	p->9	r->2	s->20	t->4	u->3	v->2	å->2	ö->2	
ätta!	D->1	
ätta,	 ->4	
ätta.	D->1	H->1	V->1	
ättad	 ->1	e->8	
ättan	d->24	
ättar	 ->8	e->14	h->1	n->1	
ättas	 ->17	,->4	.->3	
ättat	 ->6	.->1	s->3	
ätte 	m->1	o->1	p->10	r->6	ö->2	
ätte,	 ->1	
ätted	e->1	
ätteg	å->1	
ättel	i->1	s->3	
ätten	 ->46	)->1	,->10	.->19	;->1	H->1	s->7	
ätter	 ->64	,->1	.->1	
ättes	 ->1	
ättet	 ->21	,->1	:->1	
ättfr	a->1	
ättfä	r->7	
ättfö	r->1	
ätthå	l->9	
ättig	a->19	h->103	
ättil	l->2	
ättli	g->1	
ättmä	t->1	
ättna	d->1	
ättni	n->213	
ättra	 ->42	d->5	n->1	r->4	s->6	t->2	
ättre	 ->66	,->3	.->6	
ättri	n->18	
ätts 	a->1	f->6	i->1	n->1	p->1	u->1	
ätts,	 ->2	
ätts.	D->1	
ättsa	k->4	
ättsf	ö->1	
ättsh	j->2	
ättsi	n->2	
ättsk	a->1	i->7	u->1	
ättsl	i->115	ä->3	
ättso	m->1	r->3	s->2	
ättsp	r->2	
ättsr	e->1	
ättss	e->1	k->3	t->9	y->20	ä->20	
ättst	i->2	j->1	r->1	
ättsv	ä->4	
ättvi	k->2	s->72	
ättän	k->1	
ätver	k->11	
äv me	d->1	
äva 4	0->1	
äva a	n->2	t->5	v->1	
äva d	e->2	u->2	
äva e	f->3	n->5	u->1	
äva f	a->1	i->1	ö->1	
äva i	 ->1	m->1	
äva j	u->1	
äva k	o->1	
äva m	e->2	
äva s	a->1	
äva t	e->1	i->2	
äva å	t->2	
äva ö	k->1	
ävade	 ->4	
ävan 	a->3	e->3	m->1	o->1	
ävan.	D->1	
ävand	e->7	
ävans	v->1	
ävar 	e->2	j->1	ä->1	
ävare	 ->1	
ävas 	a->3	e->3	f->1	i->1	o->3	
ävas,	 ->1	
ävas.	G->1	
ävat 	e->1	
ävda 	a->6	d->1	
ävdad	e->3	
ävdar	 ->10	,->1	.->1	
ävdat	 ->4	.->1	
ävde 	e->1	
ävde,	 ->1	
ävdes	 ->2	
ävdvu	n->1	
även 	-->1	E->2	G->1	R->2	a->16	b->3	d->18	e->10	f->19	g->2	h->5	i->41	j->3	k->9	l->3	m->12	n->9	o->62	p->7	r->3	s->10	t->11	u->7	v->5	y->1	ä->2	ö->2	
ävent	y->9	
äver 	a->14	d->2	e->9	i->1	j->2	k->3	m->2	n->4	o->2	p->1	s->1	v->2	y->1	
äver.	J->1	V->1	
äves 	h->1	
ävigt	,->1	
ävjas	 ->1	
ävlad	e->1	
ävlar	 ->1	
ävlin	g->1	
ävnad	 ->2	e->2	
ävnin	g->10	
ävs a	v->2	
ävs b	e->1	
ävs d	e->10	r->1	
ävs e	n->11	t->1	
ävs f	r->1	ö->7	
ävs h	a->1	
ävs i	 ->1	n->1	
ävs k	r->1	
ävs m	e->2	
ävs o	c->1	
ävs p	r->1	
ävs r	a->1	
ävs s	k->1	p->1	t->1	å->1	
ävs u	p->1	
ävs v	e->1	i->2	
ävs ä	r->1	
ävs, 	m->1	s->2	
ävs.E	t->2	
ävt e	n->1	
ävt s	i->1	
ävts 	ä->1	
ävts.	E->1	
ävule	n->1	
ävuls	k->1	
äxa u	t->1	
äxa.H	ä->1	
äxa.M	e->1	
äxan?	V->1	
äxand	e->6	
äxat 	u->1	
äxelk	u->1	
äxelv	e->2	
äxer 	d->1	f->1	o->2	s->2	
äxer,	 ->1	
äxlan	d->1	
äxlar	 ->1	
äxlin	g->2	
äxor.	D->1	
äxt a	v->1	
äxt o	c->4	
äxt s	o->1	
äxt ä	r->1	
äxt, 	i->1	s->1	
äxt.K	o->1	
äxt.O	c->1	
äxtbr	a->1	
äxten	 ->6	,->2	
äxter	 ->1	.->1	
äxthu	s->7	
äxtsk	y->3	
å "me	l->1	
å - a	t->1	
å - d	e->1	
å - i	n->1	
å - m	a->1	
å - o	c->2	m->1	
å - s	o->1	
å 10 	p->1	
å 100	 ->1	
å 13 	p->2	
å 140	 ->1	
å 199	9->1	
å 20 	p->1	
å 200	0->2	
å 22,	5->1	
å 24 	n->1	
å 33 	0->1	
å 34 	å->1	
å 37 	p->1	
å 40 	p->1	
å 5 m	i->1	
å 50 	p->1	
å 50-	 ->1	
å 7,2	 ->1	
å 75 	m->1	
å 80 	p->2	
å 86 	p->1	
å 90 	p->1	
å 95 	m->1	
å All	a->2	
å Ass	a->1	
å Atl	a->1	
å BSE	-->1	
å Bal	k->5	
å Bel	g->1	
å CEN	 ->1	
å CSU	-->1	
å Da 	C->1	
å EG-	d->2	k->1	r->1	
å EU-	n->1	r->1	
å EU:	s->2	
å Eri	k->2	
å Eur	o->18	
å Fla	u->1	
å För	e->1	
å Gen	e->1	
å Gol	a->2	
å Hol	l->1	
å ISP	A->1	
å Int	e->6	
å Irl	a->1	
å Isr	a->1	
å Kin	n->1	
å Mal	t->1	
å Mor	g->1	
å Oli	v->1	
å PPE	-->1	
å Pap	a->1	
å Ric	h->2	
å Roi	s->1	
å Tys	k->1	
å Väs	t->2	
å abs	o->1	
å acc	e->1	
å akt	a->1	i->2	u->1	
å alb	a->1	
å all	a->16	d->1	m->2	t->7	v->14	
å alt	e->1	
å amb	i->1	
å an 	a->1	
å and	r->22	
å ang	å->1	
å anl	e->1	
å anm	ä->1	
å ann	a->1	
å ans	e->2	j->1	l->1	t->1	v->4	å->1	
å ant	a->1	i->2	
å anv	ä->1	
å arb	e->9	
å arg	u->1	
å art	i->5	
å asp	e->2	
å asy	l->1	
å att	 ->353	
å av 	E->1	a->2	d->5	e->1	f->1	k->1	n->1	r->2	u->1	v->2	å->1	
å avf	a->1	
å avg	a->1	e->1	ö->2	
å avs	l->1	p->1	
å avt	a->1	
å bal	a->2	
å bar	 ->1	a->5	
å bas	i->2	k->1	
å be 	k->1	
å bef	a->2	o->2	
å beg	ä->1	
å beh	a->1	o->5	ä->1	ö->3	
å bek	l->1	o->1	r->1	y->1	
å ber	e->1	i->1	o->1	ä->1	
å bes	l->3	t->1	v->1	
å bet	r->1	y->6	ä->2	
å bid	r->1	
å bil	a->3	b->1	i->1	å->1	
å ble	v->1	
å bli	 ->2	r->6	
å blo	m->1	
å bly	g->1	
å bol	a->1	
å bor	d->5	g->1	t->2	
å bos	n->1	
å bra	 ->2	,->1	
å bre	d->4	t->1	
å bri	t->1	
å bro	m->1	t->2	
å byg	g->2	
å bär	 ->1	a->2	
å bäs	t->8	
å bät	t->2	
å båd	a->1	e->2	
å bör	 ->7	j->3	
å cen	t->1	
å civ	i->1	
å cri	c->1	
å dag	 ->1	a->1	e->2	o->5	
å dan	s->1	
å de 	2->1	a->6	b->1	c->1	e->3	f->8	h->4	i->3	j->1	k->2	m->7	n->6	o->5	p->1	r->4	s->8	t->1	u->4	v->1	å->1	ö->1	
å deb	a->2	
å def	i->2	
å del	a->2	t->2	v->2	
å dem	 ->5	.->1	o->3	
å den	 ->98	.->1	n->25	
å der	a->4	
å des	s->16	
å det	 ->92	,->1	.->2	?->1	a->2	t->68	
å dir	e->2	
å dis	k->2	
å dju	p->6	r->1	
å dom	s->2	
å dra	m->1	
å dru	n->1	
å dub	b->3	
å dum	p->1	
å dyl	i->1	
å där	 ->1	f->2	
å dål	i->1	
å eff	e->5	
å eft	e->2	
å ege	n->1	t->2	
å eko	n->5	s->1	
å ele	k->1	
å ell	e->3	
å emb	r->1	
å en 	a->14	b->7	c->1	d->4	e->6	f->6	g->7	h->9	i->1	j->1	k->6	l->9	m->13	n->2	o->5	p->2	r->5	s->10	t->6	u->3	v->7	ä->2	å->1	ö->3	
å ena	 ->11	d->1	
å end	a->1	
å eng	e->1	
å enh	e->1	ä->2	
å eni	g->1	
å enk	e->1	
å enl	i->2	
å eno	r->1	
å ens	t->1	
å er 	e->1	s->1	ä->1	
å er,	 ->1	
å era	 ->1	
å erk	ä->1	
å ers	ä->1	
å ert	 ->1	
å eta	p->1	
å ett	 ->172	
å eur	o->14	
å exa	k->1	
å exe	m->2	
å fak	t->2	
å fal	l->4	
å fam	i->2	
å far	l->1	t->3	
å fas	t->9	
å fel	 ->1	
å fem	 ->1	t->1	
å fen	o->1	
å fin	n->11	s->1	
å fis	k->2	
å fle	r->3	
å fly	g->2	
å fok	u->1	
å fol	k->2	
å for	d->1	t->4	
å fra	m->22	
å fre	d->1	s->1	
å fri	 ->1	v->1	
å frå	g->17	n->13	
å ful	l->2	
å fun	d->1	
å fyr	a->2	
å fäl	t->5	
å fär	r->1	
å få 	h->1	k->1	m->1	
å får	 ->7	
å fåt	t->2	
å föl	j->4	l->1	
å för	 ->42	b->4	d->2	e->47	h->8	k->1	l->4	m->1	n->2	o->1	p->1	s->14	t->1	u->1	
å föt	t->2	
å gar	a->2	
å gat	o->1	
å ge 	e->1	m->1	
å gem	e->16	
å gen	a->1	e->1	o->6	
å geo	g->1	
å ger	 ->1	
å giv	e->1	
å gla	d->1	
å glo	b->1	
å god	a->1	k->1	t->1	
å got	t->1	
å gra	v->3	
å gru	n->82	p->1	
å grä	n->1	
å gäl	l->2	
å gär	n->2	
å gå 	m->1	
å gån	g->5	
å går	 ->3	
å gör	 ->3	,->1	.->1	a->2	
å ha 	e->1	h->1	k->1	r->1	v->1	
å had	e->2	
å han	 ->1	d->4	
å har	 ->11	
å hat	t->1	
å hav	 ->1	e->4	
å hel	a->1	h->1	t->7	
å hem	 ->1	.->1	m->1	
å het	a->1	t->1	
å hin	d->1	
å hjä	l->2	r->4	
å hom	o->1	
å hop	p->1	
å hos	 ->1	
å hot	 ->1	
å hur	 ->19	
å huv	u->1	
å hän	d->1	v->1	
å här	 ->4	.->1	
å häv	t->1	
å hål	l->1	
å hög	 ->1	a->2	
å i A	l->1	
å i S	c->1	
å i T	i->1	
å i b	u->1	
å i c	i->1	
å i d	a->2	e->8	i->1	
å i e	g->1	n->7	t->1	
å i f	e->1	r->1	ö->3	
å i g	å->1	
å i k	a->1	o->2	u->1	
å i l	e->1	j->1	
å i n	o->1	
å i p	r->1	
å i r	a->1	
å i s	i->1	t->2	y->4	
å i v	i->1	ä->1	å->1	
å iak	t->1	
å ick	e->1	
å idé	n->1	
å ige	n->4	
å igå	n->1	
å iho	p->1	
å ill	a->1	e->1	
å imp	o->1	
å in 	f->1	i->1	p->13	
å inf	o->2	r->1	ö->2	
å ing	e->2	i->1	å->1	
å ini	t->1	
å inl	e->1	ä->1	
å inn	a->1	e->5	
å ino	m->1	
å inr	e->1	ä->4	
å ins	e->3	p->2	t->4	
å int	e->27	r->2	
å inv	e->2	o->1	
å irl	ä->1	
å ita	l->1	
å jag	 ->7	
å jak	t->1	
å jor	d->2	
å ju 	p->1	
å jus	t->2	
å jär	n->3	
å kad	m->1	
å kal	l->11	
å kam	p->2	
å kan	 ->23	d->1	s->2	
å kat	a->2	
å kla	r->6	s->1	
å kli	m->1	
å knu	t->1	
å kol	d->1	l->4	
å kom	 ->1	m->40	p->2	
å kon	c->1	j->1	k->8	s->10	t->4	
å kor	r->1	t->9	
å kra	f->1	v->1	
å kri	t->4	
å krä	v->1	
å kun	n->2	s->1	
å kva	l->1	r->2	
å kvi	n->2	
å kän	d->1	
å kär	n->2	
å kör	n->1	s->1	
å lag	a->1	s->2	t->1	
å lan	d->13	
å lig	g->1	
å lik	a->2	n->1	
å lis	t->3	
å lit	e->3	
å lob	b->1	
å lok	a->2	
å los	s->1	
å lov	 ->1	
å lyc	k->1	
å läg	g->2	
å läm	n->1	p->3	
å län	d->2	g->23	
å läs	a->1	
å lät	t->2	
å låg	 ->4	a->1	
å lån	g->18	
å låt	 ->1	
å lör	d->1	
å maj	o->1	
å man	 ->2	d->1	
å mar	k->13	
å mas	s->1	
å med	 ->20	b->2	e->4	l->13	v->2	
å mel	l->3	
å men	 ->1	a->2	
å mer	 ->6	
å mig	,->1	:->1	
å mil	i->1	j->12	
å min	 ->11	a->1	d->1	i->3	n->1	s->2	u->2	
å mis	s->1	
å mit	t->1	
å mod	e->2	
å mon	o->1	
å mot	i->1	s->2	t->1	
å myc	k->43	
å män	g->1	n->1	
å mål	 ->1	.->1	e->1	
å mån	a->3	g->21	
å mås	t->17	
å måt	t->2	
å möj	l->10	
å nat	i->3	t->1	
å ned	e->1	l->1	
å nog	a->1	
å nor	d->1	m->1	r->1	
å not	e->3	
å ny 	k->2	
å nya	 ->4	
å nyc	k->1	
å nys	s->1	
å nyt	t->21	
å näm	n->2	
å när	 ->6	a->2	
å näs	t->4	
å nät	e->1	
å någ	o->24	r->7	
å nåt	t->1	
å nöd	v->4	
å oac	c->2	
å obe	r->1	s->1	
å obl	i->1	
å och	 ->48	
å ock	s->6	u->1	
å oen	s->1	
å off	r->1	
å oft	a->5	
å ogy	n->1	
å oli	k->3	
å olj	e->3	
å om 	1->1	a->4	d->2	e->1	f->1	g->1	h->1	m->1	n->2	ö->1	
å omf	a->1	
å omk	r->1	
å omr	å->15	ö->1	
å omt	a->1	
å ons	d->2	
å ord	e->1	f->2	n->1	
å org	a->1	
å ors	a->1	
å oss	 ->7	
å pap	p->1	
å par	l->4	
å pas	s->2	
å pen	g->2	
å per	m->1	r->1	s->3	
å pes	t->1	
å pla	c->1	n->1	t->9	
å pol	i->2	
å pos	i->2	
å poä	n->1	
å pre	s->1	
å pri	n->3	o->2	s->3	
å pro	b->3	c->1	d->2	g->1	
å pun	k->9	
å på 	8->1	I->1	a->5	d->1	e->2	g->1	j->1	m->1	o->1	s->1	t->1	
å påm	i->3	
å påp	e->2	
å påt	a->1	
å påv	e->1	
å ran	n->1	
å ras	i->1	
å rat	i->1	
å rea	g->1	
å red	a->4	
å ref	o->2	
å reg	e->14	i->1	l->1	
å rek	o->1	
å res	a->1	o->1	p->3	u->7	
å rik	l->1	t->3	
å ris	k->2	
å ryg	g->2	
å räc	k->2	
å räd	s->1	
å räk	n->2	
å rät	t->12	
å råd	e->9	f->1	
å röd	a->1	
å rös	t->2	
å sad	e->1	
å sak	e->5	
å sam	a->2	b->1	m->26	s->2	
å san	t->2	
å sat	s->1	
å se 	d->1	e->1	f->2	h->2	i->1	p->1	r->1	s->1	t->1	v->1	ö->1	
å sed	e->1	
å sek	r->2	t->1	
å sem	e->1	
å sen	a->7	t->1	
å ser	 ->1	b->1	
å ses	 ->1	
å sif	f->1	
å sig	 ->7	.->1	
å sik	t->7	
å sin	 ->7	a->10	
å sis	t->1	
å sit	t->4	u->1	
å sjä	l->3	
å ska	d->1	l->11	n->1	p->3	t->1	
å ske	 ->1	r->2	
å ski	l->1	
å sko	g->2	
å sku	l->10	t->1	
å sky	d->1	
å skä	l->2	
å slu	t->2	
å slå	 ->1	
å smi	d->1	
å små	 ->3	n->4	
å sna	b->15	r->16	
å soc	i->2	
å som	 ->38	
å spe	c->1	l->9	
å spr	å->1	
å spå	r->1	
å sta	b->1	d->3	l->1	n->4	r->1	t->3	
å ste	g->2	
å sto	r->13	
å str	a->1	i->1	u->3	ä->2	ö->1	
å stu	d->1	g->1	
å stä	l->1	r->1	
å stö	d->8	r->1	
å sub	v->2	
å sva	g->1	
å svå	r->4	
å syd	k->1	
å syf	t->1	
å sys	s->2	t->1	
å säg	a->13	e->2	
å säk	e->5	r->2	
å sär	s->2	
å sät	t->17	
å så 	f->1	k->1	l->3	m->2	s->15	t->1	v->2	ä->1	
å såd	a->3	
å såv	ä->2	
å ta 	a->1	d->3	e->1	h->2	i->1	s->2	u->2	
å tac	k->7	
å tal	 ->1	,->1	.->1	a->7	m->3	
å tan	k->1	
å tar	 ->1	
å tas	 ->2	
å tek	n->1	
å tem	a->1	
å ter	r->1	
å tex	t->1	
å tid	e->3	i->3	p->1	
å til	l->57	
å tim	m->3	
å tjä	n->1	
å tog	 ->1	
å top	p->1	
å tor	p->2	s->7	
å tra	n->3	v->1	
å tre	 ->4	d->2	
å tro	r->3	v->1	
å trö	s->3	
å tvi	n->1	
å tvä	r->1	
å två	 ->5	:->1	
å tyc	k->1	
å tyd	l->1	
å tys	k->1	
å tän	k->3	
å und	e->9	v->1	
å ung	a->1	
å uni	o->6	
å upp	 ->3	d->1	e->1	g->2	h->1	k->1	l->1	m->4	n->4	r->2	s->1	
å ut 	a->1	h->1	m->2	ö->2	
å ut,	 ->1	
å uta	n->3	
å utf	l->1	o->1	
å utg	ö->2	
å uto	m->2	
å utr	e->1	
å uts	k->1	u->1	
å utt	r->1	
å utv	e->1	i->2	
å utö	v->1	
å vad	 ->12	
å vak	t->1	
å val	d->2	
å van	l->1	
å var	 ->4	a->14	f->5	g->1	i->3	
å vat	t->1	
å vec	k->1	
å ved	e->4	
å vem	 ->2	
å ver	k->5	
å vet	 ->2	a->6	e->3	
å vi 	a->1	b->1	h->2	k->2	s->3	t->1	ä->1	
å via	 ->1	
å vic	e->1	
å vid	 ->1	a->13	t->1	
å vik	t->18	
å vil	j->9	k->14	l->6	s->1	t->1	
å vis	 ->2	a->2	s->5	u->2	
å vit	t->1	
å vre	d->1	
å väg	 ->10	,->8	.->1	N->1	a->4	e->5	
å väl	 ->2	.->1	k->1	
å vär	d->1	l->2	
å väs	e->1	t->1	
å vår	 ->6	a->13	d->1	t->6	
å ytt	e->3	
å zig	e->2	
å Öst	e->2	
å ägn	a->1	
å än 	e->1	k->1	
å änd	a->1	l->1	r->5	
å änn	u->2	
å änt	l->1	
å är 	a->2	b->3	d->14	e->6	f->3	i->1	j->2	k->2	n->3	o->1	p->2	r->1	s->2	v->2	
å äve	n->3	
å åhö	r->1	
å år 	2->1	e->1	h->1	l->1	s->2	
å år,	 ->1	
å års	 ->1	
å åsi	k->1	
å åt 	d->1	
å åta	g->1	
å åte	r->4	
å åtg	ä->4	
å åtm	i->2	
å öka	t->2	
å ön 	N->1	
å öns	k->1	
å öpp	e->6	
å öve	r->6	
å, al	l->1	
å, at	t->3	
å, bö	r->2	
å, dä	r->1	
å, el	l->1	
å, en	l->1	
å, et	t->1	
å, fr	a->1	u->1	å->1	
å, fö	r->4	
å, ge	n->1	
å, he	r->2	
å, hu	r->1	
å, i 	l->1	s->1	
å, lö	n->1	
å, me	n->7	
å, nu	 ->1	
å, nä	m->2	r->1	
å, ob	e->1	
å, oc	h->8	
å, of	t->1	
å, om	 ->3	
å, ri	k->1	
å, rä	t->1	
å, rö	r->1	
å, so	m->1	
å, st	ö->1	
å, så	 ->2	
å, ti	l->1	
å, vi	l->1	
å, vå	g->1	
å, är	 ->1	
å. De	t->2	
å....	(->1	
å.Att	 ->2	
å.Bet	ä->1	
å.Bis	t->1	
å.Bri	s->1	
å.De 	k->1	
å.Den	 ->2	
å.Det	 ->7	t->3	
å.Doc	k->1	
å.Där	f->1	i->1	
å.En 	g->1	
å.Eur	o->2	
å.FPÖ	 ->1	
å.Fru	 ->1	
å.För	 ->2	
å.Gen	o->1	
å.Gra	t->1	
å.Her	r->2	
å.I s	t->1	
å.Int	e->1	
å.Jag	 ->8	
å.Jus	t->1	
å.Jäm	f->1	
å.Men	 ->1	
å.Ni 	h->1	
å.Nor	m->1	
å.När	 ->2	
å.Och	 ->1	
å.Om 	l->1	
å.Ord	f->1	
å.På 	d->2	
å.Slu	t->1	
å.Soc	i->1	
å.Uni	o->1	
å.Vi 	b->1	m->2	t->1	
å.Är 	d->1	s->1	
å: at	t->1	
å: de	n->2	
å: fö	r->2	
å: Öp	p->1	
å: å 	e->1	
å; de	t->1	
å?. (	E->1	
å?Int	e->1	
å?Jag	 ->1	
å?Ser	i->1	
åbar 	v->2	
åbero	p->1	
åbjud	e->1	
åbörj	a->11	
åd (a	r->1	
åd - 	m->1	
åd an	t->1	
åd at	t->1	
åd be	h->1	
åd fr	å->2	
åd fö	r->1	
åd i 	s->1	
åd nä	r->1	
åd oc	h->2	
åd om	 ->3	
åd so	m->3	
åd, b	o->1	
åd, m	e->1	
åd, o	c->2	
åd.De	t->1	
åd.Ja	g->1	
åd.Ka	n->1	
åd.Lå	t->1	
åd.Me	n->1	
åd?Är	 ->1	
åda a	v->1	
åda b	e->1	o->2	
åda d	e->3	o->3	
åda e	n->1	t->4	
åda f	a->1	ö->6	
åda g	ä->1	
åda h	a->1	
åda i	n->1	
åda l	ä->2	
åda m	e->2	ä->1	
åda n	å->1	
åda o	m->2	r->1	
åda p	a->2	
åda s	i->3	
åda, 	h->1	
ådad 	s->1	
ådade	 ->2	
ådan 	-->1	a->3	b->2	d->3	e->3	f->5	h->5	i->3	j->1	k->4	l->1	m->5	n->2	o->2	p->2	r->3	s->4	u->3	v->2	ä->2	ö->1	
ådan,	 ->2	
ådan.	D->1	S->1	
ådan?	H->1	
ådana	 ->49	
ådand	e->5	
ådant	 ->53	,->1	
ådar 	s->1	
ådar.	D->1	
ådare	 ->1	
ådarn	a->1	
ådd m	e->1	
ådda 	k->1	m->1	r->2	
ådde 	4->1	f->1	i->1	
åddes	 ->1	
åde -	 ->1	
åde D	a->1	
åde S	v->1	w->1	
åde a	n->1	v->4	
åde b	r->1	u->1	
åde d	e->5	j->1	ä->4	
åde e	f->1	l->1	t->1	x->1	
åde f	i->1	r->1	å->1	ö->6	
åde g	o->1	
åde h	a->2	ä->2	
åde i	 ->5	n->4	
åde k	a->2	r->1	u->1	
åde m	a->1	e->9	i->1	ä->2	ö->1	
åde n	a->1	ä->1	
åde o	c->7	
åde p	a->1	o->1	r->1	å->1	
åde r	e->2	
åde s	e->1	k->1	o->5	t->2	å->1	
åde t	i->1	
åde v	a->2	e->1	i->1	
åde ä	r->5	
åde å	s->1	
åde ö	v->1	
åde, 	a->2	d->1	h->2	i->2	m->1	o->4	t->1	ä->1	
åde. 	V->1	
åde.D	e->4	
åde.F	r->1	ö->3	
åde.I	 ->1	d->1	
åde.J	a->3	
åde.M	e->2	i->1	å->1	
åde.O	c->2	
åde.P	l->1	
åde.T	a->1	
åde.V	a->1	
åde: 	h->1	
åde; 	m->1	
åde?D	e->1	
ådefö	r->1	
åden 	-->2	a->1	b->2	d->5	e->1	f->5	g->1	i->10	k->3	m->3	o->8	r->1	s->17	t->1	ä->1	
åden)	 ->1	
åden,	 ->10	
åden.	D->4	F->2	I->1	J->1	K->1	M->3	O->1	P->1	S->2	V->3	Ä->1	
åden:	 ->2	
åden;	 ->1	
åden?	D->2	
ådena	 ->18	,->10	.->7	s->1	
ådens	 ->1	
åder 	b->2	d->2	e->5	f->3	i->6	m->3	s->2	t->3	
åder)	 ->2	F->2	J->1	K->1	T->1	
ådera	d->1	r->2	
ådet 	(->7	-->2	A->1	B->1	S->1	a->17	b->5	d->2	e->4	f->22	g->7	h->19	i->16	j->1	k->15	l->3	m->10	n->2	o->33	r->3	s->14	t->5	u->8	v->7	ä->7	
ådet)	N->1	
ådet,	 ->47	
ådet.	 ->4	(->1	.->1	D->6	E->4	F->1	H->1	I->2	J->9	L->1	M->4	N->3	O->1	P->3	S->1	T->1	U->1	V->5	Ä->1	Å->2	
ådet:	 ->1	
ådet?	.->2	H->1	I->1	
ådets	 ->98	,->1	
ådfrå	g->6	
ådgiv	a->23	n->3	
ådgör	 ->1	
ådlig	 ->4	a->1	t->2	
ådnin	g->1	
ådrag	 ->1	
ådsbe	s->1	
ådska	 ->1	n->18	r->1	
ådsla	g->3	
ådsme	d->1	
ådsmi	n->1	
ådsmö	t->1	
ådsor	d->20	
ådsrä	t->1	
ådsto	p->1	
åelig	 ->1	a->1	t->4	
åelse	 ->7	n->1	
ående	 ->103	,->1	.->5	:->21	n->3	t->3	
åer g	e->1	
åer i	 ->2	n->1	
åer o	c->1	
åer s	o->1	
åer, 	e->1	i->1	n->1	
åer.D	e->2	
åer.K	o->1	
åer.M	i->1	
åer: 	d->1	
åerna	.->1	
ået.D	e->1	
åfres	t->1	
åfölj	a->1	d->3	
åföre	t->6	
åg Ir	l->1	
åg ar	b->1	
åg at	t->15	
åg av	 ->2	
åg de	 ->1	m->1	t->3	
åg dä	r->1	
åg el	l->1	
åg et	t->1	
åg hö	j->1	
åg in	k->1	t->1	
åg ni	v->2	
åg nå	g->1	
åg om	 ->1	
åg re	g->1	
åg si	g->1	t->1	
åg so	m->1	
åg ti	l->1	
åg ut	 ->2	
åg Ös	t->1	
åg är	 ->1	
åg, v	i->1	
åg.Eu	r->1	
åga -	 ->1	
åga a	n->1	t->14	v->3	
åga b	e->1	i->1	o->1	
åga e	f->1	r->1	
åga f	o->1	ö->6	
åga g	e->2	r->1	ä->3	
åga h	a->5	u->2	ö->2	
åga i	 ->7	n->2	
åga j	a->1	
åga k	a->2	o->6	
åga m	e->5	i->1	å->1	
åga n	i->1	r->24	ä->2	
åga o	b->1	c->8	m->71	s->3	
åga p	a->1	å->2	
åga r	e->1	å->2	ö->1	
åga s	i->4	k->4	o->37	p->1	ä->1	
åga t	a->1	e->1	i->2	o->1	
åga v	a->1	e->1	i->4	
åga ä	r->9	
åga ö	p->1	
åga!F	r->1	
åga, 	a->2	d->3	e->2	f->3	h->1	k->2	n->1	o->4	s->5	v->3	
åga. 	M->1	
åga.-	 ->1	
åga.A	n->1	
åga.D	e->7	ä->1	
åga.E	n->1	t->1	
åga.F	r->1	ö->1	
åga.H	e->3	
åga.I	 ->2	
åga.J	a->8	
åga.M	e->2	
åga.N	i->1	
åga.O	c->1	m->1	
åga.S	o->1	
åga.T	i->1	
åga.U	t->1	
åga.V	i->5	
åga.Ä	v->1	
åga: 	N->1	h->2	o->1	v->3	
åga?.	 ->1	
ågade	 ->6	,->1	s->1	
ågan 	-->2	1->1	a->4	c->1	d->3	f->7	g->5	h->2	i->11	j->1	k->2	m->1	n->3	o->98	p->1	r->1	s->6	t->1	u->2	v->3	y->1	ä->16	å->1	
ågan,	 ->14	
ågan.	D->1	E->1	F->3	H->2	I->1	J->4	K->1	S->2	U->1	
ågan:	 ->5	
ågan;	 ->1	
ågan?	J->1	
ågand	e->1	
ågar 	d->1	h->1	i->1	j->4	k->1	m->4	n->1	o->6	s->4	ä->1	
ågar.	V->1	
ågasa	t->1	
ågasä	t->19	
ågat 	e->2	m->1	
ågat,	 ->1	
ågata	 ->1	
ågats	 ->1	.->1	
ågava	r->1	
ågeko	m->1	
ågell	i->1	
ågels	k->1	
ågelv	ä->1	
ågen 	a->1	
ågeri	.->1	
ågerp	o->1	
ågest	u->7	ä->3	
åget 	i->1	
ågete	c->2	
ågick	 ->3	
ågkra	s->2	
åglar	 ->4	,->2	
åglän	g->1	
ågnin	g->8	
ågoly	c->1	
ågon 	a->13	b->5	c->1	d->3	e->5	f->4	g->7	i->4	j->1	k->8	l->3	m->5	n->5	o->3	p->4	r->8	s->18	t->7	u->3	v->2	å->1	
ågon,	 ->2	
ågon.	I->1	
ågons	i->11	t->4	
ågont	i->39	
ågor 	-->1	a->10	b->6	d->3	e->4	f->4	g->4	h->6	i->11	k->1	l->1	m->3	o->41	p->3	s->54	t->10	u->2	v->8	ä->5	
ågor)	 ->1	
ågor,	 ->37	
ågor.	 ->1	.->1	D->10	F->4	H->1	J->2	K->2	M->1	N->2	S->1	V->3	
ågor:	 ->4	
ågor;	 ->1	
ågor?	,->1	
ågorl	u->1	
ågorn	a->28	
ågot 	E->1	K->1	a->22	b->3	d->3	e->3	f->15	h->1	i->4	j->4	k->2	l->6	m->10	o->10	p->5	r->2	s->75	t->4	u->2	v->10	å->1	
ågot,	 ->2	
ågot.	A->1	D->2	J->1	S->1	Ä->1	
ågot?	N->1	
ågra 	-->1	a->24	b->5	d->4	e->5	f->10	g->6	h->1	i->6	k->11	m->9	n->3	o->5	p->9	r->2	s->19	t->7	u->3	v->7	ä->3	å->8	ö->1	
ågrup	p->3	
ågräl	,->1	
ågs i	 ->1	
ågs m	e->1	
ågs.J	a->1	
ågs.L	å->1	
ågt s	t->1	
ågt v	ä->1	
ågver	k->1	
ågå i	 ->1	
ågåen	d->6	
ågår 	d->1	e->1	f->1	i->2	p->1	s->1	
ågår.	 ->1	I->1	J->1	
ågått	 ->1	
åhund	r->1	
åhänd	a->6	
åhär.	V->1	
åhöra	r->1	
åja, 	d->1	
åk fö	r->1	
åk på	 ->3	
åk ti	l->1	
åk. D	e->1	
åka e	n->1	
åkar 	f->1	s->2	v->2	
åkare	 ->2	.->1	
åkarn	a->1	
åket 	a->1	m->1	
åket.	I->1	N->1	
åkigt	 ->3	
åklag	a->37	
åklig	 ->1	a->2	
åkomr	å->2	
åkrat	e->2	i->28	
åktag	a->1	
åkte 	t->1	
ål (B	r->1	
ål 1 	o->2	
ål 1,	 ->2	
ål 1-	o->4	r->5	s->2	
ål 1.	J->1	
ål 2 	-->1	b->1	e->1	o->1	s->1	
ål 2,	 ->1	
ål 2-	o->2	s->1	
ål 2.	M->1	
ål 5b	 ->1	.->1	
ål at	t->3	
ål av	t->1	
ål be	t->2	
ål en	l->1	
ål fi	n->1	
ål fö	r->19	
ål gå	 ->1	
ål he	l->1	
ål hi	n->1	
ål i 	1->1	k->1	s->5	
ål ja	g->1	
ål li	g->1	
ål nå	g->1	
ål oc	h->5	
ål om	 ->3	
ål på	 ->2	
ål rö	r->1	
ål sk	a->1	
ål so	m->13	
ål sä	t->1	
ål ti	l->1	
ål up	p->2	
ål är	 ->4	
ål, R	e->1	
ål, f	r->1	ö->1	
ål, g	e->1	
ål, h	a->1	
ål, m	e->2	
ål, n	ä->1	
ål, o	c->1	
ål, p	r->1	
ål, s	o->4	å->2	
ål, u	t->1	
ål-2-	o->1	
ål.Bä	s->1	
ål.De	n->2	
ål.Dä	r->1	
ål.Et	t->1	
ål.Fr	u->1	
ål.He	r->2	
ål.I 	e->1	f->1	
ål.Ja	g->1	
ål.Ku	l->1	
ål.Ma	r->1	
ål.Me	n->1	
ål.Nä	r->2	
ål.Äv	e->1	
ål: V	i->1	
ål: a	t->1	
åla b	i->1	
åla f	o->1	
åla, 	a->1	
ålagd	 ->1	
ålago	r->1	
ålagt	s->2	
ålamo	d->2	
ålare	 ->2	
ålarf	ä->1	
åld i	 ->1	
åld o	c->1	
ålder	 ->5	.->3	d->2	n->2	
åldet	 ->1	,->1	
åldra	d->3	
åldsa	m->3	
åldsh	a->2	
åldsu	t->1	
åldta	 ->1	g->1	
ålede	s->44	
ålen 	E->1	a->1	b->1	e->1	f->3	h->1	i->2	n->1	s->2	ä->1	å->1	
ålen.	 ->1	D->1	
ålens	 ->1	
ålet 	a->3	e->1	f->1	i->1	k->2	m->11	o->1	ä->3	
ålet,	 ->2	
ålet.	A->1	F->1	H->1	J->2	
ålför	e->5	
ålgem	e->1	
ålig 	f->2	g->1	l->1	s->1	
åliga	 ->8	
åligg	e->5	
åligh	e->1	
åligt	 ->6	,->1	.->1	
ålind	u->25	
ålinr	i->4	
ålitl	i->1	
ålkas	t->1	
åll a	v->1	
åll f	ö->2	
åll h	a->1	
åll i	 ->3	
åll k	a->1	u->1	
åll o	c->3	
åll r	å->1	
åll s	o->3	ä->1	
åll t	i->1	
åll v	a->1	
åll, 	m->1	o->2	t->1	ä->1	
åll.D	e->2	
åll.F	ö->1	
åll.I	 ->1	
åll.J	a->2	
åll.V	i->1	
åll: 	"->1	
åll?.	 ->1	
ålla 	a->1	b->1	d->11	e->12	f->9	g->1	h->3	i->2	k->3	l->2	m->8	n->2	o->2	p->2	r->2	s->8	t->11	u->1	v->3	ä->1	
ålla,	 ->1	
ållan	d->84	
ållar	 ->1	
ållas	 ->9	,->1	.->1	
ållba	r->25	
ållen	 ->1	
åller	 ->92	,->2	
ållet	 ->19	,->5	.->3	
ållit	 ->16	,->1	s->6	
ållna	,->1	
ållni	n->66	
ålls 	a->1	e->1	f->1	i->1	
ålls,	 ->1	
ålls.	D->1	
ållsa	m->2	
ållsl	i->1	ö->1	
ållsm	ä->2	
ållsr	i->2	
ållst	i->7	
ållsv	i->1	
ålmed	v->1	
ålnin	g->3	
ålsdo	m->1	
ålsek	t->5	
ålsen	l->2	
ålsky	d->1	
ålssi	d->1	
ålsti	l->1	
ålsät	t->17	
ålund	a->4	
ålver	k->5	
ålägg	a->4	e->2	
åmind	e->1	
åminn	a->21	e->8	
ån (H	-->21	
ån - 	d->1	Ö->1	
ån 10	5->1	
ån 15	 ->1	
ån 19	6->1	9->4	
ån 28	 ->1	
ån 3,	8->1	
ån 5 	0->2	
ån 50	-->1	
ån 89	 ->1	
ån 95	 ->1	
ån Af	r->1	
ån Al	b->1	t->1	
ån Am	s->4	
ån At	a->2	
ån Au	t->1	
ån BS	E->1	
ån Ba	s->1	
ån Bo	n->1	
ån Br	e->1	y->1	
ån CE	N->2	
ån Ca	n->1	
ån Da	l->1	
ån De	 ->1	
ån EG	-->2	
ån EU	?->1	
ån Er	i->2	
ån Eu	r->24	
ån FM	I->1	
ån Fl	o->3	
ån Fr	a->1	
ån Fö	r->1	
ån GU	E->1	
ån Ga	l->1	
ån Go	l->1	
ån Gö	t->1	
ån He	l->2	
ån IR	A->1	
ån In	d->1	t->2	
ån Is	r->1	
ån Ja	p->1	
ån Ko	r->1	
ån Ky	o->2	
ån Kö	l->1	p->1	
ån La	n->1	
ån Li	s->1	
ån Lo	i->1	
ån Ma	r->1	
ån Na	t->3	
ån OS	S->1	
ån PP	E->2	
ån PS	E->1	
ån Pa	r->1	
ån Po	l->1	r->2	
ån Ro	t->1	
ån Sa	m->3	
ån Sh	a->1	
ån Sy	d->1	r->1	
ån Ta	m->4	
ån Te	r->1	
ån Ty	s->1	
ån UN	I->1	
ån US	A->1	
ån Ve	n->1	
ån Wi	e->1	
ån Wu	r->1	
ån al	l->4	
ån an	d->3	
ån at	t->26	
ån av	 ->2	f->1	
ån be	f->1	
ån bi	d->1	l->3	
ån bo	n->2	
ån bu	d->2	
ån bö	r->5	
ån da	g->3	
ån de	 ->25	c->2	m->2	n->36	p->1	r->2	t->21	
ån di	k->1	r->2	s->1	
ån do	m->1	
ån dr	a->1	
ån dä	r->1	
ån en	 ->16	e->1	k->1	s->1	
ån er	 ->1	,->1	a->1	
ån et	t->17	
ån eu	r->1	
ån ex	t->3	
ån fa	r->2	
ån fl	a->1	e->1	
ån fr	a->1	å->1	
ån fö	n->1	r->38	
ån ge	m->3	r->1	
ån ha	m->1	n->1	r->1	v->1	
ån he	l->1	
ån hö	g->2	
ån i 	d->1	f->1	m->1	
ån ju	l->1	n->1	s->2	
ån ka	m->1	n->1	r->1	
ån ko	l->1	m->31	n->2	
ån la	n->1	
ån le	d->3	
ån li	k->1	
ån lä	n->4	
ån ma	j->1	r->3	
ån me	d->7	
ån mi	l->5	n->3	
ån mo	r->1	t->1	
ån må	l->2	
ån na	t->1	
ån ny	h->1	l->1	
ån nå	g->3	
ån ob	e->1	
ån oc	h->11	
ån of	f->1	
ån ol	i->4	
ån om	 ->1	
ån op	p->1	
ån or	d->2	
ån os	s->2	
ån pa	r->13	
ån pe	d->1	
ån pr	i->1	o->3	
ån på	 ->3	
ån ra	p->1	
ån re	d->1	g->2	
ån rå	d->13	
ån sa	m->3	
ån se	r->1	
ån si	g->1	n->5	t->2	
ån sk	a->2	r->1	
ån so	c->2	
ån st	a->1	r->3	
ån sy	s->1	
ån sä	g->1	k->2	
ån så	d->1	
ån sö	d->1	
ån t.	e->1	
ån ti	d->1	l->4	
ån to	p->2	
ån tr	a->1	e->15	
ån tu	n->1	
ån un	i->2	
ån ut	l->1	s->17	t->2	
ån va	r->2	
ån ve	r->1	
ån vi	c->1	l->1	s->3	
ån vä	n->1	
ån vå	g->1	l->1	r->8	
ån Ös	t->1	
ån är	 ->1	
ån år	 ->1	
ån öv	r->4	
ån, d	u->1	
ån, f	r->1	
ån, n	ä->1	
ån, o	c->1	
ån.De	 ->1	t->2	
ån.Dä	r->1	
ån.Hä	r->1	
ån.Än	d->1	
åna m	i->1	
åna o	m->3	
ånad 	-->1	d->1	k->1	m->1	o->2	s->1	u->1	ö->1	
ånad,	 ->2	
ånad.	D->1	J->1	P->1	
ånade	 ->1	n->3	r->55	
ånads	l->1	
ånand	e->2	
ånar 	d->1	
ånare	 ->6	
ånarn	a->5	
ånas 	ö->1	
ånbok	e->1	
ånd a	n->1	t->4	
ånd d	e->2	
ånd e	f->1	n->6	
ånd f	r->6	ö->1	
ånd h	a->2	
ånd i	 ->5	
ånd k	a->1	o->1	
ånd m	e->3	
ånd n	ä->1	
ånd o	c->6	m->1	
ånd p	å->1	
ånd s	o->4	t->1	
ånd t	i->4	
ånd v	i->1	
ånd ä	r->1	
ånd å	t->1	
ånd, 	E->1	d->1	k->1	m->1	o->2	r->1	s->1	
ånd. 	V->1	
ånd.A	t->1	
ånd.D	e->3	
ånd.F	r->1	
ånd.H	e->1	
ånd.J	a->1	
ånd.V	a->1	i->1	
ånd?.	 ->1	
ånd?J	a->1	
åndag	 ->1	s->2	
åndar	e->4	n->1	
ånde.	U->1	
åndel	s->1	
ånden	 ->6	,->2	.->1	?->1	
åndet	 ->16	,->2	s->1	
åndig	a->1	
åndpu	n->97	
ånds 	o->1	
åndsd	e->12	
åndsp	o->2	
åndsr	ö->1	
åndss	y->1	
åndst	a->2	
åner 	o->1	
åner.	Ä->1	
ång -	 ->1	
ång a	j->1	l->2	n->1	t->1	v->4	
ång b	e->4	ö->1	
ång d	e->4	i->1	ä->1	
ång e	l->1	n->3	t->2	
ång f	r->1	å->1	ö->10	
ång h	a->5	e->1	
ång i	 ->5	n->1	r->1	
ång k	a->1	o->3	
ång l	i->1	
ång m	e->2	
ång n	i->1	
ång o	c->6	
ång p	e->2	r->2	å->2	
ång r	a->1	e->1	i->1	ä->1	
ång s	a->1	e->1	i->9	k->3	o->4	t->1	ä->1	
ång t	a->2	i->30	r->1	y->1	
ång u	n->2	p->1	r->1	t->2	
ång v	a->1	e->1	i->1	o->1	ä->2	
ång ä	r->4	
ång ö	k->1	
ång".	N->1	
ång, 	a->1	e->1	f->1	i->1	l->1	o->2	r->1	t->1	u->1	v->1	
ång.D	e->4	ä->1	
ång.F	r->1	
ång.H	ö->1	
ång.J	a->1	
ång.N	u->1	ä->1	
ång.O	c->1	
ång.T	r->1	
ång.V	i->2	
ånga 	-->1	a->36	b->8	c->1	d->8	e->3	f->12	g->6	h->2	i->4	k->4	l->3	m->11	n->3	o->9	p->2	r->1	s->13	t->8	u->2	v->4	ä->6	å->9	ö->1	
ånga,	 ->2	
ånga.	J->2	
ångar	 ->7	,->1	.->3	e->3	n->2	
ångas	 ->1	
ångdr	a->1	
ångel	 ->1	
ången	 ->38	,->3	.->4	
ånger	 ->19	,->4	.->3	
ånget	 ->1	
ångfa	l->15	
ångfr	i->1	
ångfu	n->1	
ångfä	r->2	
ångkö	r->1	
ångli	g->1	
ångmå	l->1	
ångna	 ->2	
ångra	n->2	
ångre	m->1	
ångs 	s->3	
ångsa	m->6	r->2	
ångsb	e->3	
ångsf	i->1	
ångsi	d->3	k->7	
ångsp	e->3	r->1	u->11	
ångsr	i->15	
ångss	t->1	y->2	ä->6	
ångst	 ->3	e->2	m->2	r->1	
ångsä	t->1	
ångt 	b->3	d->5	f->2	h->1	i->7	k->2	m->4	n->2	s->4	u->2	v->1	ö->1	
ångt.	D->1	M->1	V->1	
ångtg	å->11	
ångti	d->4	
ångva	r->6	
ångår	 ->1	
åning	 ->1	,->1	e->1	o->4	
ånkom	l->3	
ånspa	k->1	
åntar	 ->1	
åntas	 ->1	
åntog	 ->1	
ånvar	a->4	o->4	
ånvän	d->1	
ånyo 	s->1	
åolja	 ->1	
åpeka	 ->14	,->1	d->7	n->9	r->6	s->3	t->10	
åpsla	g->1	
år - 	o->1	
år 19	7->1	8->1	9->17	
år 20	0->31	1->2	
år Ba	r->1	
år Ma	r->1	
år OL	A->1	
år ad	m->1	
år ak	t->1	
år al	d->1	l->4	
år an	s->2	t->1	
år ar	b->1	
år at	t->32	
år av	 ->14	.->1	
år ba	l->1	
år be	d->3	g->1	h->1	s->3	t->3	
år bi	l->1	
år bo	r->2	
år br	a->1	o->1	
år bu	d->1	
år de	 ->4	b->2	l->8	m->2	n->8	s->3	t->22	
år di	a->1	r->1	s->2	t->1	
år dj	u->1	
år do	c->1	
år dr	a->1	
år du	g->1	
år dä	r->5	
år då	 ->2	
år ef	t->4	
år eg	e->2	
år el	l->3	
år em	e->1	
år en	 ->23	e->1	h->1	
år er	 ->2	,->1	.->1	f->1	
år et	t->9	
år fa	k->1	m->1	r->1	s->1	
år fe	l->1	
år fi	n->2	
år fo	r->3	
år fr	a->8	e->2	ä->1	å->11	
år få	 ->1	
år fö	r->26	
år ge	m->4	n->4	
år gi	v->1	
år gl	ö->1	
år gr	u->16	
år gö	r->2	
år ha	n->1	r->4	
år he	d->1	l->7	
år hä	n->1	r->2	
år hå	l->1	
år hö	g->1	
år i 	E->4	O->1	a->3	d->8	e->4	f->1	h->2	i->1	k->2	m->4	o->2	p->1	r->5	u->1	v->2	Ö->1	
år ib	l->1	
år id	é->1	
år if	r->2	
år ig	e->3	
år in	f->14	g->3	i->1	l->1	n->1	o->3	s->5	t->44	
år ja	g->13	
år ju	 ->1	
år ka	m->1	n->1	r->1	
år kl	a->9	
år ko	l->2	m->9	n->3	
år kr	ä->1	
år ku	l->1	
år kv	ä->1	
år la	g->2	
år le	d->1	v->1	
år li	g->1	k->1	t->2	
år lo	k->1	t->1	
år ly	s->1	
år lä	n->1	
år lå	n->1	t->1	
år ma	n->2	
år me	d->4	l->1	n->3	r->2	s->1	
år mi	g->5	l->4	n->1	
år mo	g->1	r->6	t->1	
år my	c->4	
år må	l->1	n->1	
år mö	j->2	
år na	t->1	
år ni	 ->1	
år no	r->1	
år nu	 ->2	
år ny	a->1	
år nä	r->1	
år nå	g->2	
år nö	d->1	j->1	
år oc	h->8	k->9	
år of	t->2	
år om	 ->2	p->1	
år or	d->2	o->2	
år os	s->1	
år pa	r->1	
år pe	r->1	
år pl	a->1	i->2	
år po	l->3	s->1	
år pr	i->1	o->2	
år på	 ->19	
år re	d->1	g->1	k->2	s->4	
år ro	l->3	
år rä	t->2	
år rö	s->2	
år sa	k->1	m->2	
år se	 ->1	d->14	g->2	n->1	
år si	d->1	n->3	t->1	
år sj	u->1	ä->1	
år sk	a->1	r->3	y->2	
år sl	u->1	
år sn	a->2	ä->1	
år so	l->3	m->10	
år sp	e->1	
år st	i->1	r->3	y->1	å->5	ö->4	
år sv	a->1	
år sä	r->1	
år så	 ->1	v->1	
år ta	 ->4	l->1	s->1	
år ti	d->1	l->31	
år tr	o->2	
år tv	e->1	
år un	d->3	i->4	
år up	p->7	
år ut	 ->9	a->1	f->1	ö->4	
år va	d->2	g->1	r->2	
år ve	r->1	t->1	
år vi	 ->28	,->1	l->1	s->3	t->1	
år vä	g->2	l->1	n->1	
år yt	t->1	
år äg	n->1	
år än	 ->1	n->1	
år är	 ->3	
år äv	e->2	
år å 	e->1	
år ås	i->3	
år åt	 ->2	e->1	g->1	s->1	
år ön	s->2	
år öp	p->1	
år öv	e->2	
år".J	a->1	
år)? 	H->1	
år, E	u->1	
år, a	l->1	
år, d	e->2	
år, e	l->1	n->1	
år, f	i->1	
år, i	n->1	
år, k	a->2	o->1	
år, m	e->3	å->1	
år, n	ä->2	
år, o	a->1	c->5	
år, p	r->1	
år, s	o->1	å->1	
år, t	r->1	
år, u	n->1	t->2	
år, v	i->1	
år, ä	r->1	
år. E	n->1	
år. J	a->1	
år.De	 ->5	s->1	t->6	
år.En	b->1	
år.Fö	r->2	
år.He	r->2	
år.Hu	r->1	
år.Hä	n->1	
år.I 	g->1	v->1	
år.Ja	g->4	
år.Kä	r->1	
år.La	n->1	
år.Ly	c->1	
år.Ma	r->1	
år.Om	 ->1	
år.Re	v->1	
år.Sa	m->1	
år.Ty	 ->1	
år.Ve	m->1	
år.Vi	 ->4	
år.Vå	r->1	
år.Än	d->1	
år?Nä	s->1	
år?So	m->1	
åra a	f->1	m->1	n->4	r->2	t->4	
åra b	a->2	e->2	
åra d	a->1	e->3	i->1	
åra e	g->4	k->1	n->3	r->2	
åra f	a->5	r->6	ö->8	
åra g	r->7	
åra h	a->1	e->1	u->1	
åra i	n->5	
åra k	a->3	o->4	r->4	u->2	
åra l	a->3	i->3	o->1	ä->5	ö->1	
åra m	e->15	i->1	o->1	å->2	
åra n	a->1	y->1	
åra o	l->1	m->1	
åra p	a->1	l->1	o->4	r->3	
åra r	e->12	i->2	u->1	ä->1	
åra s	a->2	i->1	k->1	l->1	t->8	y->1	
åra t	i->1	j->1	r->1	u->1	v->2	
åra u	p->1	
åra v	ä->4	
åra ä	n->5	
åra å	t->6	
åra ö	g->1	r->1	s->1	v->1	
åra, 	i->1	
årand	e->1	
årar 	e->1	
årare	 ->3	.->1	
åras,	 ->1	
årata	l->1	
årbar	a->1	h->1	t->1	
årbed	ö->1	
årbeg	r->1	
ård g	r->1	
ård k	a->1	
ård o	c->2	
ård p	r->1	
ård t	i->1	
ård),	 ->1	
ård, 	o->1	s->1	
årda 	a->1	k->1	n->1	r->2	v->2	
årdag	e->2	
årdar	 ->1	,->1	e->3	
årdas	t->2	
ården	 ->1	
årdna	c->2	
årds-	 ->1	
årdsl	ö->2	
årdsm	y->1	
åren 	2->1	d->1	f->1	g->1	h->9	m->2	o->3	s->5	t->1	u->2	ä->1	
åren,	 ->5	
åren.	D->1	I->1	J->1	K->1	M->1	Ö->1	
årens	 ->2	
året 	-->2	1->10	a->2	f->2	g->2	i->2	k->2	o->1	r->1	s->2	t->1	u->1	ä->1	ö->1	
året,	 ->8	
året.	 ->1	D->1	J->1	
årets	 ->4	
århun	d->7	
åriga	 ->6	.->1	
årigh	e->31	
årigt	 ->7	
åring	a->1	
årkly	v->1	
årköt	t->1	
årlig	a->6	e->2	
årlös	t->2	
årnin	g->2	
års E	G->1	
års b	u->3	
års e	r->1	
års p	r->1	
års s	k->1	
års t	i->3	
års ö	v->1	
årsaf	t->1	
årsbe	l->1	r->1	
årspe	r->1	
årspr	o->1	
årsra	p->2	
årssk	i->2	
årsti	d->1	
årt E	u->2	
årt a	g->1	n->4	r->8	t->19	v->4	
årt b	e->1	o->1	u->1	
årt d	e->4	r->2	
årt e	g->3	k->3	n->1	u->3	
årt f	ö->14	
årt g	e->1	r->2	
årt h	e->1	
årt i	n->2	
årt k	o->1	r->1	u->2	
årt l	a->3	o->1	ö->1	
årt m	e->1	å->4	ö->1	
årt n	u->1	y->1	
årt o	r->3	
årt p	a->8	o->1	r->4	
årt r	e->2	ä->1	
årt s	a->4	p->1	t->6	v->3	y->1	
årt t	a->2	
årt u	p->1	t->11	
årt v	a->1	e->1	ä->1	
årt y	t->1	
årt, 	a->1	b->1	c->1	
årt.M	e->1	
årtal	 ->1	
årtio	n->1	
årtus	e->3	
åröve	r->1	
ås al	l->1	
ås at	t->2	
ås av	 ->1	
ås bl	.->1	i->1	
ås bä	s->1	
ås de	t->2	
ås dä	r->1	
ås en	 ->2	
ås fa	l->1	
ås fö	r->3	
ås ge	n->2	
ås gö	r->1	
ås i 	L->1	d->4	f->1	r->2	s->1	v->3	ä->1	
ås ig	e->1	
ås in	o->1	
ås ko	m->1	
ås mo	t->1	
ås oc	h->1	
ås på	 ->1	
ås sk	u->1	
ås ti	l->2	
ås up	p->1	
ås va	r->1	
ås, i	n->1	
ås.De	t->1	
ås.Fö	r->1	
ås.La	n->1	
ås: a	t->1	
åsamk	a->3	
åsatt	,->1	
åser 	e->1	f->1	i->1	
åsikt	 ->23	,->3	.->2	e->22	
åskal	i->1	
åskyn	d->7	
åskåd	a->1	n->1	
åsom 	"->1	3->1	A->1	C->1	D->1	P->1	T->1	W->1	a->4	b->1	d->3	e->2	f->6	j->1	k->3	n->1	r->1	v->2	ä->1	ö->1	
åss m	e->1	
åst s	i->1	
åsta 	f->1	t->1	
åstad	 ->1	k->24	
åste 	-->2	E->6	F->1	I->1	a->32	b->45	c->1	d->51	e->12	f->46	g->39	h->14	i->32	j->10	k->27	l->9	m->30	n->16	o->28	p->9	r->17	s->69	t->36	u->29	v->106	ä->11	å->6	ö->8	
åste,	 ->3	
åstri	d->1	
åstå 	a->3	o->1	
åstå,	 ->2	
åståe	n->8	
åstår	 ->4	
åstås	 ->2	
åståt	t->1	
åsyft	a->5	
åt Eu	r->1	
åt Fö	r->1	
åt an	v->1	
åt at	t->7	
åt be	s->1	
åt de	 ->6	m->3	n->9	s->1	t->8	
åt eg	n->1	
åt en	 ->3	
åt er	 ->2	
åt et	t->2	
åt fo	r->1	
åt fr	å->1	
åt ge	n->1	
åt hu	r->1	
åt i 	s->4	t->3	v->1	
åt im	m->1	
åt in	f->1	t->1	
åt jä	m->1	
åt ko	m->3	n->1	
åt kv	a->1	
åt li	v->1	
åt ma	r->1	
åt me	d->2	
åt mi	g->55	
åt mo	t->1	
åt nu	.->1	
åt ny	b->1	
åt oc	h->2	
åt os	s->26	
åt pa	r->1	
åt på	 ->1	
åt re	g->1	
åt rä	t->3	
åt sa	m->1	
åt si	d->2	n->1	t->1	
åt sy	f->1	
åt ti	l->1	
åt tv	å->1	
åt tä	n->1	
åt un	d->1	
åt ve	t->1	
åt vå	r->1	
åt Ös	t->1	
åt äm	n->1	
åt är	 ->2	
åt åt	e->1	
åt", 	d->1	
åt, i	 ->1	
åt, k	o->1	
åt, m	e->2	
åt, u	t->1	
åt.Da	g->1	
åt.De	t->1	
åt.Dä	r->1	
åt.Fr	a->1	
åt.He	r->1	
åt.Ja	g->1	
åt.Ko	m->1	
åt.Nä	r->1	
åt.Va	d->1	
åta E	u->1	
åta J	ö->1	
åta a	n->1	t->1	
åta b	l->3	
åta d	e->9	i->1	
åta e	n->1	t->1	
åta f	o->1	ö->1	
åta h	e->1	
åta j	u->1	
åta k	o->1	
åta l	ä->1	
åta m	e->3	i->1	
åta n	u->1	
åta o	s->2	
åta p	a->2	
åta r	e->1	i->1	
åta s	i->6	k->1	
åta t	u->1	
åtaga	n->28	
åtagi	t->2	
åtagl	i->4	
åtal 	i->3	m->1	o->1	s->1	
åtal.	I->1	
åtala	 ->2	?->1	d->1	s->2	t->4	
åtals	f->1	p->6	
åtand	e->3	
åtank	e->1	
åtar 	a->1	g->1	h->1	s->4	
åtar,	 ->2	
åtarn	a->1	
åtas 	a->2	j->1	o->1	p->1	t->1	
åte s	o->1	
åten 	f->1	r->1	t->2	
åtenh	e->2	
åtens	 ->1	
åter 	E->1	K->1	a->5	b->2	d->3	e->1	f->2	g->3	h->1	i->5	j->1	m->1	n->1	o->5	r->1	s->3	t->3	v->1	ä->1	
åter,	 ->1	
åter.	Å->1	
återa	n->18	
återb	e->1	
återe	r->1	
återf	i->3	u->2	ö->8	
återg	a->2	e->4	å->1	
återh	ä->2	å->2	
återi	g->19	n->6	
återk	o->7	r->1	
återl	ä->2	
återn	a->11	
åters	a->1	k->2	p->3	t->27	
återt	a->9	
återu	p->32	
återv	e->1	i->65	u->2	ä->3	
åtet 	a->1	
åtföl	j->12	
åtgär	d->240	
åtgån	g->1	
åtill	v->1	
åtit 	a->1	f->1	
åtits	 ->1	
åtlig	.->1	a->1	t->3	
åtmin	s->27	
åtna 	b->1	f->1	s->1	t->2	
åtna.	S->1	
åtnju	t->1	
åtryc	k->3	
åts e	n->1	
åts f	r->1	
åts m	e->1	
åts å	t->1	
åtsas	 ->2	
åtski	l->3	
åtstr	a->2	ä->1	
ått -	 ->1	
ått 8	 ->1	
ått 9	8->1	
ått E	U->1	
ått K	y->1	
ått a	n->1	r->1	t->3	v->2	
ått b	e->3	
ått d	e->4	å->1	
ått e	n->13	r->2	t->7	
ått f	e->1	o->1	r->4	
ått g	o->1	
ått h	u->1	ö->4	
ått i	 ->4	g->3	n->5	
ått j	u->1	
ått k	l->1	r->1	u->1	
ått l	u->1	
ått m	e->5	i->2	å->2	ö->1	
ått n	y->1	å->6	
ått o	c->3	t->1	
ått p	r->1	å->1	
ått s	a->1	e->2	t->2	
ått t	a->4	i->7	
ått u	p->3	t->1	
ått v	e->4	i->2	ä->1	å->1	
ått y	t->3	
ått ä	r->1	
ått å	t->1	
ått, 	t->1	ä->1	
ått.D	e->2	
ått.F	ö->1	
ått.I	 ->2	
ått.P	a->2	
åtta 	m->1	p->1	r->1	ä->1	
åtta,	 ->1	
åttfu	l->1	
åtto 	a->1	f->1	
åtton	d->1	
åttor	 ->1	
åtts 	a->3	h->1	i->1	m->1	v->1	
åtts.	D->1	R->1	
åtvin	g->4	
åvar 	i->1	
åvara	n->1	
åverk	a->37	
åvida	 ->3	
åvila	r->1	
åvisa	t->2	
åvisb	a->1	
åvor 	t->1	
åvor.	L->1	
åväl 	S->1	a->3	b->1	d->3	e->2	f->2	i->7	k->1	m->3	p->2	s->8	u->5	v->2	å->1	
åzon 	o->1	
ça Mo	u->5	
çois 	M->1	
ère k	o->1	
ète s	o->1	
ève 1	9->1	
ève, 	å->1	
èveko	n->1	
é - f	å->1	
é - o	c->1	m->1	
é att	 ->2	
é ave	c->1	
é ell	e->1	
é för	 ->3	
é har	 ->1	
é jag	 ->1	
é kom	m->1	
é med	 ->1	
é och	 ->3	
é om 	h->1	
é per	i->1	
é som	 ->5	
é uta	n->1	
é är 	a->1	
é, me	n->1	
éavta	l->1	
ébeto	n->1	
ébé a	v->1	
échar	d->1	
ée, v	i->1	
éer a	n->1	
éer i	 ->1	n->1	
éer m	å->1	
éer o	m->2	
éer s	k->1	o->2	
éer t	i->1	
éer, 	e->1	s->1	u->1	
éer.D	e->1	
éerna	 ->5	,->1	s->1	
éfére	n->1	
éförf	a->2	
ékonv	e->1	
én (C	E->2	
én at	t->6	
én ba	k->1	
én be	s->1	
én bö	r->1	
én fö	r->3	
én i 	e->1	
én ko	m->1	
én la	g->1	
én me	d->1	
én oc	h->4	
én om	 ->11	
én sa	d->1	
én si	n->1	
én va	d->1	
én vi	l->1	
én är	 ->1	
én, k	o->1	
én, o	c->1	
én, s	o->1	
én, u	t->1	
én, v	i->1	
én.Hu	r->1	
én.Me	n->1	
én.Wo	r->1	
én?Vi	l->1	
éns a	n->2	
éns g	e->6	
éns r	a->2	
éns s	a->1	
érend	a->1	
érys 	o->1	
és Ru	i->1	
ésyst	e->2	
étain	,->1	
éunio	n->2	
ête o	c->3	
êts (	u->1	
í är 	i->1	
íez G	o->1	
íncip	e->1	
ón Cr	e->2	
ón i 	C->1	
ón ti	l->1	
ón vi	s->1	
ónio 	V->1	
ône-A	l->1	
ö för	 ->2	
ö i d	e->1	
ö i e	n->1	
ö kan	 ->1	
ö mot	 ->1	
ö sak	n->1	
ö som	 ->1	
ö vin	n->1	
ö!Det	 ->1	
ö, fo	l->7	
ö, fö	r->1	
ö, hä	l->1	
ö, li	v->1	
ö, sm	å->1	
ö, up	p->1	
ö- oc	h->2	
ö.Det	 ->2	t->1	
ö.Då 	k->1	
ö.Men	 ->1	
ö.Und	e->1	
ö.Vil	k->1	
öanpa	s->1	
öansv	a->2	
öar s	o->1	
öarna	 ->2	,->1	.->1	s->1	
öavta	l->1	
öbela	s->1	
öbesk	a->1	
öbest	ä->1	
öbler	 ->1	i->1	
öbo v	i->1	
öbrot	t->1	
öcker	 ->1	,->2	
öd - 	e->1	v->1	
öd an	t->1	
öd av	 ->3	s->1	
öd bi	d->1	
öd de	 ->1	t->1	
öd dä	r->1	
öd ef	f->1	
öd en	l->2	
öd fr	å->7	
öd fö	r->20	
öd ge	n->1	
öd ha	r->1	
öd ho	s->1	
öd i 	E->2	h->1	k->1	l->1	t->1	
öd ib	l->1	
öd in	 ->1	n->1	o->2	t->1	
öd ka	n->4	
öd ko	m->1	
öd lö	p->1	
öd me	d->2	
öd må	s->3	
öd oc	h->14	
öd om	 ->4	
öd pe	r->1	
öd pr	i->1	
öd på	 ->5	
öd sk	u->1	
öd so	m->18	
öd så	 ->1	
öd ti	l->43	
öd va	d->1	r->1	
öd vi	 ->2	d->1	s->1	
öd än	 ->2	
öd åt	 ->2	
öd ök	a->1	
öd, d	e->1	
öd, e	f->1	
öd, m	i->1	
öd, o	c->2	m->1	
öd, s	o->3	p->1	t->2	å->1	
öd, u	t->1	
öd."J	a->1	
öd.- 	(->1	
öd..(	D->1	
öd.Al	l->1	
öd.At	t->1	
öd.De	n->2	t->8	
öd.Dä	r->1	
öd.Då	 ->1	
öd.Eu	r->1	
öd.Fö	r->2	
öd.Ha	d->1	
öd.He	r->4	
öd.I 	d->1	v->1	
öd.Ja	g->3	
öd.Me	n->1	
öd.Mo	t->1	
öd.Ni	 ->1	
öd.Or	d->1	
öd.Re	g->1	
öd.Så	 ->1	
öd.Tr	o->1	
öd.Ut	g->1	
öd.Vi	 ->2	
öd.Än	d->1	
öd.Äv	e->1	
öd.Å 	a->1	
öd.År	 ->1	
öd; d	e->1	
öd?- 	(->1	
öda o	c->1	s->2	
öda s	i->1	
öda t	r->2	
öda" 	b->1	
öda, 	ä->1	
ödade	 ->2	s->1	
ödand	e->5	
ödas 	i->1	
ödas,	 ->1	
ödats	 ->1	
ödbed	d->1	
ödd.M	e->1	
ödde 	V->1	
öddes	 ->2	
öde i	 ->1	
öde u	t->1	
öde, 	b->1	d->1	h->1	v->1	
öde.D	e->1	
öde?H	e->1	
ödela	g->1	
ödels	d->1	e->4	
ödema	r->1	
öden 	b->1	d->1	f->1	i->5	k->2	m->4	o->1	p->1	t->6	ö->1	
öden,	 ->2	
öden.	A->1	F->1	H->1	L->1	
ödena	 ->1	
ödens	 ->4	
ödepa	r->1	
öder 	E->1	U->1	a->3	d->15	e->1	f->1	g->1	h->5	i->5	j->2	k->3	l->1	m->2	p->1	r->4	s->3	t->1	v->8	ä->1	
öder,	 ->1	
öder.	U->1	
öderm	a->2	
ödesb	e->1	
ödesd	i->2	
ödesg	e->1	
ödet 	-->1	a->1	b->3	f->5	i->1	o->1	p->3	s->1	t->11	u->1	ä->1	
ödet,	 ->1	
ödet.	I->1	T->1	
ödets	 ->2	
ödföd	d->1	
ödgrö	n->1	
ödig 	b->1	f->1	
ödig.	E->1	
ödiga	 ->3	
ödigt	 ->6	,->1	
ödins	a->1	
ödire	k->1	
ödja 	-->1	D->1	H->1	a->1	d->28	e->4	f->4	i->1	k->4	l->1	m->1	o->3	p->1	r->1	s->4	u->1	v->1	Ö->1	å->3	
ödja.	H->1	J->1	
ödjas	 ->5	,->2	
ödjer	 ->1	
ödmed	l->1	
ödmot	t->1	
ödnin	g->1	
ödniv	å->1	
ödor.	K->1	
ödosa	m->1	
ödoäm	n->1	
ödpol	i->1	
ödra 	E->1	L->2	a->1	d->2	
ödram	 ->1	a->1	
ödrar	 ->1	
öds a	v->5	
öds b	l->1	
öds e	f->1	
öds g	e->1	
öds j	u->1	
öds t	r->1	
ödsdö	m->1	
ödsfa	l->1	
ödsit	u->1	
ödspo	l->1	
ödsys	t->4	
ödvän	d->125	
ödåtg	ä->5	
öende	 ->1	
öer f	ö->1	
öer i	 ->1	
öer s	a->1	
öerna	.->1	
öfakt	o->1	
öfarl	i->1	
öfart	,->1	s->7	
öfråg	o->4	
öfte 	d->1	i->1	s->1	
öften	 ->5	.->3	
öförb	ä->1	
öförh	å->1	
öförs	t->2	
ög ar	b->1	
ög be	v->1	
ög fe	l->1	
ög gr	a->6	
ög in	t->1	
ög kv	a->1	
ög ni	v->2	
ög pr	e->1	o->1	
ög se	i->1	
ög sk	y->1	
ög so	c->1	
ög st	a->2	
ög sy	s->1	
ög, d	e->1	
öga f	ö->1	
öga g	r->1	
öga k	o->1	r->2	
öga m	e->1	
öga n	i->1	
öga p	r->1	
öga r	e->2	ä->1	
öga s	k->1	
öga t	j->1	r->1	
öga å	t->2	
öga, 	i->1	
öga.M	e->1	
ögakt	u->1	
ögat.	V->1	
öge k	o->1	
öge r	e->1	
ögelm	e->1	
öger 	o->1	s->1	
öger,	 ->1	
ögere	x->6	
ögerm	a->1	
ögern	 ->7	,->2	.->3	s->7	
ögerp	o->1	
ögerv	r->1	
öghet	 ->1	,->1	.->1	
öglju	d->1	
ögna 	a->1	
ögniv	å->3	
ögon 	b->1	e->1	h->1	p->1	ä->1	
ögon,	 ->1	
ögonb	l->13	
ögra 	h->1	
ögre 	b->1	c->1	g->3	i->1	n->1	o->1	p->1	s->3	t->3	u->2	ä->1	
ögre.	D->1	
ögsko	l->1	
ögst 	a->2	b->1	g->1	k->2	o->1	p->1	r->1	t->1	u->1	
ögst,	 ->1	
ögsta	 ->16	
ögt f	ö->1	
ögt i	 ->1	n->1	
ögt p	r->3	
ögt s	a->1	
ögt u	p->1	
ögt v	ä->1	
ögt, 	o->1	
ögt.S	e->1	
ögtek	n->2	
ögtid	l->4	
öinfo	r->1	
öja J	ö->1	
öja d	e->4	
öja f	ö->1	
öja k	o->1	
öja l	e->1	
öja m	i->1	
öja o	s->5	
öja s	i->2	
öja t	i->1	
öja.V	i->1	
öjade	 ->1	
öjakt	i->2	
öjand	e->2	
öjar 	d->1	e->2	
öjare	 ->1	
öjas.	M->2	N->1	
öjd -	 ->1	
öjd a	t->1	
öjd g	a->1	
öjd m	e->1	
öjd p	å->1	
öjd s	ä->1	
öjd u	t->1	
öjda 	m->6	
öjda,	 ->3	
öjde 	b->1	s->1	
öjden	 ->1	
öjder	n->3	
öjdpu	n->2	
öje B	a->1	
öje E	u->1	
öje f	ö->1	
öje o	c->1	
öjels	e->1	
öjer 	j->1	l->1	m->2	s->1	
öjet 	a->2	
öjevä	c->3	
öjlig	 ->8	.->2	a->31	e->6	g->12	h->131	t->119	
öjnin	g->2	
öjor.	F->1	
öjs t	i->1	
öjsmå	l->2	
öjt o	s->1	
öjt s	i->1	
öjts 	t->1	
öjts,	 ->1	
ök at	t->4	
ök be	t->1	
ök i 	A->1	K->1	L->1	W->1	r->1	
ök om	 ->1	
ök so	m->1	
ök, d	e->1	
ök, o	c->1	
ök, s	o->1	
öka F	l->1	
öka a	l->3	n->7	r->1	
öka b	e->1	i->1	u->1	
öka d	e->4	
öka e	f->1	r->1	t->1	
öka f	a->1	i->1	r->1	å->2	ö->7	
öka g	e->2	
öka h	a->1	i->1	u->1	
öka i	 ->1	n->1	
öka j	ä->1	
öka k	o->4	v->3	ä->1	
öka m	i->1	y->1	ö->2	
öka o	c->1	m->2	
öka s	a->1	e->1	i->3	y->3	
öka t	r->1	
öka u	n->5	
öka v	a->3	ä->1	
öka å	t->1	
öka, 	m->1	
öka.O	c->1	
öka.R	å->1	
öka.T	a->1	
ökad 	a->4	d->1	e->1	f->2	i->2	j->1	k->4	p->3	s->7	t->1	u->1	ö->1	
ökade	 ->9	
ökand	e->11	
ökar 	1->1	a->1	d->1	e->1	f->1	i->3	m->1	n->1	o->1	v->1	
ökar,	 ->3	
ökar.	D->1	
ökarl	a->1	ä->5	
ökas 	e->1	i->1	o->1	t->1	u->1	
ökas,	 ->2	
ökas.	D->1	H->1	I->1	
ökast	a->1	
ökat 	a->3	d->1	e->1	h->1	i->3	m->2	o->1	s->1	u->1	y->1	ä->1	
ökat.	D->1	
ökata	s->10	
öke d	y->1	
öke.M	e->1	
öken 	a->1	t->1	
öker 	E->1	a->2	b->1	e->1	i->1	m->2	n->1	s->3	t->1	u->2	v->4	ä->1	ö->1	
öket 	a->2	m->1	p->1	
ökmod	e->1	
öknin	g->43	
ökonf	e->1	
ökons	e->5	
ökrav	 ->4	,->1	e->3	
öks, 	d->1	
öksbo	r->1	
ökstä	d->1	
ökt F	r->1	
ökt a	n->1	t->4	
ökt b	a->1	
ökt d	e->1	
ökt e	r->1	
ökt f	å->1	
ökt h	u->1	
ökt o	m->1	
ökt u	p->1	
ökt v	i->1	
ökte 	E->1	k->1	s->3	t->1	
ökval	i->1	
öl nä	r->1	
öl oc	h->1	
öl, s	å->1	
ölags	t->1	
ölar.	J->1	
öld m	i->1	
öld, 	m->1	
öldbe	s->1	
öldgr	ä->1	
ölja 	F->1	d->6	e->6	g->1	h->3	k->1	o->3	r->1	u->7	v->2	
ölja,	 ->1	
ölja.	M->1	
öljak	t->14	
öljan	d->37	
öljar	n->1	
öljas	 ->5	,->1	
öljd 	a->18	
öljd.	J->1	
öljde	 ->3	r->16	s->2	
öljdr	i->1	
öljds	k->2	
öljdå	t->1	
öljel	s->3	
öljer	 ->17	
öljni	n->10	
öljs 	a->1	k->1	u->2	
öljs,	 ->1	
öljt 	i->1	v->1	
öljts	 ->2	
öll K	i->1	
öll a	l->2	r->1	
öll d	e->2	ä->1	
öll e	l->1	n->3	
öll i	 ->2	
öll m	å->1	
öll n	ä->1	
öll o	c->2	
öll s	i->1	
öll t	i->1	
öll ö	v->1	
öll.H	a->1	
ölls 	a->1	d->1	i->1	p->1	
öln a	t->1	
öln i	 ->1	
öm av	 ->2	
öm be	r->1	
öm in	t->1	
öm ta	n->1	
öm, s	o->1	
öm: N	ä->1	
öma H	a->2	
öma a	l->2	v->1	
öma d	e->4	
öma e	n->2	
öma f	r->1	ö->1	
öma h	a->1	u->1	
öma i	 ->1	
öma o	m->2	s->1	
öma p	å->1	
öma r	i->1	
öma s	i->1	o->1	
öma t	y->1	
öma v	a->1	i->1	
öma, 	s->1	
öma.D	e->1	
ömand	e->7	
ömas 	b->1	p->1	
ömbar	a->1	
ömd, 	e->1	h->1	
ömde.	D->1	
ömdes	 ->1	
öme.K	o->1	
ömer 	J->2	a->1	f->2	o->2	p->1	s->1	
ömesg	i->1	
ömini	s->1	
ömlig	a->2	
ömma 	-->1	a->5	b->3	d->4	o->1	p->1	
ömma:	 ->1	
ömman	d->3	
ömmar	 ->1	,->1	n->1	
ömmas	 ->1	
ömmen	 ->1	,->2	.->1	
ömmer	 ->5	
ömnin	g->34	
öms e	f->2	
öms v	a->1	
ömses	i->5	
ömska	n->1	
ömt A	u->1	
ömt W	a->1	
ömt a	t->1	
ömt b	a->1	i->1	o->1	
ömt e	t->1	
ömt p	a->1	
ömt s	i->1	
ömt v	a->1	
ömts 	a->1	i->1	
ömtål	i->1	
ömvär	d->1	
ömän 	e->1	s->1	
ömäss	i->11	
ömål 	o->1	ä->1	
ömåls	ä->1	
ön No	i->1	
ön el	l->1	
ön en	 ->1	
ön fö	r->2	
ön hå	l->1	
ön i 	s->1	
ön oc	h->6	
ön på	 ->1	
ön so	m->2	
ön ti	l->1	
ön vä	n->2	
ön är	 ->1	
ön!De	n->1	
ön, a	t->1	
ön, d	e->1	
ön, h	a->1	
ön, m	e->1	
ön, o	c->3	
ön, s	k->1	
ön, u	t->1	
ön.De	n->1	t->1	
ön.Dä	r->1	
ön.En	 ->1	
ön.Fr	u->1	
ön.Ja	g->1	
ön.Lå	t->1	
ön.Ma	n->1	
ön.Un	i->1	
ön.Vi	 ->1	
ön.Vå	r->1	
öna e	l->1	
öna f	ö->1	
öna g	e->1	l->1	
öna h	a->2	
öna i	n->1	
öna m	ä->1	
öna n	ä->1	
öna o	c->1	
öna p	o->1	
öna s	t->1	ä->1	
öna/E	u->1	
önar 	d->1	
önare	.->1	
önas 	f->1	m->1	
önas,	 ->1	
önbok	 ->1	
önder	 ->2	.->1	d->4	
öne- 	o->1	
önear	b->1	
önen 	(->1	-->1	E->1	
öner 	o->1	s->1	
önhet	.->1	
önitz	 ->1	
önk h	o->1	
önk r	a->1	
önk u	t->1	
önk.D	e->1	
önorm	e->2	
öns f	l->1	
öns s	k->1	
önsam	 ->2	m->2	t->1	
önsgr	u->1	
önska	 ->11	.->2	d->4	n->13	r->20	t->4	
önske	m->3	
önskn	i->2	
önskv	ä->10	
önste	r->2	
önstr	e->1	
önt a	t->1	
önt l	j->1	
öntag	a->3	
öområ	d->4	
öovän	l->1	
öp av	 ->2	
öpa d	e->1	
öpa e	n->1	
öpa u	t->1	
öpand	e->6	
öpare	 ->1	,->1	.->1	
öparn	a->1	
öpenh	a->1	
öper 	E->1	d->2	e->2	o->1	r->3	u->3	
öper.	F->1	
öpers	p->1	
öpkra	f->1	
öpoli	c->1	t->7	
öppen	 ->6	h->59	
öppet	 ->13	.->1	
öppna	 ->8	,->2	d->1	r->3	s->2	
öppni	n->4	
öprob	l->3	
öprog	r->1	
öpsbe	s->1	
öpsla	g->1	
öpt i	 ->1	
öpt u	t->5	
öpte 	d->1	u->2	
öpåve	r->1	
ör "K	u->1	
ör "a	n->2	
ör "f	o->1	
ör "i	n->1	
ör "n	a->1	
ör - 	a->3	h->1	s->1	v->1	
ör -,	 ->1	
ör 19	9->17	
ör 20	 ->2	0->3	
ör 27	 ->1	
ör 29	 ->1	
ör 3 	0->1	
ör 33	 ->1	
ör 5 	m->1	
ör 5,	8->1	
ör 75	 ->1	
ör 76	 ->1	
ör 81	 ->1	
ör Ag	r->1	
ör Al	t->3	
ör Be	l->1	
ör Bi	s->1	
ör Bo	u->1	
ör Br	e->3	
ör CS	U->1	
ör Ce	n->1	
ör Da	n->2	
ör De	u->1	
ör EC	H->1	
ör EG	-->4	
ör EU	 ->1	,->1	-->1	.->2	:->4	
ör Er	i->1	
ör Eu	r->60	
ör FP	Ö->1	
ör Fo	U->1	l->1	
ör Fö	r->2	
ör Ge	n->1	
ör Go	l->1	
ör Ha	i->1	
ör IM	O->1	
ör IN	T->1	
ör In	t->1	
ör Is	r->1	
ör Ka	n->3	
ör Ko	s->1	
ör Ku	l->2	
ör Ky	o->1	
ör La	n->1	
ör Le	i->1	
ör Mo	r->1	
ör OL	A->1	
ör PP	E->1	
ör Pa	c->1	
ör Po	r->2	
ör Sa	v->2	
ör Sã	o->1	
ör Ta	c->1	
ör Ti	b->6	
ör Tu	r->1	
ör Vo	l->1	
ör WT	O->1	
ör Wa	l->1	
ör ab	s->2	
ör ac	c->1	
ör ai	d->1	
ör al	l->141	
ör am	b->2	
ör an	d->4	g->1	n->8	s->23	t->5	v->5	
ör ar	b->12	r->1	t->2	
ör as	y->3	
ör at	t->778	
ör av	 ->3	f->2	g->1	s->17	t->1	u->1	v->1	
ör ba	k->1	r->2	
ör be	a->1	d->5	f->5	g->6	h->7	k->4	m->1	r->7	s->3	t->3	v->2	
ör bi	d->1	l->5	s->5	
ör bj	u->1	
ör bl	.->1	a->1	i->3	y->1	
ör bo	m->1	s->1	t->1	
ör br	o->4	
ör bu	d->13	s->1	
ör bä	t->1	
ör bå	d->3	
ör bö	r->6	
ör ce	n->2	
ör ch	o->1	
ör ci	r->1	v->3	
ör da	g->3	n->1	
ör de	 ->132	b->1	c->1	f->1	l->1	m->27	n->180	r->14	s->24	t->303	
ör di	r->2	s->9	
ör dj	u->1	
ör do	c->2	k->1	m->1	
ör du	 ->2	
ör dä	r->7	
ör då	 ->2	l->2	
ör dö	r->1	
ör ef	f->1	
ör eg	e->4	
ör ek	o->16	
ör el	e->2	l->3	
ör em	e->1	
ör en	 ->136	b->1	d->1	e->6	l->1	o->1	s->3	
ör er	 ->12	,->5	.->2	a->4	i->2	k->2	t->7	
ör et	t->57	
ör eu	r->1	
ör ev	i->2	
ör ex	p->1	t->2	
ör fa	c->1	n->1	r->7	s->2	
ör fe	l->1	m->2	
ör fi	n->7	s->5	
ör fj	o->1	
ör fl	e->3	y->1	ä->1	
ör fo	d->3	l->2	r->5	
ör fr	a->7	e->5	i->9	ä->5	å->7	
ör fu	l->1	n->2	
ör fy	s->1	
ör få	 ->5	,->1	.->1	r->1	
ör fö	l->2	r->66	
ör ga	n->1	
ör ge	 ->1	m->8	n->14	
ör gi	v->3	
ör gl	ä->1	
ör go	d->4	
ör gr	a->5	u->8	ä->3	
ör gu	d->2	
ör gä	r->1	
ör gö	r->8	
ör ha	 ->5	n->28	r->6	
ör he	l->11	m->5	n->7	
ör hi	s->1	
ör hj	ä->3	
ör ho	n->4	p->1	t->1	
ör hu	m->1	n->1	r->9	v->1	
ör hä	l->3	n->2	r->4	s->1	
ör hå	l->2	r->1	
ör hö	g->4	j->1	
ör i 	E->1	a->2	d->6	e->1	f->2	g->1	p->2	s->3	Ö->1	
ör ic	k->1	
ör ih	o->2	
ör ik	r->1	
ör il	l->1	
ör in	 ->1	d->9	f->5	g->4	i->1	k->1	n->5	r->3	s->6	t->24	v->3	
ör ja	g->14	
ör jo	r->11	
ör ju	 ->1	r->2	s->1	
ör jä	m->2	r->1	
ör ka	l->1	m->3	n->11	p->1	r->1	t->2	
ör kl	a->1	
ör kn	a->1	
ör ko	l->2	m->58	n->34	r->4	s->6	
ör kr	a->3	i->2	ä->5	
ör ku	l->19	n->2	s->2	
ör kv	a->1	e->2	i->6	
ör kä	n->1	r->5	
ör la	g->3	n->4	s->2	
ör le	d->3	
ör li	k->4	t->8	v->16	
ör lo	b->1	g->1	k->1	
ör lä	g->4	n->10	s->1	
ör lå	n->7	
ör lö	n->1	
ör ma	n->32	r->1	t->1	
ör me	d->46	l->1	n->2	r->2	t->1	
ör mi	g->19	l->21	n->18	t->2	
ör mo	t->6	
ör my	c->15	
ör mä	n->14	
ör må	l->4	n->11	s->14	
ör mö	j->3	
ör na	m->1	r->1	t->9	
ör ne	d->2	
ör ni	 ->2	
ör no	r->6	t->3	
ör nu	 ->2	.->1	
ör ny	 ->1	a->6	
ör nä	r->39	s->3	
ör nå	g->19	
ör nö	d->3	
ör oc	h->10	k->9	
ör of	f->2	t->11	
ör ol	i->2	j->2	y->1	
ör om	 ->4	f->5	r->5	
ör op	i->1	
ör or	d->6	s->1	
ör os	s->55	t->1	
ör ot	r->1	
ör ov	a->1	ä->1	
ör pa	r->23	
ör pe	n->4	r->21	s->1	
ör pl	a->1	
ör po	l->5	t->1	
ör pr	e->2	i->2	o->15	
ör pu	n->1	
ör på	 ->4	t->1	
ör ra	m->1	s->1	
ör re	a->2	f->4	g->39	h->1	k->2	l->2	p->1	s->5	t->1	v->3	
ör ri	s->4	
ör ro	s->1	
ör rä	k->1	t->27	
ör rå	d->9	
ör rö	r->1	s->5	
ör sa	k->1	m->13	t->2	
ör se	 ->4	d->1	n->4	x->1	
ör si	g->21	n->21	s->4	t->8	
ör sj	ä->5	
ör sk	a->9	e->1	i->1	o->4	r->3	u->9	y->3	ä->1	
ör sl	ä->2	
ör sm	å->5	
ör sn	a->4	
ör so	c->2	m->3	
ör sp	e->1	r->2	ä->1	
ör st	a->10	e->2	o->16	r->9	u->2	y->1	ä->1	å->3	ö->15	
ör sv	a->3	
ör sy	d->1	s->19	
ör sä	g->1	k->15	l->1	
ör så	 ->4	d->5	v->4	
ör t.	e->2	
ör ta	 ->3	g->1	l->1	n->2	
ör te	k->2	
ör ti	b->1	d->3	l->49	
ör tj	u->1	ä->6	
ör to	b->1	
ör tr	a->19	e->3	o->3	y->1	
ör tu	n->1	r->2	
ör tv	i->2	u->1	ä->1	å->4	
ör ty	c->1	d->2	n->1	
ör tå	g->1	
ör un	d->10	g->4	i->26	
ör up	p->12	
ör ur	 ->2	
ör ut	 ->1	a->1	b->4	e->2	f->5	g->3	n->1	r->4	s->25	t->3	v->18	
ör va	d->6	k->1	r->32	
ör ve	r->7	t->5	
ör vi	 ->38	d->6	k->2	l->17	n->1	r->1	s->8	t->3	
ör vo	t->1	
ör vu	x->1	
ör vä	l->4	n->1	
ör vå	r->43	
ör yn	g->1	
ör yr	k->1	
ör yt	t->2	
ör Ös	t->2	
ör äg	n->1	
ör än	 ->1	d->5	n->2	
ör är	 ->26	
ör äv	e->4	
ör åk	l->1	
ör år	 ->10	e->2	
ör åt	 ->1	a->2	e->19	g->4	
ör öa	r->1	
ör ög	o->7	
ör ök	a->3	
ör öp	p->5	
ör ör	e->1	
ör ös	t->1	
ör öv	e->7	r->27	
ör".O	m->1	
ör, 1	6->1	
ör, B	u->1	
ör, a	t->6	
ör, e	f->1	n->1	
ör, f	r->2	ö->1	
ör, h	e->1	
ör, i	 ->2	
ör, k	o->3	
ör, m	i->1	
ör, o	c->4	
ör, s	o->2	å->1	
ör, t	r->1	
ör, u	t->1	
ör, v	a->1	
ör, ä	r->1	v->1	
ör. D	e->1	
ör. E	n->1	
ör.(L	i->1	
ör...	(->1	
ör.De	t->6	
ör.Di	r->1	
ör.Et	t->1	
ör.Fö	r->1	
ör.He	r->1	
ör.Ja	g->1	
ör.Ko	m->1	
ör.Ma	n->1	
ör.Me	n->2	
ör.Vi	 ->4	
ör.Vå	r->1	
ör: D	e->1	
ör: F	i->1	
ör: a	t->1	
ör; d	e->1	
ör?Dä	r->1	
ör?Fr	u->1	å->1	
ör?I 	m->1	
ör?Är	 ->1	
öra -	 ->1	
öra E	U->1	u->2	
öra a	f->1	g->1	l->8	n->2	r->1	t->11	v->3	
öra b	a->1	e->6	
öra d	e->98	i->2	y->1	
öra e	g->1	n->50	r->3	t->18	
öra f	l->1	o->1	r->4	ö->18	
öra g	a->1	e->4	r->2	ä->1	
öra h	a->1	e->1	o->1	u->2	ä->1	
öra i	 ->7	n->5	
öra k	l->6	o->7	v->1	
öra l	a->2	i->2	ä->1	
öra m	a->1	e->24	i->11	o->1	y->2	ä->1	å->1	
öra n	a->1	e->1	u->1	y->2	ä->1	å->19	
öra o	c->3	m->4	
öra p	a->2	o->2	r->4	å->2	
öra r	e->5	ö->1	
öra s	a->3	i->20	j->1	k->1	l->1	o->3	t->5	y->2	å->2	
öra t	a->1	i->4	r->3	v->2	
öra u	n->4	p->8	r->1	t->3	
öra v	a->7	i->5	å->3	
öra y	t->2	
öra ä	n->1	r->4	
öra å	t->2	
öra ö	k->1	v->1	
öra, 	a->1	f->1	h->1	k->1	m->1	o->2	v->1	å->1	
öra.D	e->4	ä->1	
öra.E	G->1	n->1	
öra.H	e->1	
öra.I	n->1	
öra.J	a->4	
öra.L	å->1	
öra.N	a->1	
öra.O	c->1	
öra.P	e->1	
öra.S	ä->1	
öra?J	a->1	
örakt	a->1	
örall	t->1	
örand	e->389	
örank	r->4	
öranl	e->2	
örans	l->1	
örarb	e->1	
örarl	ä->1	
örarn	a->1	
öras 	a->3	b->2	e->2	f->5	g->1	h->1	i->5	j->2	k->1	m->7	n->3	o->3	r->3	s->5	t->4	u->6	v->3	å->1	ö->3	
öras!	D->1	G->1	
öras,	 ->5	
öras.	A->1	B->1	D->3	G->2	I->1	J->1	M->2	N->1	U->1	V->3	
öras;	 ->1	
örban	d->2	
örbar	 ->2	.->1	a->5	m->1	t->3	
örbeh	å->6	
örber	e->27	
örbi 	d->1	
örbif	a->2	
örbig	å->6	
örbin	d->22	
örbis	e->1	
örbju	d->14	
örble	v->1	
örbli	 ->8	r->6	
örbru	k->1	
örbry	t->2	
örbrä	n->2	
örbud	 ->11	,->2	.->3	e->8	s->2	
örbun	d->12	
örbät	t->78	
örd a	r->1	v->1	
örd f	r->1	
örd k	a->1	
örd m	i->1	
örd o	c->1	
örd, 	s->1	
örd.D	e->1	ä->1	
örda 	a->3	d->1	e->1	f->2	k->5	l->2	m->3	n->1	o->1	p->5	s->4	u->1	
örda,	 ->2	
örda.	D->1	H->2	
örda?	D->1	
ördad	e->2	
ördag	 ->1	
ördan	 ->5	.->3	d->1	
ördar	e->1	
ördat	 ->1	s->1	
örde 	K->1	a->1	e->3	g->1	i->3	j->2	k->1	m->1	n->1	p->1	r->1	s->1	t->1	v->1	
örde,	 ->1	
örde.	J->1	L->1	
ördel	 ->3	,->2	.->2	a->13	e->1	n->21	
örden	 ->6	.->1	
ördes	 ->9	,->1	.->1	
ördhe	t->1	
ördju	p->11	
ördna	d->1	
ördom	a->1	s->1	
ördor	 ->1	n->1	
ördra	g->164	
ördrö	j->1	
ördub	b->2	
ördun	k->1	
ördär	v->4	
ördöm	a->13	e->5	t->2	
öre 2	0->1	
öre A	m->1	
öre K	i->1	
öre d	e->5	
öre e	n->1	
öre m	a->1	e->1	i->1	
öre n	ä->2	
öre o	c->1	m->1	s->1	
öre s	l->1	t->1	
öre u	t->4	
öre v	a->2	
öre å	t->1	
öre ö	v->1	
örebi	l->1	
örebr	å->2	
öreby	g->23	
öredr	a->165	o->1	
öredö	m->2	
örefa	l->20	
örefö	l->1	
öregi	c->1	o->7	
öregr	i->1	
öregå	e->15	n->2	
öreha	v->1	
öreko	m->22	
örele	g->1	
öreli	g->26	
örels	e->21	
öremå	l->13	
ören 	o->1	
ören,	 ->1	
örena	 ->8	d->16	r->1	
öreni	n->12	
örenk	l->8	
örenl	i->9	
örens	 ->1	
örent	a->28	
örer 	h->1	o->2	s->3	
örer,	 ->3	
örer.	D->3	P->1	
örern	a->10	
öresa	t->6	
öresk	r->28	
öresl	a->24	o->11	å->69	
öresp	e->1	r->9	
örest	ä->9	å->6	
öresä	t->1	
öreta	,->2	g->198	
öretr	ä->73	
örfal	s->1	
örfar	a->76	
örfat	t->7	
örfin	i->1	
örfjo	l->1	
örflu	t->14	
örfly	t->4	
örfog	a->18	
örfry	s->1	
örfrå	g->4	
örfäk	t->1	
örfär	a->1	l->1	
örfån	g->1	
örföl	j->5	
örg H	a->14	
örglö	m->2	
örgru	n->3	
örgäv	e->1	
örhan	d->92	
örhas	t->3	
örhin	d->31	
örhop	p->12	
örhål	l->56	
örhöl	l->1	
örig 	i->1	p->1	
öriga	 ->2	
örigh	e->15	
örigt	 ->1	.->1	
öring	 ->6	,->3	;->1	a->1	e->5	
örint	e->5	
örirr	a->1	
örja 	a->7	d->1	e->2	f->8	k->2	m->37	o->1	p->3	r->1	s->1	t->3	u->1	å->1	
örjad	e->8	
örjan	 ->17	,->2	
örjar	 ->16	.->1	
örjat	 ->9	.->2	s->1	
örjde	 ->1	
örjer	 ->2	
örjni	n->4	
örk d	a->1	
örkas	t->9	
örkla	r->76	
örklä	g->1	
örkni	p->3	
örkor	t->2	
örkro	m->1	
örkun	n->2	
örlag	e->1	o->2	
örleg	a->2	
örlig	 ->7	.->1	a->2	e->1	h->24	t->4	
örlik	a->1	n->44	
örlin	g->1	
örlis	t->2	
örlit	a->6	l->4	
örliv	a->19	
örlor	a->20	
örlus	t->10	
örläg	g->2	
örlän	g->4	
örlåt	a->1	e->1	l->2	
örmed	l->3	
örmen	a->2	
örmid	d->3	
örmod	l->12	
örmyn	d->1	
örmå 	b->1	r->1	
örmåg	a->31	
örmån	 ->11	e->2	s->1	
örmår	.->1	
örmög	n->1	
örn d	ä->1	
örn f	ö->1	
örnam	n->1	
örned	r->2	
örnek	a->8	
örnin	g->7	
örnst	e->1	
örnuf	t->14	
örnya	 ->1	n->1	r->1	s->1	
örnyb	a->39	
örnye	l->6	
örolä	m->2	
öron,	 ->1	
öronm	ä->2	
örord	a->2	n->42	
örore	n->28	
örors	a->6	
örpac	k->5	
örpas	s->1	
örpli	k->21	
örr d	å->1	
örr e	l->2	
örr ö	p->1	
örr, 	i->1	m->1	
örra 	k->6	m->2	p->1	r->1	v->13	å->19	
örrar	 ->2	n->1	
örre 	-->2	a->6	b->4	d->3	e->2	f->4	h->2	i->2	j->2	k->1	l->2	m->3	o->5	p->4	r->4	s->8	t->1	u->8	v->6	ä->2	ö->6	
örren	 ->1	,->3	
örres	t->2	
örrgå	r->3	
örrin	g->1	
örräd	e->1	
örrän	 ->4	
örråd	e->1	
örs a	t->1	v->16	
örs b	a->1	
örs d	e->1	
örs e	n->4	t->2	
örs f	l->1	o->1	r->1	u->2	ö->2	
örs i	 ->8	
örs k	a->1	
örs m	e->2	
örs o	c->1	
örs p	å->5	
örs t	i->1	
örs u	n->1	
örs ä	r->1	
örs ö	v->2	
örs, 	a->1	f->2	i->1	k->1	m->1	o->1	
örs. 	E->1	
örs..	(->1	
örs.D	e->2	
örs.H	e->1	
örs.J	a->2	
örs.O	n->1	
örs.V	å->1	
örsam	l->12	
örse 	d->1	f->1	
örsen	 ->1	a->14	i->13	
örser	 ->1	n->1	
örses	 ->1	
örsik	t->67	
örska	p->2	
örski	n->2	
örskj	u->1	
örsko	n->1	t->1	
örskr	ä->4	
örskä	m->1	
örskå	r->1	
örsla	g->492	
örsom	r->1	
örson	a->1	i->4	
örspo	r->1	
örst 	a->8	d->2	e->4	g->2	h->2	i->4	k->1	m->3	n->2	o->23	r->3	s->11	t->3	u->1	v->6	
örst.	M->2	
örsta	 ->205	,->10	:->5	;->2	b->1	i->22	k->1	
örste	 ->1	
örstk	l->1	
örsto	d->3	
örstä	l->1	r->29	
örstå	 ->20	,->1	.->2	d->2	e->13	n->9	r->23	s->4	t->9	
örstö	r->21	
örsum	b->1	m->8	
örsva	g->21	r->41	
örsvi	n->15	
örsvu	n->4	
örsvå	r->2	
örsäk	r->44	
örsäl	j->5	
örsäm	r->10	
örsän	k->1	
örsåg	s->1	
örsök	 ->5	,->2	a->22	e->18	t->14	
örsör	j->4	
ört -	 ->2	
ört D	u->1	
ört a	r->1	
ört d	e->4	y->1	
ört e	k->1	n->2	r->2	t->2	
ört f	a->1	r->4	ö->1	
ört i	 ->2	n->1	
ört k	l->1	
ört l	i->1	
ört m	e->10	y->1	å->1	
ört n	y->1	å->1	
ört o	m->1	s->1	
ört p	o->2	å->1	
ört s	a->2	i->1	t->1	v->1	y->1	
ört t	a->2	
ört u	n->2	
ört v	i->1	å->1	
ört, 	h->2	t->1	
ört.J	a->1	
ört.K	o->1	
örtec	k->3	
örtid	s->6	
örtju	s->1	
örtjä	n->20	
örtni	n->1	
örtro	e->56	g->1	s->2	t->1	
örtry	c->2	
örträ	f->2	n->1	
örtrö	t->1	
örts 	a->7	d->2	f->2	h->2	i->4	m->1	o->4	p->2	s->1	t->1	v->1	
örts,	 ->3	
örts.	D->1	S->1	T->1	V->1	
örtvi	v->1	
örtyd	l->3	
örtäc	k->1	
örund	e->1	
örut 	a->1	o->1	
örut.	D->1	
örutb	e->1	
öruto	m->15	
öruts	a->1	e->8	ä->54	
örutv	a->2	
örval	t->49	
örvan	d->4	s->2	
örvar	n->1	
örver	k->22	
örvir	r->12	
örvis	a->1	s->8	
örvrä	n->1	
örväg	 ->5	,->4	.->2	r->3	
örvän	t->29	
örvär	r->4	v->7	
örvån	a->6	
öränd	e->1	r->73	
öråde	t->1	
öråld	r->3	
öröda	n->3	
öröde	l->2	
öröre	l->2	
öröva	d->1	r->2	
ös - 	o->1	
ös da	g->1	
ös de	b->1	
ös en	 ->1	
ös kä	l->1	
ös oc	h->2	
ös po	l->1	
ös ra	m->1	
ös sk	o->1	
ös su	b->1	
ös ut	v->1	
ös, k	o->1	
ös.De	t->1	
ösa a	r->1	
ösa d	e->9	
ösa e	n->2	
ösa f	r->1	
ösa g	e->1	r->1	
ösa h	i->1	
ösa i	 ->1	
ösa k	o->2	
ösa m	a->1	e->2	o->1	å->4	
ösa n	å->1	
ösa o	c->2	r->1	
ösa p	r->7	å->1	
ösa r	e->1	
ösa s	i->2	k->1	t->1	
ösa u	n->1	p->1	
ösa v	a->1	e->1	i->2	
ösa, 	5->1	d->1	l->1	v->1	
ösa.A	n->1	
ösa.F	ö->1	
ösa.I	 ->1	
ösa.M	e->1	
ösar 	m->1	
ösare	 ->1	.->1	
ösas 	b->1	o->3	p->1	
ösas.	D->1	
ösekt	o->1	
öser 	i->1	
öseri	 ->2	.->1	
öses 	t->1	
ösgör	 ->1	
öshet	 ->10	,->3	.->3	e->25	s->3	
ösida	n->1	
öskad	l->2	
öskel	n->3	
öskyd	d->11	
öskäl	 ->1	.->1	
ösnin	g->52	
ösryc	k->1	
öss o	c->1	
öss p	å->1	
öss ä	r->1	
öss) 	o->1	
össor	,->1	
öst -	 ->2	
öst a	r->1	t->1	
öst d	e->1	r->1	
öst f	r->1	ö->1	
öst h	a->2	ö->1	
öst i	 ->2	n->2	
öst l	e->1	
öst m	e->1	
öst o	c->3	m->2	
öst p	l->1	r->1	
öst r	a->1	
öst s	o->1	ä->2	
öst t	i->2	
öst v	e->1	
öst, 	a->1	e->1	i->1	
öst.J	a->1	
öst.Ä	r->1	
östa 	d->1	e->6	f->26	h->1	i->3	m->3	o->4	p->2	v->1	
östa,	 ->1	
östa.	)->1	-->1	D->1	V->1	
östad	e->15	
östar	 ->15	
östat	 ->14	s->1	
östbl	o->1	
östed	t->4	
östen	 ->1	
öster	 ->1	,->2	n->20	r->49	
östes	 ->1	
östeu	r->3	
östfö	r->7	
östlä	n->1	
östni	n->57	
östra	 ->3	
östrä	t->3	
östs.	S->1	
östto	n->1	
östut	v->2	
östvi	k->3	
östöd	 ->1	
ösynp	u->6	
öt 93	 ->1	
öt at	t->1	
öt de	m->1	
öt ha	n->1	
öt lo	j->1	
öt ta	l->4	
öt vi	 ->1	
öt.De	 ->1	
öta E	u->1	
öta d	e->8	
öta e	t->1	
öta m	e->1	i->1	
öta p	å->1	
öta s	i->3	
öta v	e->1	
ötand	e->1	
ötar 	i->1	
ötas 	v->1	
öte d	ä->1	
öte i	 ->4	
öte k	o->1	
öte m	e->4	
öte o	c->1	
öte p	å->1	
öte s	ä->1	
ötebo	r->1	
öten 	m->1	o->1	
ötena	 ->2	
öter 	-->1	a->7	d->2	e->2	g->1	h->3	i->7	l->1	m->1	o->6	p->1	s->7	v->4	
öter!	 ->12	M->1	V->1	
öter,	 ->7	
öter.	D->1	
ötern	a->24	
öters	 ->1	
ötes 	m->1	
ötes.	K->1	
ötesg	å->3	
ötest	e->1	
ötet 	(->1	f->1	i->13	m->3	u->1	
ötet.	E->1	V->1	
ötfån	g->1	
ötköt	t->3	
ötran	s->1	
öts a	v->1	
öts b	e->1	
öts i	n->1	
öts k	l->2	
öts m	e->1	
öts.V	i->1	
ötsel	 ->4	.->1	
ötska	l->1	
ötsli	g->4	
ött B	e->1	
ött F	N->1	
ött d	e->2	
ött k	o->1	
ött o	c->1	
ött p	å->2	
ött s	i->1	o->1	t->1	
ött t	i->1	
ött u	t->1	
ött v	i->1	å->1	
ött ä	n->1	
ött.D	e->2	
ött.J	a->1	
ötta 	p->1	
ötta,	 ->1	
öttat	 ->2	
ötte 	d->1	o->1	
ötter	 ->4	,->1	n->3	
öttes	 ->1	
öttkr	i->1	
öttra	r->1	
ötts 	a->1	u->1	
ötts-	 ->1	
öttsp	r->1	
öutsk	o->1	
öva E	u->1	
öva a	v->1	
öva d	e->1	
öva e	n->3	
öva f	ö->1	
öva g	ö->3	
öva h	u->1	
öva k	l->1	o->1	
öva l	e->1	
öva n	å->1	
öva p	a->1	å->2	
öva r	å->1	
öva s	i->2	
öva t	v->1	
öva u	p->1	r->1	
öva v	å->1	
öva ö	k->1	
övade	 ->1	s->1	
övand	e->1	
övar 	d->1	e->1	o->1	s->2	
övare	n->2	
övas 	a->4	h->1	o->1	
övas.	C->1	H->1	V->1	
övat 	u->1	
övats	 ->1	
övde 	f->1	g->1	
över 	-->2	1->1	2->1	3->2	4->1	5->1	7->1	8->1	9->1	B->1	E->5	H->1	a->38	b->3	d->46	e->25	f->11	g->14	h->37	i->6	j->2	k->6	l->3	m->11	n->3	o->9	p->6	r->8	s->20	t->5	u->5	v->29	Ö->1	ä->4	å->1	
över,	 ->5	
över.	 ->1	D->2	H->1	M->1	O->1	S->2	T->1	V->1	
övera	l->9	
överb	e->4	l->1	r->4	
överc	e->1	
överd	r->14	
övere	n->71	
överf	a->3	i->1	l->3	ö->16	
överg	e->10	i->2	r->14	å->15	
överh	a->1	ä->1	ö->2	
överi	n->1	
överk	l->6	
överl	a->1	e->5	ä->21	å->8	
överm	o->2	
övern	a->3	i->1	
övero	r->1	
överp	r->1	
överr	a->1	e->2	ö->1	
övers	a->1	i->18	k->23	t->9	v->7	y->1	ä->11	
övert	a->6	o->2	r->7	y->38	ä->1	
överv	a->25	i->8	u->1	ä->37	
övitt	 ->1	
övlad	e->1	
övlig	a->1	
övnin	g->12	
övoår	 ->1	
övrad	e->1	
övran	d->1	
övrar	,->1	
övrig	 ->1	a->32	t->32	
övs d	e->3	
övs e	g->1	n->4	t->1	
övs f	ö->2	
övs i	 ->1	n->2	
övs m	y->1	
övs n	å->1	
övs o	c->1	
övs p	å->1	
övs s	ä->1	å->1	
övs, 	f->1	o->1	
övs.D	e->1	
övs.F	r->1	
övs.I	 ->1	
övs.S	a->1	l->1	
övsko	g->1	
övsta	 ->1	
övt f	ö->1	
övt s	t->1	
övt t	a->1	
övts 	d->1	
övänl	i->7	
övärd	e->2	i->1	
öw fö	r->1	
öy - 	s->1	
ööw f	ö->1	
øn, i	n->1	
øn, m	e->1	
ørgen	s->2	
ührko	p->1	
ünche	n->1	
ürkda	m->1	
üssel	 ->2	,->1	.->1	
