 	"->99	'->1	(->215	,->5	-->565	0->31	1->443	2->230	3->86	4->71	5->47	6->28	7->40	8->67	9->41	:->1	A->149	B->188	C->95	D->223	E->1104	F->214	G->99	H->152	I->175	J->191	K->193	L->130	M->135	N->60	O->47	P->176	Q->1	R->78	S->217	T->179	U->38	V->111	W->61	X->3	Y->2	Z->3	[->3	a->13183	b->4761	c->161	d->11542	e->7033	f->11742	g->3644	h->5121	i->8091	j->1522	k->6112	l->2384	m->8171	n->2924	o->9147	p->4785	q->4	r->3591	s->14142	t->5952	u->4024	v->6975	w->3	y->158	z->8	º->1	Ä->18	Å->7	Î->1	Ö->87	ä->3699	å->1117	ö->1078	
!	 ->374	"->4	(->1	.->3	A->5	D->21	E->5	F->5	G->1	H->11	I->1	J->18	K->1	L->2	M->9	N->4	O->2	P->1	R->1	S->2	T->6	U->1	V->5	Ä->2	
"	 ->38	!->1	)->1	,->23	.->29	;->1	A->2	B->1	D->6	E->4	I->1	J->4	K->7	L->1	M->3	O->3	P->1	T->3	U->1	a->8	b->1	c->1	d->6	e->9	f->2	g->2	h->2	i->4	j->1	k->4	l->3	m->1	n->4	o->3	p->2	r->6	s->5	t->1	u->2	v->2	å->1	ö->2	
'	V->1	e->1	
(	"->1	1->15	5->1	8->2	9->4	A->42	B->7	C->34	D->5	E->43	F->22	G->1	H->22	I->8	K->10	L->2	N->4	P->34	S->7	T->8	U->2	a->9	d->2	e->4	f->8	h->1	i->4	k->6	m->3	o->1	r->2	s->2	t->2	u->1	Ö->5	å->1	
)	 ->189	(->11	)->22	,->12	.->28	0->6	:->19	;->2	?->1	A->5	B->8	D->1	F->10	G->1	H->3	J->4	K->1	N->3	O->1	R->1	S->1	T->1	U->1	]->3	o->1	Å->1	
,	 ->6144	0->1	2->3	3->1	4->3	5->3	6->1	7->1	8->4	9->1	
-	 ->672	(->1	,->12	0->89	1->4	2->24	4->1	9->1	A->5	B->7	C->2	D->9	E->1	F->5	H->2	I->3	J->2	K->1	L->2	M->3	N->1	P->5	R->2	S->8	a->15	b->14	d->32	e->4	f->31	g->22	h->1	i->11	k->33	l->13	m->9	n->4	o->13	p->28	r->17	s->30	t->12	u->2	v->2	z->3	
.	 ->349	"->5	(->57	)->32	,->3	-->15	.->79	0->14	1->17	2->8	3->6	4->3	5->2	8->1	9->1	?->1	A->141	B->71	C->5	D->1567	E->268	F->370	G->43	H->378	I->277	J->786	K->172	L->77	M->388	N->157	O->201	P->102	R->59	S->242	T->129	U->67	V->683	W->1	Y->3	a->28	d->3	e->20	g->1	k->5	m->8	o->7	Ä->73	Å->24	Ö->9	
/	0->26	1->43	2->28	3->5	4->2	5->4	6->1	7->4	9->32	E->11	N->4	O->1	d->1	e->1	h->1	i->1	r->1	s->1	å->2	
0	 ->184	"->5	(->5	)->26	,->13	-->32	.->28	/->12	0->397	1->38	2->21	3->26	4->11	5->12	6->36	7->23	8->21	9->9	N->1	
1	 ->71	(->2	)->1	,->13	-->12	.->22	/->16	0->45	1->21	2->38	3->24	4->21	5->25	6->17	7->15	8->17	9->286	:->1	
2	 ->62	(->2	)->4	,->27	-->4	.->21	/->13	0->172	1->13	2->13	3->6	4->12	5->22	6->9	7->10	8->14	9->8	
3	 ->50	(->3	,->10	-->5	.->9	/->11	0->16	1->8	2->7	3->15	4->11	5->16	6->3	7->12	8->7	9->4	:->1	;->1	?->2	
4	 ->55	(->2	,->8	-->7	.->12	/->12	0->26	1->8	2->5	3->4	4->7	5->13	6->3	7->1	8->8	
5	 ->82	(->3	)->1	,->10	-->63	.->13	/->20	0->20	1->2	2->7	3->1	4->1	5->10	6->2	7->4	8->4	9->4	b->3	
6	 ->66	(->2	)->1	,->13	.->16	/->12	0->6	1->1	2->6	4->1	5->1	6->3	7->12	8->2	9->4	
7	 ->70	(->1	)->2	,->18	.->18	/->20	0->10	1->6	2->1	3->2	4->1	5->4	6->4	7->3	8->8	9->6	?->1	N->1	
8	 ->66	(->2	)->5	,->10	-->3	.->6	/->20	0->31	1->20	2->14	3->2	5->6	6->7	7->5	8->6	9->3	:->2	
9	 ->98	"->1	(->2	)->45	,->12	-->2	.->19	/->19	0->10	1->8	2->7	3->13	4->20	5->22	6->32	7->46	8->47	9->409	:->1	
:	 ->251	A->19	D->2	F->2	a->1	e->3	s->75	
;	 ->101	
?	 ->9	"->1	,->2	-->3	.->13	A->8	B->1	D->35	E->9	F->19	H->32	I->10	J->27	K->13	M->4	N->14	O->6	P->4	R->2	S->8	T->4	U->1	V->36	Ä->13	
A	 ->9	)->2	,->3	-->2	.->3	5->36	:->1	B->4	D->1	F->20	K->1	N->1	R->1	S->2	T->1	c->2	d->5	f->4	g->2	h->8	i->1	k->4	l->88	m->48	n->54	p->6	r->15	s->5	t->35	u->3	v->51	z->2	
B	 ->3	-->2	5->4	A->1	B->3	C->1	I->1	N->16	P->1	R->1	S->6	a->47	e->103	i->13	l->10	o->19	r->47	u->5	y->4	ä->1	å->5	
C	 ->1	,->1	-->1	.->3	4->6	5->22	A->1	E->18	H->4	K->1	L->1	M->1	N->9	O->15	S->3	a->19	e->15	h->2	l->2	o->21	r->2	u->4	y->1	
D	 ->3	)->13	,->1	-->2	A->2	D->4	E->13	R->5	S->1	a->51	e->1610	i->15	o->7	u->12	ä->132	å->25	í->1	ü->1	
E	 ->7	)->5	-->28	/->2	B->1	C->4	D->3	E->3	G->71	I->2	K->13	L->7	M->7	N->47	O->3	P->2	R->4	S->5	U->147	c->1	d->1	f->55	g->2	h->2	i->1	k->5	l->8	m->9	n->117	q->10	r->38	t->51	u->851	v->8	x->8	
F	 ->7	)->2	,->8	.->4	:->2	A->1	B->1	E->3	I->3	J->3	M->1	N->11	O->1	P->19	R->19	S->1	U->1	a->11	e->4	i->21	l->26	o->14	r->195	u->1	y->1	ä->1	å->3	ö->319	
G	 ->7	(->1	,->9	-->58	.->2	:->3	?->1	A->2	F->3	L->2	O->1	U->3	a->17	e->48	i->5	o->19	r->40	u->6	ä->1	å->1	ö->3	
H	 ->1	-->21	O->3	a->83	e->363	i->17	o->9	u->69	y->1	ä->40	å->1	ö->1	
I	 ->282	)->3	,->2	-->3	.->2	:->2	C->4	F->4	I->19	K->3	L->1	M->3	N->9	P->1	R->1	S->1	T->3	V->3	X->2	b->3	d->1	h->1	l->2	m->4	n->84	r->22	s->42	t->18	z->1	
J	)->2	:->1	a->976	e->3	o->25	u->13	ä->3	ö->14	ø->2	
K	 ->2	(->4	,->2	.->2	A->1	O->10	S->8	T->1	a->49	e->1	f->1	i->39	n->1	o->241	r->3	u->27	v->7	y->7	ä->11	ö->3	
L	 ->1	)->8	,->1	-->2	A->20	D->3	F->1	L->1	T->1	a->53	e->20	i->40	l->1	o->19	u->7	y->6	ä->3	å->63	ö->1	
M	 ->2	(->10	-->1	.->1	A->1	I->4	O->3	R->2	U->6	a->102	c->6	e->293	i->67	o->47	u->1	y->5	ä->6	å->13	ö->2	ü->1	
N	 ->4	)->38	,->3	-->2	.->1	:->12	A->3	D->1	G->4	I->10	L->4	M->3	P->9	S->9	T->4	a->35	e->18	i->54	o->9	u->29	y->5	ä->109	å->6	ö->1	
O	 ->4	)->1	,->1	.->2	:->1	?->1	C->1	D->13	F->1	K->1	L->21	M->13	P->1	R->1	S->3	a->2	b->3	c->70	f->5	i->2	l->6	m->120	n->2	r->18	s->4	u->1	z->3	
P	 ->16	)->2	,->3	A->1	E->15	M->1	O->2	P->15	R->1	S->4	T->16	V->3	a->109	e->10	l->11	o->41	r->60	u->3	Ö->21	å->49	é->1	
Q	u->1	
R	 ->2	)->19	-->2	.->1	:->1	A->1	E->5	I->3	N->2	P->1	R->3	a->25	e->42	h->1	i->12	o->23	u->3	y->4	Å->2	Ö->2	ä->3	å->22	é->2	ö->1	
S	 ->2	)->13	-->3	:->1	A->10	D->1	E->17	G->8	K->1	O->1	P->5	R->1	S->3	T->2	U->3	Y->1	a->65	c->38	e->34	h->16	i->6	j->9	k->21	l->39	m->2	n->2	o->69	p->9	r->3	t->55	u->5	v->9	w->3	y->35	á->1	ã->2	ä->5	å->44	ö->2	
T	 ->1	)->19	C->1	E->4	N->2	O->1	T->1	U->1	V->5	a->85	e->7	h->26	i->73	o->18	r->27	s->3	u->38	v->6	y->39	ä->2	å->1	
U	 ->39	,->7	-->48	.->11	:->49	?->1	C->2	E->4	F->1	G->3	N->4	S->12	l->1	n->48	p->7	r->8	t->27	z->2	
V	 ->5	-->4	C->3	D->1	I->5	P->6	a->124	e->21	i->641	l->1	o->3	ä->10	å->31	
W	T->1	a->20	e->2	i->11	o->19	u->5	y->4	
X	 ->2	,->1	V->2	X->2	
Y	N->1	a->1	o->1	t->3	
Z	e->2	i->1	
[	K->2	S->1	
]	.->3	
a	 ->18237	!->18	"->13	)->2	,->721	-->4	.->838	/->3	:->32	;->12	?->39	H->1	N->2	a->16	b->310	c->379	d->2325	e->61	f->317	g->4686	h->45	i->94	j->51	k->978	l->4627	m->3443	n->11481	o->4	p->1104	r->11094	s->2546	t->10412	u->65	v->3516	w->2	x->29	y->26	z->23	ç->5	
b	 ->11	)->2	,->4	-->1	.->2	a->1037	b->161	e->3459	i->612	j->46	l->758	n->1	o->462	p->1	r->487	s->76	t->43	u->228	v->14	y->214	ä->361	å->81	é->2	ö->372	
c	 ->10	"->1	)->1	,->1	-->3	.->5	?->1	C->1	N->5	a->34	c->94	e->616	h->4776	i->656	k->2447	l->1	o->25	q->4	r->1	t->4	u->2	y->12	è->1	
d	 ->3786	!->2	)->4	,->166	-->4	.->219	:->4	;->5	?->10	a->2773	b->268	d->329	e->17773	f->267	g->306	h->32	i->1511	j->242	k->124	l->1013	m->41	n->446	o->458	p->122	r->1692	s->641	t->147	u->261	v->324	w->1	y->24	z->9	ä->526	å->236	é->35	ö->146	
e	 ->10240	!->14	"->5	(->1	)->3	,->370	-->48	.->429	:->46	;->6	?->18	E->1	F->1	H->1	N->2	P->1	a->155	b->391	c->522	d->4065	e->98	f->993	g->1634	h->462	i->753	j->41	k->1655	l->3875	m->2148	n->19085	o->25	p->294	r->16837	s->2865	t->15007	u->435	v->326	w->4	x->415	y->7	z->9	ä->2	å->1	
f	 ->32	,->5	-->4	.->6	a->1351	b->1	d->1	e->659	f->499	h->1	i->832	j->24	k->1	l->304	m->1	o->1057	p->2	r->2791	s->7	t->1089	u->277	y->99	ä->217	å->480	é->1	ö->8318	
g	 ->5596	!->3	"->8	)->7	,->416	-->1	.->470	:->11	;->8	?->16	N->1	a->4624	b->20	d->131	e->4772	f->47	g->612	h->859	i->1054	j->136	k->5	l->361	m->15	n->438	o->1061	p->6	r->1502	s->1452	t->1580	u->30	v->8	y->21	ä->770	å->665	ö->626	
h	 ->4636	!->1	)->1	,->16	-->8	.->5	/->1	:->1	?->1	I->2	a->2986	e->2589	h->1	i->201	j->136	l->4	n->13	o->391	r->26	s->1	t->13	u->326	w->3	y->28	ä->709	å->527	ô->1	ö->463	ü->4	
i	 ->6519	!->5	"->1	,->84	-->14	.->52	:->1	;->1	?->2	a->481	b->150	c->263	d->1688	e->715	f->482	g->5442	h->149	i->8	j->3	k->2354	l->5018	m->235	n->11095	o->3478	p->321	q->4	r->456	s->5758	t->2610	u->28	v->1435	w->1	x->8	z->12	ä->18	å->2	è->1	é->1	ö->24	
j	 ->24	,->13	-->1	.->8	a->1860	d->73	e->466	f->1	i->5	k->4	l->309	n->19	o->359	s->10	t->9	u->460	ä->619	ö->219	
k	 ->926	!->2	"->3	,->101	-->9	.->96	:->2	?->4	a->6520	b->23	d->11	e->2516	f->24	g->35	h->84	i->467	j->31	k->10	l->1191	m->9	n->771	o->4749	p->14	r->1222	s->891	t->3424	u->1517	v->302	y->183	ä->543	å->15	ö->75	
l	 ->4461	!->7	"->5	'->1	,->183	-->38	.->251	:->12	;->3	?->7	F->1	a->5823	b->160	d->577	e->4199	f->240	g->78	h->89	i->5662	j->834	k->666	l->9660	m->585	n->289	o->406	p->170	r->124	s->1228	t->1555	u->852	v->491	y->335	z->6	ä->1212	å->391	é->1	ö->274	ø->2	
m	 ->7285	!->4	"->1	)->2	,->164	-->2	.->192	/->1	:->7	;->2	?->5	I->1	a->2999	b->197	d->37	e->6524	f->460	g->76	h->188	i->3056	j->65	k->31	l->272	m->3339	n->400	o->957	p->622	r->418	s->753	t->438	u->127	v->30	y->619	á->1	ä->566	å->1311	é->8	ö->473	
n	 ->16123	!->251	"->18	)->14	,->1122	-->12	.->1187	/->4	:->36	;->23	?->53	F->3	H->2	I->1	J->2	N->7	a->6371	b->156	c->275	d->7798	e->3704	f->565	g->5811	h->407	i->4004	j->108	k->1507	l->436	m->63	n->2608	o->1455	p->52	r->257	s->5532	t->4890	u->429	v->395	y->481	z->26	Ä->1	ä->951	å->636	ç->1	è->3	ö->201	
o	 ->204	!->1	,->45	-->9	.->49	/->1	:->1	;->1	?->2	N->1	U->2	a->105	b->326	c->5696	d->635	e->195	f->318	g->625	h->9	i->18	j->87	k->395	l->1947	m->10157	n->5704	o->10	p->1505	r->4484	s->814	t->1359	u->65	v->295	w->13	x->19	y->4	ä->17	å->1	ö->7	
p	 ->491	"->4	,->53	-->1	.->58	:->1	?->1	a->2005	b->26	d->28	e->2459	f->131	g->99	h->41	i->69	j->1	k->19	l->490	m->148	n->233	o->1081	p->1784	r->1545	s->199	t->213	u->393	v->11	y->3	ä->14	å->2025	é->11	ö->4	
q	a->2	u->26	
r	 ->22023	!->142	"->11	)->12	,->980	-->20	.->963	:->45	;->14	?->38	H->1	J->1	M->1	N->2	a->9136	b->898	c->9	d->1824	e->6544	f->650	g->616	h->566	i->4242	j->224	k->1394	l->1379	m->745	n->2650	o->3419	p->85	q->1	r->1309	s->2786	t->2217	u->1304	v->469	w->1	y->245	z->1	ä->2046	å->2355	é->2	ê->1	í->1	ó->5	ö->458	
s	 ->6048	!->8	"->3	)->2	,->303	-->58	.->414	/->2	:->7	;->6	?->16	N->1	a->2938	b->192	c->90	d->71	e->2976	f->534	g->57	h->100	i->3207	j->266	k->6529	l->1794	m->478	n->368	o->4417	p->1002	q->2	r->258	s->3654	t->8688	u->450	v->765	w->1	y->655	ä->1591	å->1473	í->1	ö->191	
t	 ->23376	!->23	"->11	)->15	,->1019	-->17	.->1192	:->35	;->13	?->45	B->1	J->1	N->1	a->7810	b->177	c->8	d->17	e->9791	f->338	g->394	h->65	i->8132	j->233	k->72	l->674	m->99	n->918	o->1332	p->51	r->2790	s->2680	t->12537	u->1192	v->916	y->663	z->7	ä->1306	å->630	é->59	ê->3	ó->1	ö->680	ü->1	
u	 ->579	"->1	,->18	-->1	.->9	:->1	;->1	?->1	M->1	a->177	b->99	c->61	d->311	e->95	f->20	g->128	h->4	i->11	k->372	l->1115	m->425	n->2436	o->2	p->1314	q->2	r->2631	s->512	t->3192	u->2	v->138	x->13	y->2	
v	 ->3121	"->1	,->49	.->61	:->2	;->1	?->3	a->2962	b->23	d->44	e->3048	f->34	g->97	h->8	i->5079	j->5	k->29	l->50	m->2	n->61	o->158	p->2	r->109	s->617	t->242	u->82	v->46	y->1	ä->1430	å->793	ö->4	
w	 ->3	,->1	-->1	.->1	a->5	e->8	i->6	n->3	o->7	
x	 ->29	!->1	,->5	-->4	.->22	a->62	b->1	c->6	e->137	f->1	h->1	i->76	k->3	l->5	m->1	n->3	o->4	p->62	t->123	u->4	v->1	x->3	
y	 ->74	!->1	,->9	-->1	.->4	D->1	a->188	b->44	c->795	d->388	e->18	f->98	g->308	h->15	i->2	k->78	l->158	m->66	n->457	o->14	p->56	r->202	s->529	t->339	u->2	v->43	w->1	x->1	å->1	
z	 ->33	)->2	,->9	-->3	.->1	F->1	a->7	b->3	e->2	i->31	j->5	m->2	o->10	q->1	u->1	w->1	á->1	
º	 ->1	
Ä	m->1	n->27	r->33	v->46	
Å	 ->16	D->1	G->1	r->7	t->10	
Î	l->1	
Ö	 ->13	)->2	-->2	:->4	S->2	V->6	g->2	k->1	p->1	s->88	v->3	
á	l->1	n->2	
ã	o->2	
ä	 ->2	c->220	d->271	e->1	f->149	g->977	k->494	l->1775	m->1057	n->3419	p->29	r->5986	s->251	t->1720	v->515	x->58	
å	 ->3919	,->59	.->66	:->7	;->1	?->4	b->15	d->1075	e->166	f->11	g->1507	h->9	j->1	k->97	l->855	m->30	n->1577	o->1	p->51	r->1492	s->901	t->1074	v->89	z->1	
ç	a->5	o->1	
è	r->1	t->1	v->3	
é	 ->26	,->1	a->1	b->2	c->1	e->22	f->3	k->1	n->58	r->2	s->3	t->1	u->2	
ê	t->4	
í	 ->1	e->1	n->1	
ó	n->6	
ô	n->1	
ö	 ->9	!->1	,->12	-->2	.->7	a->10	b->7	c->3	d->655	e->5	f->29	g->169	i->1	j->388	k->314	l->210	m->168	n->168	o->5	p->154	r->9982	s->509	t->228	u->1	v->923	w->1	y->1	ö->1	
ø	n->2	r->2	
ü	h->1	n->1	r->1	s->4	
