 "Am	s->1	
 "At	t->1	
 "Bi	g->1	
 "De	t->4	
 "EU	-->1	
 "Eq	u->1	
 "Eu	r->2	
 "Ja	,->1	
 "Ku	l->4	
 "Kv	i->3	
 "Lo	t->1	
 "Mi	n->1	s->1	
 "Ol	j->1	
 "Om	 ->1	
 "Po	r->1	
 "Ti	b->2	
 "Ty	 ->1	
 "Ur	b->1	
 "af	f->1	
 "al	d->2	l->1	
 "an	g->3	
 "av	g->1	
 "ba	n->1	
 "co	u->1	
 "de	n->3	t->1	
 "dö	d->1	
 "eg	e->1	
 "ek	o->1	
 "en	 ->3	t->1	
 "eu	r->3	
 "fo	r->1	
 "fö	r->1	
 "ge	m->1	n->1	
 "he	l->1	r->1	
 "in	 ->1	l->1	
 "ir	r->1	
 "ja	 ->1	
 "ko	l->2	
 "kr	o->1	
 "ku	l->1	
 "lä	n->1	s->2	
 "me	l->1	
 "na	t->1	
 "ne	 ->1	
 "no	r->1	
 "nå	g->1	
 "ob	e->1	
 "or	m->1	
 "ov	i->1	
 "pa	r->1	
 "på	p->1	
 "re	f->1	s->4	
 "ri	k->1	
 "se	 ->1	
 "sh	a->1	
 "sk	a->1	
 "sp	e->1	
 "sv	a->1	
 "ti	l->1	
 "ut	v->1	å->1	
 "va	l->1	r->1	
 "åt	e->1	
 "öp	p->1	
 "öv	e->1	
 'Va	d->1	
 ("d	i->1	
 (14	0->2	
 (19	9->2	
 (57	1->1	
 (80	9->2	
 (96	1->1	
 (A5	-->35	
 (B5	-->4	
 (Be	n->1	
 (Br	y->2	
 (C5	-->7	
 (CE	N->2	R->1	
 (CO	D->1	
 (DE	)->1	
 (EG	,->1	
 (EI	F->1	
 (EL	)->1	
 (EN	)->23	
 (EU	-->1	G->2	
 (FI	)->1	P->1	
 (FP	Ö->1	
 (FR	)->12	
 (FU	F->1	
 (H-	0->21	
 (Ho	w->1	
 (IC	E->1	
 (IF	O->1	
 (IM	O->1	
 (In	t->1	
 (KO	M->8	
 (Ku	l->2	
 (PP	E->1	
 (PT	)->15	
 (SE	K->1	
 (SP	Ö->1	
 (Ut	s->2	
 (ar	t->7	
 (at	t->1	
 (av	s->1	
 (de	 ->1	t->1	
 (ef	t->1	
 (el	l->1	
 (en	 ->2	
 (fi	s->4	
 (fo	r->1	
 (fö	r->3	
 (hä	l->1	
 (i 	d->1	s->1	
 (in	f->1	r->1	
 (ko	d->2	m->1	n->1	
 (kr	i->2	
 (ma	i->2	
 (me	r->1	
 (oc	h->1	
 (re	c->1	
 (rå	d->1	
 (se	 ->1	
 (så	s->1	
 (t.	e->1	
 (ty	v->1	
 (un	g->1	
 (ÖV	P->1	
 (Ös	t->4	
 (åt	e->1	
 , a	t->1	
 , b	o->1	
 , d	e->1	
 , m	e->1	
 , v	i->1	
 - "	d->1	
 - '	V->1	
 - ,	 ->1	
 - 1	9->26	
 - 2	,->1	
 - 3	1->1	
 - 6	 ->1	
 - 8	0->1	
 - A	l->2	
 - C	4->6	5->14	a->1	
 - D	o->1	
 - E	U->1	
 - H	e->1	
 - K	a->1	o->1	
 - P	a->1	
 - R	e->1	i->1	å->1	
 - S	a->2	
 - a	l->5	n->2	r->1	t->27	v->9	
 - b	e->1	i->1	l->1	ö->1	
 - c	e->1	
 - d	e->51	o->1	v->2	ä->2	å->2	
 - e	f->2	k->1	l->5	n->12	t->3	v->1	x->2	
 - f	a->1	i->1	r->3	å->3	ö->15	
 - g	e->2	ä->1	ö->2	
 - h	a->10	o->1	u->3	ä->1	
 - i	 ->11	d->1	n->16	
 - j	a->15	u->1	
 - k	a->1	n->1	o->9	r->1	
 - l	i->2	y->1	å->2	
 - m	a->3	e->14	i->2	o->2	å->2	
 - n	a->1	y->1	ä->6	å->6	
 - o	c->62	f->1	m->9	r->1	
 - p	a->1	r->2	å->5	
 - r	a->1	e->2	i->1	å->1	ö->1	
 - s	a->5	e->3	i->1	k->3	n->2	o->25	t->3	y->2	ä->2	å->6	ö->1	
 - t	a->1	e->1	i->3	r->3	v->1	ä->1	
 - u	n->1	t->10	
 - v	a->2	e->2	i->18	ä->1	
 - Ö	s->2	
 - ä	r->7	v->10	
 - å	t->2	
 - ö	p->1	v->4	
 -(E	N->1	
 -, 	a->1	d->1	f->1	i->2	m->1	s->1	u->1	ä->1	
 -er	 ->1	
 -or	g->3	
 0 p	r->1	
 000	 ->24	.->1	
 008	 ->2	
 011	3->1	
 055	0->1	
 065	2->1	
 1 0	0->2	
 1 4	0->1	
 1 f	r->1	
 1 i	 ->1	
 1 j	a->5	u->1	
 1 m	a->2	e->1	
 1 o	c->7	
 1 p	r->4	
 1 s	e->1	
 1 u	r->1	t->1	
 1, 	2->1	4->1	a->1	o->1	s->1	
 1,2	 ->2	
 1,4	 ->1	
 1-2	 ->1	
 1-o	m->4	
 1-r	e->5	
 1-s	t->2	
 1.J	a->1	
 1/3	 ->1	
 10 	0->2	e->1	j->1	k->1	m->2	p->4	r->1	s->1	ä->2	å->1	
 10,	 ->1	
 10.	K->1	
 100	 ->9	
 105	 ->2	
 11 	i->1	j->2	m->1	o->1	s->1	
 11,	 ->3	3->1	
 11.	0->3	A->1	E->1	K->1	
 110	 ->1	
 115	 ->1	
 12 	f->1	i->1	j->1	m->2	o->1	p->1	s->1	
 12,	 ->4	
 12.	0->6	
 12/	9->3	
 120	 ->1	
 123	 ->1	
 124	4->3	
 125	 ->1	
 126	0->1	
 13 	(->1	0->1	A->1	f->1	i->2	j->1	n->1	o->1	p->2	s->1	ä->1	
 13,	 ->2	
 13.	0->1	F->1	
 130	 ->1	
 133	.->1	
 138	.->1	
 14 	f->5	m->5	o->1	s->1	t->1	
 14,	 ->1	
 140	 ->1	
 143	 ->1	
 15 	a->1	m->1	o->3	p->3	r->1	s->2	å->1	
 15,	 ->2	
 15.	0->2	
 150	 ->2	
 158	 ->2	)->1	.->1	
 16 	0->1	o->3	p->2	r->1	
 16)	 ->1	
 16,	 ->1	
 164	 ->1	
 166	 ->1	
 167	 ->3	
 17 	d->2	m->1	o->1	s->1	
 17,	 ->2	
 17.	3->1	S->1	
 170	 ->1	
 174	 ->1	
 176	2->2	
 18 	d->1	h->1	i->1	m->2	n->3	
 18,	 ->1	
 180	 ->1	
 19 	d->1	m->1	p->1	s->1	ä->1	
 19.	5->1	
 191	7->1	
 192	3->1	
 193	 ->1	0->1	
 194	.->1	5->1	8->1	
 195	 ->1	7->2	
 196	7->6	9->1	
 197	6->1	7->1	
 198	2->2	6->3	9->1	
 199	0->2	1->3	2->4	3->8	4->6	5->7	6->18	7->40	8->25	9->79	
 2 -	 ->1	
 2 0	0->1	
 2 4	0->1	
 2 b	l->2	
 2 d	e->1	
 2 e	l->1	
 2 i	 ->4	
 2 m	i->1	
 2 o	c->3	
 2 p	r->2	u->1	
 2 s	o->1	
 2, 	1->1	i->1	s->2	v->1	
 2,4	8->1	
 2,6	 ->1	
 2,8	 ->1	
 2-o	m->2	
 2-s	t->1	
 2.1	 ->1	
 2.2	 ->1	
 2.D	e->1	
 2.M	e->1	
 20 	0->1	e->1	g->1	m->2	n->1	p->3	º->1	ä->1	å->5	
 20,	 ->1	
 20.	2->1	
 200	 ->5	0->70	1->2	2->9	3->1	4->1	6->8	7->1	
 201	0->1	2->1	
 21 	j->2	o->2	s->1	ä->1	å->1	
 21.	0->1	5->1	
 21:	a->1	
 22 	a->1	r->1	
 22,	 ->3	5->1	
 22.	Ä->1	
 226	 ->1	
 23 	d->1	i->1	
 23,	7->1	
 24 	n->2	o->2	p->1	
 245	 ->1	
 248	,->1	
 25 	g->1	m->2	o->1	p->7	t->1	
 25.	D->1	
 250	 ->1	
 255	 ->4	
 26 	"->1	i->1	m->1	n->1	o->1	p->1	
 262	 ->1	
 27 	d->1	f->1	l->1	o->1	p->2	
 27,	 ->1	
 28 	f->1	j->1	n->1	p->1	
 28,	 ->2	
 280	 ->4	.->1	
 28:	e->1	
 29 	d->1	f->1	l->1	m->1	
 29,	 ->1	
 299	.->2	
 3 0	0->2	
 3 f	e->1	
 3 j	a->1	
 3 m	a->1	
 3 o	c->1	k->1	
 3 p	r->1	u->1	
 3, 	7->1	
 3,8	 ->2	
 3-4	 ->1	
 3-l	i->2	
 3.1	)->1	
 3.8	 ->1	
 3.I	 ->1	
 30 	f->1	i->2	j->1	m->2	o->1	p->3	
 30,	 ->1	
 300	 ->1	
 31 	f->1	j->1	m->2	o->2	
 314	 ->1	
 32 	m->1	
 32,	 ->2	
 32.	J->1	
 33 	0->2	a->1	f->2	i->1	o->1	
 332	,->1	
 34 	i->1	s->1	t->1	å->1	
 34,	 ->1	
 34.	1->1	
 344	 ->1	
 35 	f->1	m->5	
 35.	S->1	
 350	 ->1	
 36 	f->1	
 36,	 ->1	
 367	 ->1	
 37 	f->1	i->1	p->1	
 37,	 ->2	
 37.	2->1	
 37/	6->1	
 370	 ->1	
 38 	f->2	o->2	
 38,	 ->1	
 38:	 ->1	
 39 	f->1	i->1	p->1	
 39,	 ->1	
 3: 	f->1	
 4 0	0->1	
 4 c	 ->1	
 4 e	n->1	
 4 i	 ->5	
 4 j	u->2	
 4 l	i->1	
 4 o	c->1	
 4 p	r->1	
 4, 	1->2	6->1	o->1	
 4.2	)->1	
 4.I	 ->2	
 4.J	a->1	
 40 	f->1	m->1	p->6	å->3	
 40,	 ->1	
 400	 ->6	
 41 	f->1	p->1	r->1	u->1	
 410	 ->1	
 42 	f->1	i->1	o->2	
 43 	h->1	
 43.	F->1	
 44 	f->1	o->2	
 45 	a->1	c->1	f->1	g->1	
 45,	 ->1	
 45.	 ->1	"->1	H->1	V->1	
 46 	o->2	
 462	 ->1	
 47 	g->1	
 48 	g->1	i->3	ä->1	
 5 0	0->5	
 5 f	r->1	
 5 g	ä->1	
 5 m	i->3	
 5 o	k->1	
 5 v	i->1	
 5 å	r->1	
 5, 	d->1	o->1	u->1	
 5,5	 ->1	
 5,8	 ->1	
 5.4	 ->1	
 5.E	m->1	
 50 	0->1	i->1	m->2	p->3	
 50,	 ->1	
 50-	 ->1	t->2	
 500	 ->1	
 519	 ->1	
 52 	i->1	
 520	 ->2	
 522	 ->1	
 53 	p->1	
 540	 ->1	
 55 	m->1	p->1	
 56 	p->1	
 56,	 ->1	
 57,	5->1	
 5b 	k->1	
 5b-	o->1	
 5b.	D->1	
 6 d	e->1	
 6 f	r->1	
 6 i	 ->6	
 6 m	i->1	
 6 o	c->6	m->1	
 6, 	7->1	t->1	
 6,0	7->1	
 6.S	å->1	
 60 	0->1	f->1	
 60-	t->1	
 600	 ->1	
 62 	i->1	
 67 	i->1	
 68 	a->1	
 685	/->1	
 7 -	 ->1	
 7 d	e->1	
 7 f	ö->1	
 7 g	r->1	
 7 i	 ->8	
 7 l	e->1	
 7 n	ä->1	
 7 o	c->2	
 7 p	r->1	å->1	
 7).	.->1	
 7, 	9->1	d->1	o->2	s->1	
 7,2	 ->1	
 7,4	2->1	
 7.F	r->1	
 70 	a->1	p->1	
 700	 ->4	
 73,	9->1	
 75 	-->1	m->2	
 76 	p->1	
 77 	m->1	
 79/	4->1	
 8 4	6->1	
 8 b	e->1	
 8 f	r->1	
 8 o	c->3	
 8 r	e->1	
 8 t	i->1	
 8 ä	r->1	
 8, 	9->1	s->1	
 80 	e->1	p->11	ä->1	å->1	
 81 	o->5	p->1	
 81.	1->5	3->5	
 82 	h->1	i->1	
 82)	 ->1	
 82,	 ->4	
 82.	I->1	
 83 	p->1	
 85 	o->2	p->1	t->1	
 86 	i->2	p->1	
 87,	 ->1	
 87.	1->1	2->1	
 88 	i->1	o->1	ä->1	
 88/	5->2	
 89 	i->1	t->1	
 9 d	e->1	
 9 f	a->1	e->1	r->1	
 9 i	n->1	
 9 m	i->3	
 9, 	a->1	f->1	
 9.1	 ->1	
 90 	d->2	p->3	
 90-	t->1	
 91 	p->1	
 92/	4->1	
 93 	p->1	
 93/	7->1	
 94 	n->1	p->2	
 94,	 ->1	
 94/	5->2	7->1	
 95 	i->1	m->2	t->1	
 95/	3->1	
 96/	3->3	7->2	
 97.	S->1	
 97/	9->1	
 98 	m->1	
 : P	a->1	
 A. 	G->1	
 ABB	 ->1	-->2	
 ABC	 ->1	
 ADR	)->1	
 AKT	U->1	
 Act	.->1	
 Ada	n->1	
 Ade	n->1	
 Ado	l->2	
 Adr	i->1	
 Afr	i->4	
 Agr	i->1	
 Agu	s->1	
 Ahe	r->7	
 Aid	s->1	
 Akk	u->2	ö->1	
 Ala	v->2	
 Alb	a->2	e->1	r->1	
 Ale	x->2	
 Alg	e->1	
 Ali	c->1	
 All	a->4	t->1	
 Alp	e->1	
 Als	a->3	t->1	
 Alt	e->16	
 Ame	r->1	
 Amo	c->1	k->5	s->1	
 Ams	t->36	
 Ang	e->1	
 Ank	a->1	
 Anl	ä->1	
 Anm	ä->1	
 Ann	a->1	
 Ant	ó->1	
 Anv	e->1	
 Apa	r->1	
 Ara	b->1	f->1	
 Arb	e->1	
 Ari	 ->1	a->3	
 Art	i->1	
 Asi	e->2	
 Ass	a->2	
 Ast	u->1	
 Ata	t->2	
 Atl	a->3	
 Att	 ->3	
 Aus	c->1	
 Aut	o->1	
 Auv	e->1	
 Av 	d->1	o->1	
 Avf	a->1	
 Avi	a->1	
 Avs	e->1	
 Azo	r->2	
 B o	c->1	
 B t	a->1	
 BNI	 ->6	,->1	
 BNP	 ->7	,->2	
 BP,	 ->1	
 BRÅ	D->1	
 BSE	 ->2	-->4	
 Bal	f->1	k->7	
 Ban	k->1	
 Bar	a->9	c->2	e->1	n->15	ó->2	
 Bas	k->2	s->1	
 Bel	g->9	
 Ber	e->12	g->13	l->7	n->5	t->2	
 Bes	l->1	q->1	
 Bet	r->1	
 Bis	c->6	
 Bla	k->1	n->1	
 Blo	k->1	
 Boe	t->1	
 Bol	k->1	
 Bon	d->1	
 Bor	d->1	t->1	
 Bou	r->6	
 Bow	e->2	i->2	
 Bra	n->2	s->1	v->1	
 Bre	m->1	t->7	
 Bri	t->1	
 Bro	k->9	
 Bru	n->1	
 Bry	s->16	
 Bud	a->1	
 Bul	g->1	
 Bus	h->1	q->1	
 Byr	n->2	å->1	
 C. 	D->1	E->1	
 C4-	0->6	
 C5-	0->15	
 CEC	A->1	
 CEN	 ->4	,->2	:->4	
 CSU	-->1	:->1	
 Cad	i->5	o->1	
 Cam	r->1	u->1	
 Can	a->1	d->1	y->3	
 Cas	a->2	
 Cau	d->1	
 Cav	a->1	
 Cen	t->11	
 Cer	m->1	
 Cey	h->1	
 Cha	m->1	
 Chi	q->1	
 Cli	n->1	
 Coc	a->1	i->1	
 Col	a->1	
 Con	a->1	s->1	
 Cor	b->1	
 Cos	t->9	
 Cou	n->1	
 Cox	 ->2	!->1	,->1	
 Cre	s->2	
 Cur	i->1	
 Cus	í->1	
 Cux	h->1	
 Cyp	e->1	
 D k	r->1	
 DDR	.->1	
 Da 	C->3	
 Dag	e->1	m->1	
 Dal	a->6	
 Dam	 ->2	a->1	
 Dan	m->25	
 Dar	m->1	
 Dav	i->3	
 De 	G->1	P->1	R->1	d->2	g->6	h->1	k->1	n->1	o->1	s->3	t->1	
 Del	o->3	
 Dem	i->1	o->1	
 Den	 ->20	n->8	
 Der	a->1	
 Des	s->4	
 Det	 ->75	t->13	
 Deu	t->1	
 Dim	i->5	
 Dir	e->2	
 Dom	s->1	
 Dor	i->1	
 Dub	l->7	
 Duh	a->1	
 Dui	s->3	
 Dut	r->1	
 Där	 ->4	e->1	f->2	
 Då 	b->1	t->1	
 Díe	z->1	
 Düh	r->1	
 E-k	o->1	
 ECH	O->3	
 EDD	,->1	-->2	
 EEG	 ->1	,->2	
 EG 	t->1	
 EG-	d->21	f->8	k->16	r->3	
 EG.	V->1	
 EG:	s->3	
 EIF	 ->1	
 EKS	G->5	
 ELD	R->3	
 EMU	,->1	-->2	:->3	
 EU 	"->1	I->1	a->3	b->2	d->1	f->1	g->2	h->2	i->4	k->3	m->2	o->4	p->1	r->1	s->6	u->2	ä->1	
 EU,	 ->5	
 EU-	b->2	e->1	f->5	g->1	i->5	k->3	l->5	m->6	n->1	p->2	r->2	s->3	t->1	u->1	v->1	
 EU.	.->1	A->1	D->3	F->1	N->1	R->1	V->3	
 EU:	s->44	
 EU?	H->1	
 EUG	F->1	
 Ece	m->1	
 Edi	n->1	
 Eft	a->2	e->9	
 Egy	p->2	
 Ehu	d->2	
 Eie	c->1	
 Eko	f->2	n->1	
 Eli	s->1	
 Ell	e->3	
 Elm	a->2	
 Els	t->1	
 Emi	l->1	
 En 	a->1	b->1	d->1	p->2	v->1	
 End	a->1	
 Enl	i->5	
 Equ	a->7	q->2	
 Era	 ->1	
 Eri	k->24	t->1	
 Erk	k->2	
 Ert	 ->1	
 Eti	o->3	
 Ett	 ->2	
 Eur	a->4	o->790	
 Eva	n->7	
 Exx	o->3	
 FBI	 ->1	
 FEO	 ->2	
 FMI	 ->1	
 FN,	 ->1	
 FN-	u->1	
 FN.	H->1	
 FN:	s->8	
 FPÖ	 ->10	-->2	:->2	
 FRÅ	G->1	
 Fac	t->1	
 Far	o->1	
 Fei	r->2	
 Fin	l->6	n->1	
 Fir	m->1	
 Fis	c->4	
 Fla	u->2	
 Flo	r->16	
 Flé	c->1	
 FoU	,->1	-->1	
 Fog	 ->1	
 Fol	k->3	
 Fon	t->1	
 For	d->1	e->1	
 Fra	g->1	m->1	n->45	s->1	
 Fri	h->2	
 Fru	 ->9	t->2	
 Frä	m->2	
 Frå	g->2	
 Fun	d->1	
 Fäs	t->1	
 Får	 ->2	
 Föl	j->1	
 För	 ->12	b->3	e->40	h->1	i->2	s->12	
 GA-	s->1	
 GAS	P->1	
 GUE	/->2	
 GUS	P->1	
 Gal	e->1	i->2	
 Gam	a->3	
 Gar	g->5	
 Gaz	a->6	
 Gem	e->2	
 Gen	e->9	o->1	è->3	
 Gil	-->2	
 Gin	o->1	
 Goe	b->1	
 Gol	a->8	f->3	l->1	
 Gom	e->1	
 Gon	z->1	
 Goo	d->1	
 Gor	s->1	
 Got	t->1	
 Gra	c->4	ç->5	
 Gre	k->12	
 Gro	s->3	
 Gru	p->8	
 Grö	n->2	
 Gua	t->1	
 Gui	g->1	
 Gul	f->1	
 Gus	p->1	
 Gut	e->2	
 Göt	e->1	
 Haa	r->1	
 Had	e->1	
 Hag	u->1	
 Hai	d->36	
 Ham	b->1	
 Han	 ->1	d->1	s->1	
 Har	 ->4	
 Hat	z->2	
 Hav	e->1	
 Heb	r->1	
 Hed	g->1	k->1	
 Hei	n->1	
 Hel	i->1	s->20	
 Hen	r->1	
 Her	r->30	
 Hic	k->1	
 Hil	t->1	
 Him	a->1	
 Hit	l->6	t->1	
 Hol	l->1	z->2	
 Hon	 ->1	
 Huh	n->1	
 Hul	t->24	
 Hur	 ->1	
 Hän	s->2	
 Här	 ->3	
 Hål	l->1	
 I -	 ->1	
 I S	c->1	
 I T	u->1	
 I b	e->1	u->1	ö->2	
 I d	a->5	e->6	
 I e	g->3	n->1	
 I g	å->1	
 I l	i->1	
 I m	o->2	
 I o	c->2	
 I r	e->1	
 I s	i->1	l->1	t->1	
 I u	t->1	
 I-p	r->1	
 ICE	S->3	
 II 	-->1	h->1	i->1	
 II,	 ->1	
 II-	p->2	
 III	 ->2	
 IMO	.->1	:->1	
 INT	E->4	
 IRA	 ->1	
 ISP	A->1	
 IV 	-->1	i->2	
 IX 	o->1	
 IX,	 ->1	
 Ile	-->1	
 Imb	e->3	
 Ind	i->5	
 Ing	a->1	e->3	l->2	
 Ini	t->1	
 Int	e->22	
 Irl	a->21	
 Isa	b->2	
 Isl	a->1	
 Isr	a->36	
 Ist	a->1	
 Ita	l->17	
 Izq	u->1	
 Ja,	 ->2	
 Jac	k->1	o->2	q->2	
 Jag	 ->140	
 Jan	-->1	
 Jap	a->3	
 Jav	e->1	
 Jea	n->1	
 Jer	u->2	
 Jon	a->2	c->13	
 Jor	d->3	
 Jos	p->1	
 Jug	o->1	
 Jun	k->1	
 Jäm	f->1	
 Jör	g->14	
 Kal	e->3	
 Kan	 ->1	a->1	t->3	
 Kar	a->3	l->6	t->2	
 Kas	p->1	
 Kau	f->1	k->3	
 Kaz	a->1	
 Kfo	r->1	
 Kin	a->10	n->21	
 Kir	g->5	
 Koc	h->14	
 Kom	m->12	
 Kon	k->1	v->1	
 Kor	e->2	
 Kos	o->59	t->1	
 Kou	c->12	
 Kul	t->11	
 Kum	a->1	
 Kun	g->1	
 Kvi	n->1	
 Kvä	k->1	
 Kyo	t->7	
 Kän	n->1	
 Kär	a->1	n->2	
 Köl	n->2	
 Köp	e->1	
 LTC	M->1	
 La 	R->1	
 Laa	n->7	
 Lam	a->7	
 Lan	d->1	g->29	k->3	
 Lap	p->2	
 Lea	d->5	
 Led	a->1	
 Lei	n->8	
 Leo	n->1	
 Lib	a->5	e->2	y->1	
 Lii	k->3	
 Lik	s->2	
 Lil	l->1	
 Lis	s->8	
 Lit	a->1	
 Llo	y->1	
 Loi	r->2	
 Lom	é->2	
 Lon	d->4	
 Lor	d->2	r->2	
 Lot	h->2	
 Lou	s->1	
 Loy	o->2	
 Lut	t->1	
 Lux	e->6	
 Lyn	n->3	
 Låt	 ->12	
 Löö	w->1	
 MAR	P->1	
 Maa	s->6	
 Mac	a->1	
 Mad	a->1	e->2	r->3	
 Mai	n->1	
 Mal	t->5	
 Man	 ->3	
 Mar	g->1	i->8	k->1	p->1	s->1	t->1	
 McC	a->1	
 McN	a->5	
 Med	 ->2	e->3	
 Mel	l->17	
 Men	 ->14	,->1	
 Mex	i->1	
 Mic	h->1	
 Mid	d->1	l->1	
 Min	 ->4	a->1	i->1	u->1	
 Mis	t->1	
 Mit	r->1	t->3	
 Mon	t->19	
 Mor	a->4	b->1	g->4	
 Mos	k->1	
 Mou	r->8	s->1	
 Mul	d->1	
 Mün	c->1	
 Nan	a->1	
 Nap	o->1	
 Nar	k->1	
 Nat	i->4	o->5	
 Ned	e->9	
 Nej	,->1	
 New	 ->1	
 Ni 	b->1	h->3	s->1	v->1	
 Nie	l->5	
 Nik	i->2	
 Nog	u->1	
 Noi	r->1	
 Nor	d->1	g->2	
 Nu 	f->1	
 Nya	 ->2	
 Nyt	t->1	
 När	 ->13	
 Näs	t->1	
 Någ	o->1	
 OCH	 ->1	
 OFS	R->1	
 OLA	F->15	
 OLF	A->1	
 OM 	A->1	
 OSS	E->1	
 Obe	r->1	
 Och	 ->4	:->1	
 Off	e->1	i->1	
 Oil	 ->1	
 Oli	v->1	
 Olj	e->1	
 Oly	m->1	
 Om 	E->1	i->1	m->1	n->1	o->1	
 Oma	g->1	
 One	s->1	
 Ora	n->1	
 Osl	o->3	
 Osm	a->1	
 Ouv	r->1	
 Oz 	d->1	
 Oz,	 ->1	
 PPE	 ->2	-->10	
 PR-	e->1	
 PSE	)->1	-->3	
 PVC	,->1	-->1	.->1	
 Pac	k->3	
 Pad	d->2	
 Pak	i->5	
 Pal	a->15	e->11	
 Pap	a->2	
 Par	i->3	l->4	
 Pat	t->23	
 Pay	s->2	
 Pea	k->1	
 Pei	j->2	
 Pek	i->1	
 Pet	e->1	r->1	
 Pla	n->1	t->1	
 Plo	o->1	
 Poe	t->5	
 Poh	j->1	
 Pol	e->1	l->1	
 Pom	é->1	
 Pon	n->1	
 Poo	s->1	
 Por	t->24	
 Pow	e->3	
 Pre	u->1	
 Pri	o->1	
 Pro	c->1	d->25	v->3	
 Prí	n->1	
 Pur	v->1	
 På 	d->2	g->1	s->1	
 Pås	t->1	
 Pét	a->1	
 Que	c->1	
 REP	 ->2	
 RIN	A->2	
 Rac	k->2	
 Raf	a->3	
 Ran	d->4	
 Rap	k->11	
 Ras	c->1	
 Rea	d->1	
 Red	i->8	
 Reg	e->1	
 Rep	u->1	
 Rev	i->2	
 Rhô	n->1	
 Ric	h->3	
 Rii	s->2	
 Rik	t->1	
 Rio	f->1	
 Rob	e->1	
 Roi	s->1	
 Roj	o->1	
 Rom	-->1	a->2	á->1	
 Roo	 ->1	
 Rot	h->5	t->2	
 Rov	e->2	
 Roy	a->1	
 Rui	z->1	
 Rus	h->1	
 Rys	s->4	
 Råd	e->5	s->1	
 Réu	n->2	
 SEK	 ->1	(->2	
 SEM	-->1	
 SOL	A->1	
 SPÖ	 ->1	
 SS 	o->1	
 Sag	e->1	
 Sai	n->1	
 Sal	a->1	
 Sam	m->15	
 San	 ->1	t->3	
 Sav	e->7	
 Sch	e->10	r->17	u->2	w->2	ö->1	ü->3	
 Sea	t->4	
 Seb	a->1	
 Sed	a->4	
 Seg	n->1	u->1	
 Sei	x->5	
 Sha	r->5	
 She	l->2	p->3	
 Sim	p->1	
 Sju	k->1	
 Sjä	t->1	
 Sjö	s->4	
 Sko	g->1	t->4	
 Sku	l->1	
 Skä	l->1	
 Slo	v->1	
 Soa	r->1	
 Soc	i->1	
 Sok	r->1	
 Sol	a->4	b->2	
 Som	 ->9	
 Sou	l->1	
 Spa	n->7	
 Spe	n->1	r->1	
 Sri	 ->3	
 St.	V->1	
 Sta	d->1	t->1	
 Sto	c->3	r->14	
 Str	a->6	
 Stö	d->1	
 Sua	n->1	
 Sud	r->2	
 Sve	r->7	
 Swo	b->3	
 Syd	a->2	k->1	o->2	
 Syr	i->22	
 Sán	c->1	
 São	 ->2	
 Så 	l->1	r->1	
 Söd	e->2	
 TV 	a->1	
 TV-	k->1	p->1	s->1	
 Tac	i->2	k->7	
 Tad	z->4	
 Tai	w->1	
 Tal	m->1	
 Tam	m->22	
 Tan	g->1	i->1	
 Tau	e->1	
 Ter	r->3	
 Tes	a->1	
 Tex	a->2	
 The	a->19	
 Thy	s->4	
 Tib	e->19	
 Tid	n->1	
 Til	l->8	
 Tod	i->1	
 Tom	 ->1	é->2	
 Tor	r->3	
 Tot	a->6	
 Tra	n->1	
 Tre	d->1	
 Tri	t->1	
 Tro	t->1	
 Tsa	t->3	
 Tur	k->37	
 Tys	k->20	
 Tåg	k->1	
 UCK	 ->1	
 UCL	A->1	
 UEN	-->1	
 UNI	F->1	
 UNM	I->3	
 USA	 ->5	,->2	.->2	:->1	
 USD	 ->1	
 Uls	t->1	
 Und	e->6	
 Uni	o->3	
 Upp	d->1	
 Urb	a->1	
 Urq	u->1	
 Urs	ä->1	
 Utn	ä->1	
 Uts	k->2	
 Utv	ä->1	
 Uzb	e->2	
 V -	 ->1	
 VD 	b->1	
 VI 	i->1	
 VII	I->2	
 Vad	 ->9	
 Val	d->3	l->3	
 Van	 ->2	d->1	
 Vap	e->1	
 Var	e->1	f->1	j->2	k->1	
 Vat	a->3	
 Vel	z->1	
 Vem	 ->3	
 Ven	d->1	e->1	s->2	
 Ver	h->2	s->1	
 Vi 	b->1	f->6	h->10	k->4	m->3	s->4	u->1	v->7	ä->3	
 Vi,	 ->1	
 Vic	h->1	
 Vid	 ->2	
 Vil	k->1	
 Vis	s->1	
 Vit	o->7	
 Viv	i->1	
 Vla	a->1	
 Vod	a->1	
 Vol	k->1	
 Vär	l->3	
 Väs	t->4	
 Vår	 ->2	a->1	t->2	
 WTO	?->1	
 Waf	f->2	
 Wal	e->11	l->4	
 Was	h->3	
 Web	,->1	
 Wes	t->1	
 Wid	e->1	
 Wie	b->1	l->4	n->4	
 Wil	h->1	
 Wog	a->18	
 Wul	f->2	
 Wur	t->3	
 Wye	 ->1	-->2	
 Wyn	n->1	
 X o	c->1	
 XXV	I->2	
 Yas	s->1	
 Yor	k->1	
 Zee	l->2	
 Zim	e->1	
 [KO	M->2	
 [SE	K->1	
 a p	r->3	
 a) 	a->1	b->1	
 abs	o->41	t->1	u->3	
 acc	e->57	
 acq	u->1	
 ad 	h->2	i->1	
 add	i->1	
 ade	k->5	
 adj	e->2	
 adm	i->23	
 adr	i->1	
 adv	o->5	
 aff	ä->4	
 age	n->1	r->42	
 agg	r->1	
 agi	t->1	
 agr	a->1	o->1	
 aid	s->5	
 ajo	u->1	
 akt	 ->7	a->4	e->1	i->27	u->31	ö->10	
 aku	t->1	
 al-	S->1	
 alb	a->9	
 ald	r->29	
 ali	b->1	
 alk	e->1	o->2	
 all	 ->36	a->362	d->22	e->12	i->9	m->121	o->1	r->9	s->18	t->364	v->74	
 alt	a->1	e->11	
 amb	a->1	i->26	u->1	
 ame	r->11	
 an 	a->3	d->2	f->2	p->1	t->1	å->1	
 ana	 ->4	l->43	m->4	
 anb	l->1	u->4	
 and	 ->1	a->12	e->12	l->1	r->314	
 anf	ö->16	
 ang	a->1	e->31	i->2	r->14	å->28	
 anh	ä->4	
 ani	n->5	
 ank	l->3	n->1	o->1	
 anl	e->48	i->1	ä->5	ö->4	
 anm	ä->28	
 ann	a->127	o->4	
 ano	n->4	r->8	
 anp	a->12	
 ans	a->5	e->204	i->1	j->17	k->2	l->46	p->6	t->75	v->276	å->12	ö->10	
 ant	a->135	e->4	i->29	o->23	y->2	
 anv	i->1	ä->158	
 app	a->1	e->1	l->6	
 apr	i->3	o->1	
 ara	b->8	
 arb	e->407	
 arg	u->16	
 ark	i->2	
 arm	o->1	é->3	
 arr	a->6	e->2	o->2	
 art	 ->1	.->2	e->2	i->101	o->1	
 arv	.->2	e->2	
 as"	.->1	
 asp	e->30	
 ass	i->2	o->1	
 ast	r->1	
 asy	l->21	
 atl	a->1	
 ato	m->4	
 att	 ->6121	,->8	.->1	:->1	a->1	e->4	i->5	r->1	
 auc	t->1	
 auk	t->6	
 aut	o->9	
 av 	"->3	-->5	1->4	2->1	5->2	A->5	B->20	C->1	D->7	E->91	F->12	G->6	H->3	I->2	J->4	K->13	L->5	M->4	O->5	P->4	R->2	S->7	T->8	U->1	V->3	W->3	a->177	b->84	c->9	d->587	e->209	f->217	g->50	h->33	i->39	j->11	k->147	l->53	m->103	n->35	o->63	p->79	r->71	s->200	t->73	u->64	v->95	y->5	Ö->2	ä->8	å->23	ö->14	
 av,	 ->5	
 av.	D->3	E->1	J->1	M->1	O->1	
 ava	n->2	
 avb	r->11	
 avd	e->8	
 ave	c->1	u->1	
 avf	a->22	o->1	ö->3	
 avg	a->2	e->10	i->6	j->4	r->3	å->5	ö->55	
 avh	j->2	ä->2	å->1	
 avi	s->4	
 avk	l->1	r->1	u->1	
 avl	a->2	e->2	i->1	o->1	ä->10	
 avm	a->1	
 avp	r->1	
 avr	a->1	e->2	u->1	ä->1	
 avs	a->7	e->83	i->37	k->29	l->74	n->3	p->5	t->32	ä->5	
 avt	a->55	v->1	
 avu	n->1	
 avv	a->6	e->9	i->22	ä->3	
 axe	l->1	
 axl	a->1	
 b) 	i->1	m->1	
 bac	i->1	k->1	
 bad	 ->4	a->1	
 bag	a->2	
 bai	n->1	
 bak	 ->1	d->1	g->31	o->21	å->3	
 bal	a->25	
 ban	a->5	b->1	d->4	k->5	n->1	o->2	t->2	
 bar	 ->1	a->228	b->2	k->1	n->12	r->2	t->1	
 bas	 ->2	,->1	a->2	e->10	i->3	k->5	t->1	
 bax	a->1	
 be 	P->1	e->5	f->1	h->2	k->6	o->2	p->1	s->1	
 bea	k->30	r->2	
 beb	y->1	å->1	
 bed	r->48	ö->44	
 bef	a->11	i->41	l->1	o->72	r->13	ä->12	
 beg	a->4	r->83	ä->60	å->11	
 beh	a->73	o->65	ä->1	å->12	ö->166	
 bei	v->1	
 bek	a->3	l->42	o->2	r->30	v->15	y->16	ä->34	
 bel	a->6	g->8	o->11	y->4	ä->5	ö->2	
 bem	a->1	y->1	ä->5	ö->10	
 ben	e->1	h->1	s->1	ä->1	å->1	
 beo	r->1	
 ber	 ->38	,->1	e->38	i->8	o->40	y->1	ä->31	ö->45	
 bes	e->2	i->4	k->32	l->198	p->2	t->173	v->29	y->1	ä->2	ö->8	
 bet	a->68	e->8	j->1	o->44	r->96	t->2	u->1	v->3	y->122	ä->248	
 beu	n->3	
 bev	a->26	e->1	i->86	
 bib	e->11	l->2	
 bid	r->109	
 bie	f->2	
 bif	a->3	
 big	o->1	
 bil	 ->10	,->2	-->1	.->3	a->83	b->2	d->31	e->6	i->30	j->1	k->4	l->6	m->1	p->7	s->5	t->15	v->6	ä->1	å->1	
 bin	d->14	
 bio	 ->1	l->4	p->1	s->3	
 bis	t->20	
 bit	 ->1	e->1	t->3	
 bju	d->2	
 bl.	a->27	
 bla	m->1	n->56	
 ble	k->1	v->14	
 bli	 ->121	,->1	.->1	c->2	n->2	r->109	v->27	x->1	
 blo	c->4	m->6	t->3	
 blu	n->4	
 bly	 ->1	,->2	.->1	g->4	
 blå	 ->1	
 bo 	i->1	k->1	
 boe	n->1	
 bog	s->1	
 boj	k->1	
 bok	 ->3	s->2	
 bol	a->5	
 bom	b->9	u->1	
 bon	d->2	
 bor	 ->6	d->71	g->3	t->47	
 bos	a->3	n->2	t->5	ä->4	
 bot	 ->2	a->2	t->9	
 bov	a->1	e->1	
 bra	 ->64	!->1	,->8	.->6	n->8	
 bre	d->13	t->7	v->6	
 bri	e->1	n->3	s->60	t->16	
 bro	 ->1	a->1	d->2	k->2	m->10	r->1	t->42	
 bru	k->7	n->1	t->4	
 bry	r->2	t->12	
 brä	n->12	s->2	
 brå	d->20	k->1	
 brö	d->2	s->1	t->1	
 bud	d->1	g->102	o->1	s->10	
 bur	i->1	
 bus	s->1	
 byg	g->50	
 byr	å->34	
 byt	a->1	e->1	t->1	
 byx	f->1	
 bär	 ->16	a->12	s->2	
 bäs	t->42	
 bät	t->75	
 båd	a->23	e->46	
 båt	a->8	e->1	
 béb	é->1	
 böc	k->3	
 böd	e->1	
 böj	e->1	t->1	
 bör	 ->208	,->1	.->1	d->7	j->104	s->1	
 böt	e->1	
 c i	 ->1	
 c) 	l->1	
 ca 	3->1	
 ca.	 ->1	
 cal	v->1	
 can	c->2	n->1	
 cap	i->10	
 cas	e->1	
 cem	e->2	
 cen	t->55	
 cer	t->5	
 cha	n->12	p->1	r->2	
 che	c->1	f->5	
 cho	c->4	k->1	
 cir	k->9	
 cit	a->1	e->7	
 civ	i->19	
 com	b->1	m->1	p->1	
 con	d->1	t->2	
 cop	y->1	
 cor	p->4	r->1	
 cos	t->5	
 cri	c->1	
 d) 	i->1	
 da 	C->5	F->1	
 dag	 ->151	,->28	.->28	:->1	a->17	e->27	l->6	o->52	s->18	
 dam	 ->1	e->41	m->2	
 dan	s->24	
 dat	a->4	o->3	u->13	
 de 	"->1	1->7	2->5	8->1	9->1	C->2	P->6	a->87	b->63	c->4	d->29	e->104	f->165	g->56	h->60	i->83	j->4	k->96	l->42	m->123	n->102	o->92	p->72	r->59	s->229	t->67	u->35	v->62	y->13	ä->31	å->29	ö->23	
 de,	 ->4	
 dea	d->1	
 deb	a->167	
 dec	e->41	
 def	i->35	
 deg	e->1	r->1	
 del	 ->114	,->4	.->4	a->77	e->50	f->1	g->1	l->1	n->1	r->1	s->17	t->56	u->2	v->11	
 dem	 ->143	,->11	.->32	:->2	?->1	a->5	o->122	
 den	 ->1717	)->1	,->10	.->22	;->2	i->2	n->526	s->4	
 dep	a->5	
 der	 ->8	a->84	
 des	 ->1	a->2	s->485	t->3	
 det	 ->2869	!->2	,->44	.->61	:->2	?->3	a->34	s->5	t->828	
 dia	l->31	
 die	 ->1	k->1	
 dif	f->5	
 dig	 ->2	
 dik	e->1	t->4	
 dil	e->3	
 dim	e->12	
 dio	x->2	
 dip	l->11	
 dir	e->212	
 dis	c->14	k->159	p->4	t->3	
 dit	 ->6	h->1	
 div	e->4	
 dju	n->2	p->28	r->14	
 djä	r->7	v->2	
 doc	k->61	
 dog	 ->1	.->2	m->2	
 dok	u->39	
 dol	l->9	
 dom	 ->2	a->16	e->2	i->7	s->62	
 dra	 ->25	b->45	g->9	m->6	r->10	s->5	
 dri	c->3	f->5	v->20	
 dro	g->6	p->1	
 dru	c->2	n->3	
 dry	f->1	g->3	
 drå	p->1	
 drö	j->7	m->1	
 du 	b->2	c->1	m->1	ä->2	
 dub	b->15	
 dug	a->1	
 duk	t->1	
 dum	h->3	p->4	t->1	
 dun	a->1	
 dus	s->1	
 dvs	.->45	
 dyk	a->2	e->5	
 dyl	i->3	
 dyn	a->5	
 dyr	 ->1	a->4	t->2	
 dys	t->1	
 däc	k->1	
 däm	p->2	
 där	 ->214	!->1	,->10	.->14	?->1	a->2	e->20	f->184	h->1	i->24	m->40	p->2	t->1	v->4	
 då 	2->1	D->1	E->3	a->11	b->11	d->16	e->1	f->9	g->2	h->4	i->12	j->3	k->11	m->9	o->9	p->4	r->4	s->12	t->8	u->1	v->13	ä->2	ö->1	
 då,	 ->2	
 då.	D->1	
 då?	I->1	
 dål	i->19	
 dåv	a->1	
 dö 	i->1	
 död	 ->5	.->3	a->9	f->1	s->2	
 döe	n->1	
 döl	j->10	
 döm	a->9	d->1	t->1	
 döp	a->1	e->2	t->1	
 dör	 ->4	r->7	
 döt	t->3	
 e) 	i->1	
 e-m	a->1	
 e.d	.->1	
 ecu	 ->1	,->1	
 ed 	g->1	
 ede	n->1	
 eff	e->129	
 eft	e->358	
 ege	n->99	t->25	
 egn	a->44	
 ego	i->2	
 ej 	a->3	b->3	i->1	k->1	l->1	n->1	ä->1	
 ej,	 ->1	
 ej.	E->1	R->1	
 eko	l->13	n->243	s->4	
 ekv	a->1	
 el-	 ->2	S->4	
 ele	f->1	k->10	m->9	
 eli	m->3	
 ell	e->323	
 elm	a->1	
 elo	g->2	
 elv	a->2	
 emb	a->1	l->1	r->1	
 eme	d->1	l->63	
 emi	g->2	
 emo	t->55	
 en 	"->6	P->1	R->1	S->1	a->157	b->107	c->18	d->106	e->152	f->170	g->146	h->76	i->48	j->9	k->138	l->66	m->195	n->68	o->90	p->87	r->137	s->304	t->81	u->65	v->110	y->3	z->1	ä->13	å->16	ö->55	
 en,	 ->2	
 en.	E->1	
 ena	 ->35	d->5	s->7	t->2	
 enb	a->30	
 end	 ->1	a->120	e->1	
 ene	r->98	
 eng	a->18	e->10	
 enh	e->53	ä->32	
 eni	g->10	
 enk	e->36	l->11	
 enl	i->122	
 eno	r->32	
 ens	 ->14	a->7	e->3	i->4	k->28	t->5	
 ent	r->4	u->3	y->4	
 env	e->1	i->5	
 epo	k->4	
 er 	-->2	a->25	b->4	d->3	e->10	f->7	g->1	h->3	i->4	k->6	l->1	m->2	n->1	o->20	p->4	r->2	s->14	t->9	u->11	v->5	ä->1	å->1	
 er,	 ->25	
 er.	B->1	J->3	K->1	N->1	O->1	P->1	
 er:	 ->2	
 era	 ->37	
 erb	j->19	
 erf	a->26	o->5	
 erh	å->7	ö->3	
 eri	n->13	
 erk	ä->39	
 ers	a->1	ä->21	
 ert	 ->36	,->2	
 erö	v->1	
 et 	o->1	
 eta	b->12	p->4	
 etc	.->5	?->1	
 eti	k->1	s->1	
 etn	i->11	
 ett	 ->1363	,->2	.->2	:->1	
 eur	o->391	
 eve	n->21	
 evi	g->3	
 ex 	a->4	p->1	t->1	
 exa	k->18	m->16	
 exc	e->5	
 exe	m->116	
 exi	l->2	s->17	
 exk	l->3	
 exp	a->6	e->45	l->2	o->5	
 ext	e->7	r->30	
 f.d	.->2	
 fab	r->1	
 fac	k->4	
 fad	d->1	
 fai	l->1	
 fak	t->133	
 fal	l->160	s->3	
 fam	i->15	
 fan	n->15	t->11	
 far	 ->1	a->10	h->2	l->58	m->1	o->4	s->1	t->61	v->9	
 fas	,->1	c->7	o->1	t->111	
 fat	t->79	
 fau	n->1	
 fav	o->1	
 fax	a->1	
 feb	r->16	
 fed	e->8	
 fel	 ->10	!->1	,->3	.->4	a->13	b->1	k->1	r->1	s->1	
 fem	 ->25	,->1	:->1	p->1	t->24	å->3	
 fen	o->3	
 fic	k->26	
 fie	n->3	
 fil	m->1	o->5	
 fin	 ->1	a->77	l->5	n->381	s->6	
 fir	a->1	
 fis	k->40	
 fjo	l->3	r->9	
 fjä	r->11	
 fla	g->13	m->4	
 fle	r->98	s->25	x->27	
 fli	c->1	t->2	
 flo	d->4	r->1	t->2	
 fly	g->13	k->14	r->1	t->10	
 flä	k->1	
 flö	d->1	
 fod	e->6	
 fog	 ->1	a->1	
 fok	u->5	
 fol	k->77	
 fon	d->26	
 for	a->1	c->1	d->68	m->70	s->36	t->192	u->3	ê->1	
 fos	s->2	
 fot	b->1	f->1	s->2	
 fra	k->1	m->654	n->36	s->1	
 fre	d->64	k->1	s->4	
 fri	 ->12	,->1	-->8	a->24	g->6	h->66	k->1	s->5	t->3	v->12	
 fro	d->4	n->2	
 fru	 ->67	,->1	k->16	s->2	
 fry	s->2	
 frä	c->1	m->139	
 frå	g->675	n->578	
 ful	l->96	t->1	
 fun	d->13	g->54	k->27	n->9	
 fus	i->7	k->1	
 fut	t->1	
 fyl	l->7	
 fyr	a->25	t->3	
 fys	i->9	
 fäd	e->1	
 fäl	l->4	t->6	
 fän	g->1	
 fär	d->5	g->1	r->2	s->1	
 fäs	t->12	
 få 	1->1	E->1	G->1	a->5	b->8	d->16	e->41	f->13	g->2	h->2	i->7	k->6	l->7	m->9	n->3	o->6	p->9	r->5	s->25	t->22	u->3	v->11	ä->1	å->1	ö->1	
 få,	 ->3	
 få.	E->1	G->1	V->1	
 fåg	e->3	l->6	
 fån	g->5	
 får	 ->182	,->2	?->1	k->1	
 fås	 ->1	
 fåt	a->1	t->57	
 föd	d->1	e->4	o->1	s->1	
 fög	a->2	
 föl	j->121	l->4	
 fön	s->1	
 för	 ->3090	,->16	.->13	;->1	?->2	a->35	b->204	d->185	e->733	f->104	g->6	h->164	i->4	k->76	l->92	m->54	n->74	o->69	p->26	r->59	s->960	t->98	u->76	v->150	ä->67	å->3	ö->8	
 föt	t->3	
 gag	n->7	
 gal	e->1	l->1	n->1	
 gam	l->28	m->4	
 gan	s->26	
 gar	a->90	d->1	
 gas	k->1	
 gat	o->1	
 gav	 ->9	,->1	s->2	
 ge 	F->1	a->8	b->6	d->13	e->27	f->3	g->2	h->4	i->3	j->1	k->4	m->4	n->2	o->10	p->6	r->9	s->7	t->3	u->12	v->3	
 ge.	J->1	
 ged	i->2	
 gem	e->379	
 gen	a->11	d->6	e->38	g->1	o->378	s->1	t->27	u->1	
 geo	g->8	s->2	
 ger	 ->63	,->1	
 ges	 ->14	t->2	
 get	t->21	
 gic	k->8	
 gif	t->2	
 gig	a->5	
 gil	l->1	t->15	
 gis	s->1	
 giv	a->17	e->27	i->4	
 gjo	r->112	
 gla	d->24	s->2	
 gle	s->1	
 glo	b->12	
 glu	p->1	
 glä	d->40	
 glö	m->19	
 gnu	t->2	
 gnä	l->1	
 god	 ->23	.->1	a->37	k->88	o->3	s->38	t->46	
 gol	v->1	
 got	t->19	
 gra	d->23	n->63	t->40	v->5	
 gre	k->7	p->2	
 gri	p->8	
 gro	g->1	u->1	v->1	
 gru	n->255	p->138	v->1	
 gry	m->1	
 grä	l->2	m->1	n->57	
 grå	 ->1	z->1	
 grö	d->1	n->17	v->1	
 gud	s->2	
 gul	d->1	t->1	
 gum	m->1	
 guv	e->1	
 gyn	n->11	
 gäc	k->1	
 gäl	l->404	
 gär	n->33	
 gå 	a->2	b->2	e->1	f->7	g->2	h->1	i->20	l->5	m->3	o->3	p->1	s->4	t->10	u->5	v->4	å->1	
 gå.	O->1	V->1	
 gån	g->132	
 går	 ->83	,->4	.->2	d->3	
 gåt	t->20	
 göm	m->3	t->1	
 gör	 ->131	,->1	.->3	a->284	s->15	
 ha 	a->5	b->5	d->10	e->55	f->6	g->5	h->7	i->3	k->10	l->4	m->12	n->10	o->2	p->2	r->3	s->14	t->11	u->5	v->14	y->1	ä->2	å->1	ö->3	
 ha,	 ->1	
 ha.	A->1	
 had	e->85	
 haf	t->37	
 hak	a->1	
 hal	t->1	v->24	
 ham	b->1	m->1	n->38	
 han	 ->117	,->2	d->258	k->1	s->76	t->34	
 hap	p->1	
 har	 ->1670	,->14	.->2	:->1	?->1	m->18	
 has	t->1	
 hat	 ->1	e->1	i->1	t->1	
 hav	 ->2	,->1	e->23	s->18	
 heb	r->1	
 hed	e->3	r->3	
 hej	d->2	
 hek	t->2	
 hel	 ->11	a->105	g->1	h->29	i->1	l->52	s->47	t->143	
 hem	 ->5	.->2	b->1	f->1	l->15	m->10	s->3	v->1	
 hen	n->27	
 her	r->209	
 hes	 ->1	
 het	a->1	e->2	s->2	t->3	
 hie	r->4	
 hig	h->1	
 hin	d->43	n->2	
 his	t->33	
 hit	 ->4	,->1	t->58	
 hjä	l->99	r->18	
 hob	b->2	
 hoc	-->2	
 hom	o->4	
 hon	 ->29	o->28	
 hop	p->100	
 hor	d->2	i->3	m->1	
 hos	 ->49	p->1	
 hot	 ->11	a->18	b->1	e->8	f->1	
 hug	g->3	
 hum	a->6	l->1	ö->2	
 hun	d->11	
 hur	 ->196	.->2	u->14	
 hus	 ->3	,->2	.->1	ö->1	
 huv	u->47	
 hyc	k->5	
 hyg	i->2	
 hyl	l->2	
 hyp	o->2	
 hyr	d->1	
 hys	a->3	e->5	t->1	
 häf	t->1	
 häl	e->1	f->3	s->23	
 häm	m->1	n->2	
 hän	d->72	f->1	g->14	s->79	t->7	v->35	
 här	 ->261	,->14	.->9	;->1	?->1	e->1	i->2	j->2	l->1	m->3	r->4	t->1	v->1	
 häs	t->1	
 häv	a->1	d->28	t->1	
 hål	 ->1	,->1	l->147	
 hån	 ->1	a->1	
 hår	d->17	e->1	k->1	t->9	
 håv	a->1	
 hög	 ->21	,->1	a->16	e->18	l->1	n->3	r->20	s->29	t->17	
 höj	a->5	d->8	e->1	n->2	t->1	
 höl	l->6	
 hön	a->1	
 hör	 ->31	.->1	a->22	d->5	n->3	t->17	
 hös	t->1	
 i "	g->1	
 i -	 ->1	
 i 1	5->1	
 i 2	0->3	
 i A	B->1	d->2	f->3	k->2	l->1	m->17	s->1	u->1	v->1	
 i B	N->1	e->11	i->5	o->1	r->11	u->1	
 i C	E->1	a->1	e->6	u->1	
 i D	D->1	a->9	u->4	
 i E	C->1	G->8	K->3	M->1	U->15	k->1	t->1	u->171	
 i F	a->1	e->1	i->2	o->1	r->11	ö->14	
 i G	U->1	a->2	e->2	o->2	r->4	u->2	
 i H	a->1	e->14	
 i I	C->2	n->1	r->10	s->2	t->6	
 i J	o->1	
 i K	a->3	f->1	i->3	o->35	y->1	ä->1	ö->1	
 i L	a->3	e->1	i->6	o->6	u->5	
 i M	a->5	c->1	e->16	i->1	o->3	
 i N	e->5	o->1	
 i O	L->1	m->1	
 i P	P->3	a->3	e->1	o->5	
 i R	a->1	o->1	y->2	
 i S	a->3	c->4	e->3	h->4	k->2	r->3	t->15	v->2	y->4	
 i T	V->1	a->17	e->1	h->5	i->5	u->7	y->5	
 i U	E->1	S->3	r->1	
 i V	a->1	e->1	ä->1	
 i W	a->4	i->1	
 i Y	a->1	
 i a	b->1	i->1	k->4	l->52	n->29	r->36	t->12	v->7	
 i b	a->1	e->36	i->14	r->4	u->9	å->3	ö->6	
 i c	e->2	i->1	
 i d	a->167	e->523	i->19	o->3	r->1	
 i e	f->8	g->12	k->5	n->127	r->14	t->61	u->3	x->2	
 i f	.->1	a->7	e->10	i->1	j->2	l->5	o->31	r->141	u->3	y->2	ä->2	ö->141	
 i g	a->1	e->23	l->1	o->8	r->8	ä->1	å->23	
 i h	a->27	e->23	i->2	j->2	u->7	ä->9	å->1	ö->9	
 i i	c->2	n->10	t->1	
 i j	a->1	o->1	u->11	ä->3	
 i k	a->28	e->1	l->3	n->1	o->45	r->26	u->4	v->4	
 i l	a->16	e->2	i->15	j->5	y->1	ä->1	å->1	
 i m	a->12	e->35	i->45	j->1	o->41	y->2	ä->1	å->21	ö->1	
 i n	a->3	i->4	o->7	u->1	y->2	ä->8	å->10	ö->1	
 i o	c->16	f->4	k->2	l->6	m->18	n->1	r->8	u->1	ö->1	
 i p	a->38	e->4	l->8	o->10	r->40	u->2	
 i r	a->10	e->37	i->5	u->1	ä->11	å->34	
 i s	a->55	e->14	i->104	j->24	k->8	l->19	m->2	n->2	o->4	p->1	t->95	v->1	y->58	ä->4	å->12	ö->1	
 i t	.->1	a->7	e->1	i->21	j->1	o->5	r->10	v->6	ä->2	
 i u	n->35	p->4	r->2	t->41	
 i v	a->27	e->10	i->56	ä->20	å->60	
 i y	r->2	t->2	
 i z	o->2	
 i Ö	V->1	s->37	
 i ä	g->1	k->1	m->2	n->9	r->1	
 i å	r->12	t->5	
 i ö	r->1	s->3	v->17	
 i, 	s->1	u->1	
 i.A	n->1	
 i.D	e->2	
 i.N	ä->1	
 i.S	e->1	å->1	
 iak	t->8	
 ian	s->1	
 ibe	r->1	
 ibl	a->19	
 ick	e->34	
 ida	g->1	
 ide	a->5	e->2	n->18	o->5	
 idr	o->4	
 idé	 ->10	,->1	e->8	n->14	
 ifa	l->2	
 ifr	å->35	
 ige	n->46	
 ign	o->4	
 igå	n->7	
 ihj	ä->1	
 iho	p->10	
 ihä	r->1	
 ihå	g->16	
 ika	p->1	
 ikr	a->4	
 ill	a->6	e->8	o->2	v->1	
 ils	k->2	
 ima	g->2	
 imm	a->1	i->6	u->1	
 imp	l->1	o->9	u->6	
 in 	2->1	F->1	a->1	b->3	d->6	e->1	f->3	h->1	i->26	k->2	l->1	m->2	n->1	o->3	p->24	r->2	s->5	u->3	v->4	y->1	
 in,	 ->4	
 inb	e->12	j->7	l->14	y->1	
 inc	i->8	
 ind	e->2	i->27	u->43	
 ine	f->3	
 inf	e->2	i->3	l->11	o->89	r->15	ö->159	
 ing	a->26	e->113	i->6	r->16	å->33	
 inh	e->2	ä->6	
 ini	f->1	t->68	
 ink	l->21	o->14	r->1	ö->3	
 inl	e->72	ä->23	å->2	ö->1	
 inn	a->39	e->215	o->5	
 ino	m->283	
 inp	r->1	
 inr	e->84	i->46	y->1	ä->54	
 ins	a->42	e->38	i->10	k->11	l->6	p->11	t->221	y->13	
 int	a->12	e->1769	i->1	o->6	r->163	y->4	ä->2	
 inv	a->19	e->24	i->1	o->9	ä->13	å->8	
 inö	v->1	
 ira	k->1	
 irl	ä->8	
 iro	n->2	
 irr	a->2	g->1	i->4	
 is 	j->2	
 isc	e->1	
 iso	l->7	
 isr	a->19	
 ist	ä->1	
 isä	r->2	
 ita	l->17	
 itu	 ->20	
 ive	r->2	
 ivä	g->3	
 ja 	-->1	e->1	i->1	n->1	t->3	
 ja,	 ->5	
 jag	 ->1069	,->15	.->2	a->2	
 jak	t->3	
 jan	u->16	
 jap	a->1	
 jet	t->1	
 job	b->4	
 jon	i->1	
 jor	d->69	
 jou	r->2	
 ju 	E->1	M->1	a->11	b->2	d->5	e->2	f->2	h->1	i->11	l->1	m->5	o->8	p->3	r->2	s->6	t->1	u->1	v->1	ä->6	
 ju,	 ->2	
 jub	l->1	
 jud	a->1	e->1	i->1	
 jul	 ->1	f->1	i->10	k->1	
 jun	g->1	i->12	
 jur	i->45	
 jus	t->104	
 juv	e->1	
 jäm	f->16	k->1	l->8	n->4	s->24	v->2	
 jär	n->17	
 jät	t->1	
 kab	a->1	i->3	
 kad	m->3	
 kal	l->33	
 kam	,->1	m->58	p->28	r->1	
 kan	 ->781	,->3	a->7	d->13	i->1	o->1	s->57	
 kao	s->2	
 kap	a->5	i->20	p->1	t->2	
 kar	a->11	g->1	r->1	t->14	
 kas	k->1	t->3	
 kat	a->65	e->5	o->7	
 ked	j->4	
 kel	t->1	
 kem	i->6	
 kid	n->1	
 kil	o->5	
 kin	e->9	
 kl.	 ->20	1->1	
 kla	g->5	p->1	r->143	s->19	u->4	v->1	
 kli	b->1	e->1	m->12	
 klo	a->1	c->2	k->7	
 kly	f->5	
 km 	l->1	m->1	
 km,	 ->1	
 km.	T->1	
 kna	p->16	
 kni	p->1	
 kno	w->1	
 knu	s->1	t->7	
 kny	t->8	
 knä	c->2	
 koa	l->12	
 kod	 ->2	e->3	
 kof	f->1	
 koh	e->1	
 kok	o->1	
 kol	-->1	d->5	l->202	o->1	
 kom	 ->25	b->1	m->1965	p->85	
 kon	c->37	f->44	g->1	j->1	k->327	s->224	t->180	v->19	
 koo	p->1	
 kop	i->2	p->5	
 kor	,->1	n->1	r->39	t->73	
 kos	t->101	
 kra	f->71	s->1	v->70	
 kre	a->3	t->6	
 kri	g->14	m->7	n->16	s->24	t->62	
 kro	a->1	m->2	p->1	s->1	
 kry	p->3	s->1	
 krä	n->17	v->134	
 krå	n->2	
 krö	n->1	
 kub	i->1	
 kul	a->2	i->1	l->1	o->1	t->107	
 kum	u->2	
 kun	d->30	g->15	n->254	s->15	
 kur	s->8	
 kus	t->27	
 kva	l->42	n->7	r->35	
 kve	s->3	
 kvi	c->3	n->59	
 kvo	t->11	
 kvä	l->9	v->2	
 kyl	a->2	i->1	
 käl	l->9	
 käm	p->5	
 kän	d->7	n->58	s->35	t->8	
 kär	a->53	e->1	l->3	n->53	
 kök	s->1	
 köl	 ->1	,->1	a->1	d->2	
 kön	e->3	s->1	
 köp	 ->1	a->1	e->1	k->1	s->1	t->1	
 kör	 ->1	a->2	n->1	s->2	t->2	
 köt	t->2	
 l'e	a->1	
 la 	L->1	
 lab	o->3	
 lad	e->17	
 lag	 ->4	,->4	.->3	a->13	d->1	e->8	f->5	l->6	o->1	r->1	s->115	t->58	
 lan	d->165	s->4	t->1	
 lap	p->3	
 lar	m->4	v->1	
 las	t->7	
 law	,->1	.->1	
 le 	b->1	p->1	
 led	 ->1	a->167	d->11	e->32	n->15	s->4	
 leg	a->15	i->18	
 lej	d->1	
 lek	e->1	t->1	
 lem	.->1	l->1	
 let	a->1	t->10	
 lev	a->13	d->1	e->15	n->6	t->1	
 lib	a->1	e->25	
 lic	e->1	
 lid	a->1	e->7	i->3	
 lig	a->1	g->75	
 lik	a->59	g->2	h->16	n->20	r->3	s->49	t->2	v->8	
 lil	l->5	
 lin	b->1	d->6	j->12	o->1	
 lis	t->12	
 lit	a->8	e->56	t->8	
 liv	 ->7	,->3	.->3	e->10	s->101	
 lju	d->2	g->1	s->10	
 lob	b->5	
 loc	k->2	
 log	i->13	
 loj	a->5	
 lok	a->42	
 lop	p->2	
 los	s->2	
 lot	t->4	
 lov	 ->2	a->11	o->2	v->2	y->1	
 luc	k->5	
 lud	d->2	
 luf	t->2	
 lug	n->6	
 luk	t->1	
 lun	c->1	
 lur	a->2	
 lut	a->1	h->1	
 lyc	k->59	
 lyd	a->2	e->3	
 lyf	t->8	
 lyk	t->1	
 lys	a->6	s->29	
 läc	k->4	
 läg	e->21	g->130	l->1	r->10	s->1	
 läk	a->4	e->1	
 läm	n->56	p->46	
 län	d->114	g->101	k->1	
 lär	 ->1	a->7	d->8	o->2	t->2	
 läs	 ->1	a->3	b->2	e->6	f->1	k->1	t->5	
 lät	 ->5	t->37	
 läx	a->2	
 låg	 ->7	a->5	t->2	
 lån	g->116	
 lås	e->1	t->2	
 låt	 ->14	a->27	e->6	i->1	s->2	
 löf	t->11	
 löj	e->3	
 lök	m->1	
 lön	 ->1	e->2	s->5	t->4	
 löp	a->6	e->7	t->7	
 lör	d->1	
 lös	 ->1	a->34	e->1	g->1	n->48	r->1	t->7	
 löv	s->1	
 m.m	.->1	
 mag	e->1	n->1	
 mai	n->5	
 maj	 ->5	,->1	.->2	o->38	
 mak	r->6	t->39	
 mal	t->3	
 man	 ->621	,->13	.->1	a->2	d->23	i->1	l->1	n->1	t->2	
 mar	g->5	i->3	k->188	s->11	
 mas	k->4	o->1	s->11	t->1	
 mat	c->1	e->26	n->1	p->1	t->2	
 max	b->1	i->7	
 med	 ->1478	,->12	.->6	a->24	b->171	d->57	e->96	f->22	g->20	h->1	i->12	k->5	l->343	v->57	
 meg	a->1	
 mek	a->9	
 mel	l->199	
 men	 ->383	,->4	a->31	i->47	
 mer	 ->173	!->2	,->2	.->7	a->11	g->1	i->1	p->1	v->5	
 mes	t->44	
 met	a->4	o->23	
 mid	d->1	
 mig	 ->210	!->1	,->15	.->5	:->1	?->1	r->2	
 mik	r->4	
 mil	d->4	i->9	j->261	l->7	s->1	
 min	 ->151	,->1	a->72	d->52	i->66	n->20	o->22	s->93	u->21	
 mir	a->1	
 mis	s->76	t->2	ä->2	
 mit	t->70	
 mix	.->1	
 mju	k->1	
 mob	i->7	
 mod	 ->4	e->55	i->6	
 mog	e->2	
 mom	s->1	
 mon	e->7	i->1	o->19	s->1	t->1	
 mor	a->6	d->8	g->36	s->6	
 mot	 ->204	,->1	a->1	g->1	i->21	o->8	p->4	s->73	t->16	v->6	å->3	
 mul	t->9	
 mun	t->8	
 mur	a->1	
 mus	i->4	s->2	
 mut	o->1	
 myc	k->452	
 myg	g->1	
 myl	l->1	
 myn	d->109	n->1	
 myt	i->1	
 mäk	t->3	
 män	 ->9	.->2	g->18	n->94	s->43	
 mär	k->23	
 mät	a->3	t->1	
 må 	h->2	v->1	
 måh	ä->5	
 mål	 ->71	,->12	-->1	.->13	:->1	a->1	e->33	i->4	m->1	s->15	
 mån	 ->10	,->1	a->72	d->4	g->161	
 mår	.->1	
 mås	t->696	
 måt	t->5	
 möb	l->1	
 möd	o->1	r->1	
 möj	l->281	
 mör	d->5	k->2	
 möt	a->6	e->24	t->1	
 nac	k->6	
 nai	v->2	
 nak	n->1	
 nam	n->16	
 nar	k->6	
 nat	i->177	t->3	u->120	
 naz	i->8	
 ned	 ->21	.->2	e->9	g->2	l->4	m->3	r->1	s->7	v->1	
 neg	a->26	
 nej	 ->2	,->2	.->1	
 nek	a->5	
 neo	n->2	
 nep	o->5	
 ner	 ->5	e->3	
 neu	t->2	
 ni 	a->25	b->10	d->7	e->4	f->12	g->5	h->24	i->14	j->3	k->17	l->3	m->3	n->8	o->6	p->3	r->5	s->30	t->7	u->5	v->23	ä->7	ö->1	
 ni,	 ->11	
 ni.	D->1	
 nim	b->1	
 nio	 ->13	n->1	
 niv	å->67	
 nju	t->1	
 nog	 ->14	,->1	.->2	a->12	g->12	
 nol	l->3	
 nom	i->3	
 non	 ->2	
 nor	d->15	m->33	r->5	
 not	a->1	e->28	
 nov	e->11	
 nr 	1->5	2->2	3->10	4->7	5->1	6->1	7->1	8->1	9->1	
 nu 	-->1	3->1	E->1	a->7	b->8	d->7	e->11	f->20	g->14	h->15	i->10	k->11	l->5	m->10	n->9	o->7	p->6	r->4	s->20	t->11	u->4	v->7	ä->16	å->1	
 nu,	 ->6	
 nu.	.->1	J->1	L->1	V->1	
 nu:	 ->1	
 nu?	J->1	
 nul	l->1	ä->1	
 num	e->5	m->2	
 nun	n->1	
 nuv	a->45	
 ny 	b->1	e->1	f->4	g->1	h->1	i->2	k->8	l->3	m->1	o->2	p->2	r->2	s->6	t->1	u->1	v->3	
 nya	 ->163	,->1	;->1	n->3	s->1	
 nyb	i->2	
 nyc	k->7	
 nyd	a->1	
 nye	 ->1	t->1	
 nyf	a->1	ö->1	
 nyh	e->12	
 nyk	t->3	
 nyl	i->30	
 nyn	a->6	
 nyp	l->1	
 nys	k->1	s->13	
 nyt	t->77	
 nyv	a->1	
 nyå	r->1	
 näm	l->43	n->83	
 när	 ->349	,->1	a->20	h->5	i->12	m->36	s->1	v->46	
 näs	d->1	t->47	
 nät	 ->2	.->1	e->1	s->1	t->1	v->11	
 nå 	a->1	d->2	e->7	f->4	h->1	v->1	ä->1	å->1	
 nåb	a->2	
 nåd	 ->1	
 någ	o->357	r->147	
 når	 ->2	
 nåt	t->7	
 nöd	b->1	e->1	i->1	s->1	v->123	
 nöj	a->10	d->9	e->6	t->1	
 nöt	.->1	k->3	s->1	t->1	
 oac	c->31	
 oak	t->1	
 oan	s->5	v->1	
 oav	b->2	s->10	
 oba	l->6	
 obe	b->1	f->1	g->5	h->2	r->50	s->5	
 obj	e->1	
 obl	i->14	
 obs	e->2	
 och	 ->4549	,->9	/->1	
 ock	s->585	u->5	
 odd	s->1	
 ode	l->1	
 odi	s->1	
 odj	u->2	
 odu	g->1	
 oef	t->1	
 oeg	e->5	
 oek	o->1	
 oen	i->4	s->4	
 oer	h->12	s->1	
 oet	i->1	
 of 	t->1	
 ofa	n->2	
 ofe	l->1	
 off	e->89	i->5	r->16	
 ofr	e->1	å->3	
 oft	a->54	
 ofu	l->2	
 ofö	r->21	
 oge	n->2	
 ogr	u->2	
 ogy	n->1	
 ohj	ä->1	
 ohä	m->1	
 ohö	v->1	
 oig	e->1	
 oin	s->2	t->4	
 ojä	m->7	
 okl	a->14	
 oko	n->2	
 okr	i->1	ä->1	
 okt	o->8	
 oku	n->3	
 okä	n->2	
 ola	g->4	
 oli	k->120	
 olj	a->8	e->32	
 olo	g->1	
 oly	c->45	m->1	
 olä	m->3	
 olö	s->2	
 om 	"->3	-->5	1->4	2->1	3->5	4->2	6->1	A->3	B->2	C->1	D->1	E->18	F->2	G->4	H->4	I->3	J->1	K->6	L->3	M->2	P->1	S->2	T->7	a->259	b->44	c->1	d->338	e->131	f->83	g->20	h->67	i->53	j->28	k->82	l->28	m->90	n->40	o->23	p->20	r->61	s->91	t->37	u->44	v->115	y->2	Ö->3	ä->13	å->12	ö->9	
 om"	.->1	
 om)	;->1	
 om,	 ->21	
 om.	 ->1	A->1	D->7	E->2	I->1	J->6	M->3	N->1	O->1	S->2	V->1	
 omI	.->1	
 omb	a->1	e->5	o->1	u->12	
 omd	e->1	i->1	ö->2	
 ome	d->21	
 omf	a->83	l->1	o->3	å->2	ö->1	
 omg	e->1	i->1	å->3	
 omh	u->1	
 omi	s->1	
 omk	r->15	
 oml	a->1	o->2	
 omm	ö->1	
 omo	r->3	
 omp	l->1	r->8	
 omr	i->1	å->222	ö->35	
 oms	o->9	t->47	v->1	ä->8	
 omt	a->1	
 omv	a->5	ä->12	
 omö	j->16	
 ond	 ->1	a->3	o->1	s->1	
 one	-->1	
 ons	d->5	
 ont	 ->1	.->1	
 onö	d->11	
 opa	r->2	
 ope	r->12	
 opi	n->4	
 opp	o->7	
 opr	a->1	o->2	
 opt	i->8	
 ord	 ->40	,->2	.->1	:->2	a->6	e->37	f->193	l->1	n->22	r->3	v->2	
 ore	a->2	d->1	g->1	
 org	a->69	
 ori	e->5	g->2	k->3	m->5	
 ork	a->3	
 orm	 ->1	e->1	
 oro	 ->36	,->4	.->9	a->21	l->6	n->5	s->4	v->2	
 ors	a->29	
 ort	,->1	.->1	
 orw	e->1	
 orä	k->1	t->10	
 osa	n->1	
 oss	 ->288	,->15	.->18	:->1	?->2	
 ost	r->3	
 osv	.->6	
 osy	n->1	
 osä	k->8	
 oså	r->1	
 ota	c->1	
 oti	l->17	
 otj	ä->1	
 otr	o->2	y->1	
 otv	e->2	i->1	
 oty	d->4	
 otä	n->1	
 otå	l->1	
 oum	b->4	
 oun	d->6	
 out	h->2	n->1	
 ova	n->7	
 ove	r->1	
 ovi	l->3	s->1	
 ovä	d->2	l->1	s->1	
 oän	d->4	
 oön	s->1	
 oöv	e->6	
 p.g	.->1	
 pak	e->2	t->1	
 pal	e->12	
 pap	p->5	
 par	 ->16	a->14	c->1	k->3	l->389	t->111	
 pas	 ->1	s->17	
 pat	e->1	i->2	
 pea	n->1	
 ped	a->1	o->1	
 pek	a->19	
 pel	a->8	
 pen	g->55	n->11	s->6	
 per	 ->24	f->7	i->60	m->8	r->1	s->118	
 pes	s->2	t->4	
 pet	i->1	
 pha	r->1	
 pht	a->1	
 pil	o->3	
 pio	n->1	
 pir	a->1	
 pla	c->14	n->81	s->5	t->31	
 ple	n->9	
 pli	k->5	m->1	
 plu	n->1	r->1	s->2	
 plä	d->2	
 plå	n->1	
 plö	t->4	
 poe	t->1	
 pol	e->2	i->339	
 poo	l->1	
 pop	u->5	
 por	s->1	t->74	
 pos	i->80	t->2	
 pot	e->5	
 poä	n->12	
 pra	c->1	g->1	k->32	t->4	x->7	
 pre	c->43	f->3	j->4	l->3	m->10	r->1	s->58	
 pri	c->2	m->1	n->113	o->36	s->22	v->28	
 pro	b->156	c->134	d->62	f->10	g->153	j->54	k->1	n->1	p->11	s->1	t->31	v->15	
 prä	g->4	
 prö	v->7	
 psy	k->1	
 pub	l->7	
 pum	p->2	
 pun	d->3	k->168	
 pur	i->1	
 pyr	a->1	
 på 	-->5	1->4	2->4	3->3	4->1	5->3	7->2	8->3	9->2	A->3	B->7	C->2	E->18	F->1	G->2	H->1	I->9	M->1	O->1	P->1	R->3	T->1	V->2	a->205	b->39	c->3	d->313	e->224	f->96	g->106	h->23	i->26	j->7	k->49	l->34	m->77	n->64	o->38	p->23	r->49	s->126	t->49	u->16	v->90	y->1	z->1	Ö->2	ä->9	å->7	ö->8	
 på,	 ->16	
 på.	B->1	D->4	E->2	J->3	N->1	O->1	U->1	V->1	Ä->2	
 på:	 ->3	
 på?	.->1	J->1	
 påb	j->1	ö->11	
 påd	r->1	
 påf	r->1	ö->3	
 påg	i->3	å->18	
 pål	a->1	i->1	ä->1	
 påm	i->30	
 påp	e->49	
 pås	k->7	t->21	
 påt	a->9	r->3	v->4	
 påv	e->36	i->3	
 qua	 ->2	
 quo	 ->1	,->1	
 rad	 ->20	e->4	i->18	
 rak	 ->1	a->2	r->1	t->3	
 ram	 ->9	,->2	.->2	a->6	e->58	p->11	v->3	
 ran	d->14	n->1	
 rap	p->98	
 ras	a->3	h->1	i->25	
 rat	i->20	
 rea	g->16	k->20	l->14	
 rec	i->1	y->1	
 red	a->166	e->2	l->1	o->17	s->1	u->4	
 ree	l->4	
 ref	e->4	l->7	o->127	
 reg	e->313	i->253	l->89	
 reh	a->1	
 rej	ä->3	
 rek	l->2	o->44	r->1	
 rel	a->23	e->9	i->5	
 rem	i->1	
 ren	 ->4	a->2	g->1	o->3	s->8	t->22	
 rep	a->5	r->16	u->10	
 res	a->7	e->9	i->1	o->98	p->83	t->11	u->147	
 ret	o->3	r->12	
 rev	i->35	o->1	
 rid	a->1	
 rig	h->1	o->4	
 rik	a->11	e->10	l->2	t->156	
 rim	l->18	m->1	
 rin	g->6	
 ris	,->1	:->1	k->84	
 ro 	i->1	
 ro,	 ->2	
 roc	k->1	
 rol	i->1	l->64	
 rom	e->5	
 rop	a->2	e->1	
 ros	 ->2	e->1	t->1	
 rot	a->1	s->1	
 rub	b->3	r->1	
 rui	n->1	
 rul	l->6	
 rum	 ->27	,->1	.->4	
 run	d->4	t->6	
 rus	a->3	t->2	
 rut	i->7	t->2	
 ryc	k->1	
 ryg	g->4	
 ryk	t->8	
 rym	m->1	
 rys	k->2	s->1	
 räc	k->34	
 räd	d->20	s->8	
 räk	e->8	n->48	
 rät	a->1	t->490	
 råd	 ->11	,->1	.->2	?->1	a->10	d->1	e->308	f->6	g->13	s->27	
 råg	a->1	
 råk	a->1	
 råo	l->1	
 råt	t->1	
 réf	é->1	
 röd	a->2	g->1	
 rör	 ->37	a->26	d->1	e->5	i->2	l->24	t->1	
 rös	t->120	
 röt	t->5	
 röv	a->1	
 s.k	.->4	
 sa 	a->1	
 sad	e->75	
 saf	e->1	
 sag	t->49	
 sak	 ->32	,->2	.->3	:->1	e->42	f->1	k->2	l->1	n->35	o->2	p->1	
 sal	i->1	u->1	
 sam	a->80	b->47	e->2	f->13	h->42	l->21	m->275	o->37	r->9	s->7	t->148	v->5	
 san	k->7	n->16	s->2	t->15	
 sat	e->1	s->17	t->14	
 sce	n->6	
 sch	a->1	
 sci	e->1	
 sco	r->1	
 se 	a->12	b->1	d->8	e->4	f->5	h->6	i->5	k->1	m->2	n->1	o->6	p->8	r->2	s->5	t->68	u->5	v->9	ä->1	ö->10	
 sed	a->101	e->1	
 seg	 ->1	d->1	e->4	l->13	r->1	
 sei	s->2	
 sek	e->4	l->2	r->12	t->47	u->3	
 sel	e->1	
 sem	e->4	i->1	
 sen	 ->1	a->97	f->1	s->1	t->6	
 sep	a->1	t->15	
 ser	 ->71	b->14	i->7	v->7	
 ses	 ->10	s->6	
 set	t->49	
 sex	 ->17	,->1	i->1	m->1	t->1	u->2	v->1	
 sid	a->74	o->7	
 sif	f->17	
 sig	 ->366	,->8	.->18	;->1	n->13	
 sik	t->27	
 sim	m->1	u->2	
 sin	 ->156	a->138	e->3	n->5	o->1	s->3	
 sis	t->57	
 sit	t->104	u->116	
 sju	 ->4	,->1	k->12	n->13	t->2	
 sjä	l->173	t->19	
 sjö	f->7	m->2	n->5	s->4	t->1	v->1	
 ska	 ->2	d->56	f->5	k->2	l->672	m->7	n->7	p->175	r->4	t->33	
 ske	 ->17	!->1	,->1	d->4	p->14	r->31	t->15	
 ski	c->16	l->61	n->1	p->2	s->4	
 skj	u->25	
 sko	g->36	l->8	n->1	
 skr	a->2	e->5	i->30	o->29	ä->8	
 sku	g->3	l->498	r->1	t->3	
 sky	d->74	f->1	h->1	l->29	m->1	n->7	
 skä	l->43	m->3	n->2	r->14	
 skå	d->2	
 skö	n->1	r->6	t->17	v->1	
 sla	g->34	k->1	m->1	p->3	v->1	
 sli	p->2	r->1	t->1	
 slo	g->2	t->1	v->1	
 slu	k->3	m->5	s->2	t->172	
 slä	c->3	k->1	p->10	
 slå	 ->10	e->1	r->3	s->1	
 slö	s->4	
 sma	k->1	
 smi	d->3	t->2	
 smu	l->1	s->1	t->3	
 smä	d->1	r->3	
 små	 ->53	,->2	.->1	f->5	g->1	n->4	s->1	
 sna	b->71	r->66	
 sne	d->12	
 snä	l->1	v->1	
 snå	r->1	
 snö	v->1	
 so 	f->1	
 soc	i->203	
 sof	t->1	
 sol	a->1	d->2	i->30	s->1	
 som	 ->3365	,->21	l->3	m->3	
 sop	a->1	
 sor	g->4	t->8	
 sov	j->1	
 spa	n->11	r->9	
 spe	c->84	g->3	k->7	l->52	n->5	t->2	
 spi	l->1	
 spl	i->3	
 spo	n->5	r->1	t->1	
 spr	i->15	å->9	
 spä	n->10	r->3	
 spå	r->8	
 spö	k->4	
 sri	l->1	
 sta	b->23	c->1	d->36	g->2	l->2	n->28	r->75	t->217	
 ste	e->1	g->35	l->3	n->3	r->1	
 sti	c->5	f->1	g->6	l->4	m->11	
 sto	d->5	l->11	p->18	r->298	
 str	a->90	i->39	u->124	y->8	ä->37	å->4	ö->9	
 stu	d->13	g->1	m->1	n->10	
 sty	c->2	m->2	r->34	
 stä	d->12	l->172	m->17	n->20	r->22	v->2	
 stå	 ->25	e->3	l->40	n->117	r->95	t->4	
 stö	d->379	l->1	r->114	t->17	
 sub	j->1	s->27	v->10	
 suc	c->5	
 sud	d->1	
 sum	m->10	
 sun	d->5	
 sup	r->1	
 sus	p->1	
 sut	t->1	
 suv	e->17	
 sva	g->21	n->1	r->74	
 sve	k->2	n->2	p->2	
 svä	l->2	
 svå	g->1	n->1	r->91	
 syd	e->1	k->1	v->1	ö->1	
 syf	t->68	
 sym	b->9	p->9	
 syn	 ->6	a->4	d->8	e->4	l->7	n->51	o->1	p->21	s->5	t->1	v->12	
 syr	i->8	
 sys	s->108	t->114	
 säg	:->1	a->173	e->73	s->5	
 säk	e->224	r->19	
 säl	j->3	l->5	
 säm	r->5	s->5	
 sän	d->14	k->6	
 sär	a->1	b->1	k->1	s->156	
 säs	o->1	
 sät	e->1	t->308	
 så 	a->133	b->13	d->8	e->4	f->18	g->4	h->14	i->7	j->1	k->27	l->31	m->52	n->5	o->6	p->3	r->3	s->93	t->6	u->5	v->28	ä->16	ö->1	
 så,	 ->6	
 så.	 ->1	D->1	I->1	O->1	
 så:	 ->1	
 såd	a->163	
 såg	 ->6	v->1	
 såh	ä->1	
 sål	e->40	u->4	
 sån	g->3	
 sår	b->2	
 sås	o->31	
 såt	i->1	
 såv	i->3	ä->40	
 söd	r->6	
 sök	a->4	e->5	
 sön	d->7	e->1	
 sör	j->10	
 t.e	x->19	
 t.o	.->7	
 ta 	A->1	a->6	b->2	d->21	e->13	f->9	g->1	h->36	i->18	l->4	m->7	n->1	o->5	p->2	r->2	s->18	t->9	u->59	v->3	ö->3	
 ta.	J->1	
 ta?	D->1	
 tab	u->1	
 tac	k->144	
 tag	 ->4	e->14	i->58	n->1	
 tak	 ->1	,->1	e->1	t->7	
 tal	 ->6	,->1	.->3	a->168	e->7	m->418	r->4	s->1	
 tan	k->82	
 tap	p->3	
 tar	 ->64	v->1	
 tas	 ->32	k->1	
 tax	-->3	e->1	
 tea	t->1	
 tec	k->11	
 tek	n->45	
 tel	e->6	
 tem	a->2	p->6	
 ten	d->12	
 teo	r->2	
 ter	a->2	m->3	r->27	
 tex	t->35	
 the	 ->3	
 tib	e->9	
 tid	 ->46	,->7	.->7	e->51	i->85	n->4	p->10	s->36	t->6	
 tig	e->2	g->1	
 til	l->2539	
 tim	m->9	
 tin	g->3	
 tio	 ->10	t->6	
 tis	d->2	
 tit	e->1	t->22	
 tja	t->1	
 tjo	c->2	
 tju	g->4	
 tjä	n->118	r->1	
 tob	a->2	
 tog	 ->21	s->8	
 tol	e->14	k->24	v->1	
 tom	 ->1	m->1	r->2	
 ton	 ->14	,->1	/->2	g->1	v->4	å->1	
 top	p->12	
 tor	d->1	k->1	n->1	p->2	s->8	t->2	v->4	
 tot	a->34	
 tox	i->1	
 tra	d->18	f->7	g->10	k->1	m->1	n->107	s->3	u->1	v->2	
 tre	 ->63	,->2	:->1	d->72	k->1	m->1	n->1	t->5	v->3	
 tri	l->1	o->1	
 tro	 ->11	.->1	d->3	g->1	j->1	l->9	n->1	r->151	t->48	v->14	
 tru	p->2	s->3	
 try	c->6	g->6	
 trä	 ->2	d->23	f->9	n->3	p->1	s->1	t->7	
 trå	d->4	k->3	n->1	
 trö	g->1	s->4	t->1	
 tuf	f->2	
 tul	l->2	
 tum	m->3	
 tun	c->1	g->17	n->4	
 tur	 ->6	,->1	.->1	e->1	i->22	k->8	
 tus	e->9	
 tve	k->29	t->5	
 tvi	n->25	s->6	v->38	
 tvu	n->11	
 tvä	r->17	t->1	
 två	 ->122	.->1	:->2	h->1	n->6	
 ty 	E->1	d->4	i->1	n->2	p->2	v->2	
 tyc	k->77	
 tyd	e->6	l->104	
 tyg	e->1	
 tyn	a->1	g->10	
 typ	 ->20	,->1	.->2	e->16	f->1	g->1	
 tys	k->22	t->3	
 tyv	ä->29	
 täc	k->14	
 täm	l->3	
 tän	d->1	k->73	
 täp	p->4	
 tär	t->1	
 tät	a->2	e->2	
 täv	l->3	
 tåg	 ->1	,->1	e->1	k->1	o->1	
 tål	 ->1	a->2	
 töm	m->1	
 u-l	ä->1	
 ult	i->1	r->2	
 umg	ä->1	
 und	a->52	e->473	g->1	r->11	v->35	
 ung	 ->1	a->6	d->14	e->8	
 uni	k->2	l->2	o->432	v->4	
 upp	 ->196	,->11	.->17	b->13	d->26	e->47	f->126	g->85	h->29	k->6	l->24	m->136	n->93	r->97	s->76	t->22	v->7	
 ur 	E->2	U->1	b->4	d->4	e->12	i->1	j->1	k->2	m->8	p->2	s->3	t->1	v->1	
 ura	n->11	
 urb	a->1	
 urh	o->4	
 urm	i->1	
 urs	k->4	p->20	ä->14	
 urv	a->13	
 ut 	1->1	T->1	a->7	b->1	d->7	e->6	f->8	g->1	h->3	i->4	k->2	m->8	n->2	o->5	p->19	r->2	s->8	t->3	u->2	ö->5	
 ut,	 ->20	
 ut.	 ->1	D->5	F->3	G->1	J->4	K->1	S->1	V->1	Ä->1	
 ut:	 ->1	
 ut?	.->1	E->1	
 uta	n->319	r->41	
 utb	a->1	e->5	i->45	r->4	u->4	y->14	
 utd	e->1	
 ute	 ->4	l->3	s->23	
 utf	a->4	l->2	o->39	r->7	ä->13	ö->37	
 utg	a->1	i->16	j->4	å->29	ö->59	
 uth	ä->2	
 uti	f->16	
 utj	ä->5	
 utk	a->16	o->3	r->3	
 utl	a->5	o->3	ä->7	å->2	ö->2	
 utm	a->20	y->1	ä->32	
 utn	y->40	ä->4	
 uto	m->16	
 utp	e->1	l->2	r->2	
 utr	e->8	i->19	o->5	u->3	y->7	ä->2	
 uts	a->6	e->9	i->1	k->126	l->20	t->42	u->1	ä->7	å->3	
 utt	a->98	j->24	o->2	r->72	ö->5	
 utv	a->1	e->228	i->104	ä->31	
 utö	k->12	v->28	
 vac	k->9	
 vad	 ->238	?->1	
 vag	a->2	n->1	t->1	
 vak	a->2	s->9	t->1	u->2	
 val	 ->12	,->2	.->4	;->1	b->1	d->23	e->7	f->5	k->4	l->1	r->1	t->12	u->22	
 van	 ->32	a->1	h->2	l->11	o->1	s->1	
 vap	e->13	n->2	
 var	 ->217	,->1	.->1	a->368	d->5	e->21	f->39	g->1	i->74	j->83	k->14	m->15	n->12	o->1	s->29	t->8	v->6	
 vat	t->26	
 vec	k->40	
 ved	e->13	
 vek	h->4	
 vel	a->7	
 vem	 ->17	s->1	
 ven	t->1	
 ver	b->1	i->1	k->337	s->11	t->3	
 vet	 ->85	,->11	a->28	e->81	t->4	
 vi 	-->3	1->1	5->1	E->2	L->1	P->1	a->128	b->108	d->56	e->44	f->97	g->52	h->175	i->194	j->11	k->123	l->27	m->90	n->35	o->44	p->15	r->28	s->161	t->62	u->38	v->74	y->1	ä->47	å->7	ö->8	
 vi,	 ->16	
 vi.	V->1	
 vi?	.->1	
 via	 ->12	
 vic	e->13	
 vid	 ->204	,->2	.->2	a->39	d->2	g->2	h->5	m->1	s->1	t->64	
 vif	t->1	
 vig	v->1	ö->1	
 vik	t->352	
 vil	a->2	d->1	j->177	k->317	l->592	s->3	t->1	
 vin	 ->1	d->5	n->6	s->11	
 vir	k->3	r->1	
 vis	 ->11	,->2	.->1	a->123	d->1	e->7	i->2	k->1	s->187	t->5	u->3	
 vit	b->50	t->5	
 vol	u->4	y->3	
 von	 ->18	
 vor	e->29	
 vot	e->3	u->1	
 vra	k->4	
 vre	d->1	
 vri	d->1	
 vrä	k->1	
 vun	n->3	
 vux	i->1	n->2	
 väc	k->17	
 väd	e->1	j->9	
 väg	 ->17	,->9	.->5	N->1	a->12	b->1	e->19	l->5	m->1	n->16	r->20	s->2	
 väk	t->2	
 väl	 ->55	,->2	.->3	b->1	d->20	f->9	g->3	j->22	k->53	l->1	m->4	s->8	t->2	u->3	
 vän	 ->1	d->20	l->4	n->2	s->16	t->45	
 väp	n->2	
 vär	d->70	l->50	n->3	r->2	s->8	t->4	
 väs	e->29	t->2	
 väv	n->3	t->1	
 väx	a->9	e->10	l->3	t->12	
 våg	 ->1	a->6	e->1	l->1	
 vål	d->12	l->1	
 vån	i->2	
 vår	 ->139	,->1	a->150	d->2	t->106	
 vör	d->1	
 wal	e->1	
 web	b->1	
 wor	s->1	
 yng	r->1	s->1	
 ypp	a->1	e->1	
 yrk	a->2	e->18	
 yta	.->1	
 ytl	i->2	
 ytt	e->89	r->42	
 zig	e->4	
 zon	 ->2	e->1	i->1	
 º C	.->1	
 Ämn	a->1	
 Änd	å->1	
 Änn	u->2	
 Är 	k->1	
 Ära	d->2	
 Äve	n->11	
 Å P	S->1	
 Å k	o->1	
 Å s	o->1	
 Årl	i->1	
 Åtg	ä->3	
 Île	-->1	
 ÖVP	 ->4	
 Öpp	e->1	
 Öst	e->80	t->2	
 äck	l->1	
 äga	 ->18	n->3	r->15	
 ägd	e->1	
 äge	r->5	
 ägg	"->1	
 ägn	a->28	
 ägt	 ->9	
 äkt	e->1	
 äld	r->7	
 äls	k->2	
 ämb	e->7	
 ämn	a->4	e->25	
 än 	1->6	2->2	3->2	E->1	F->1	W->1	a->15	b->2	d->20	e->33	f->9	g->1	h->3	i->12	j->1	k->6	l->3	m->12	n->7	o->2	p->4	r->4	s->10	t->7	v->18	ä->4	
 än,	 ->1	
 än.	J->1	
 änd	a->20	l->1	p->1	r->288	å->53	
 äng	s->1	
 änn	u->77	
 änt	l->20	
 är 	"->1	-->4	1->1	2->1	3->1	E->12	F->1	P->2	W->1	a->231	b->110	c->2	d->356	e->360	f->161	g->45	h->51	i->176	j->45	k->68	l->53	m->140	n->105	o->93	p->41	r->49	s->153	t->64	u->49	v->131	y->10	ä->16	å->2	ö->31	
 är,	 ->13	
 är.	.->1	D->2	E->1	F->1	H->1	J->2	k->1	
 är:	 ->5	
 är?	H->1	
 ära	d->22	n->4	
 äre	n->18	
 ärl	i->8	
 äro	 ->1	
 äte	r->1	
 äve	n->275	
 å P	P->1	
 å a	n->7	
 å d	e->3	
 å e	n->11	
 å m	i->2	
 å r	e->1	
 å u	t->1	
 åbe	r->1	
 åhö	r->1	
 åkl	a->37	
 åkt	e->1	
 åla	g->3	
 åld	e->9	
 åli	g->5	
 ålä	g->5	
 åny	o->1	
 år 	-->1	1->19	2->33	a->7	b->1	d->2	e->6	f->8	h->2	i->4	k->3	l->1	n->1	o->7	p->2	s->26	t->3	u->2	v->1	ä->2	å->1	
 år,	 ->18	
 år.	D->9	E->1	F->2	H->2	I->1	J->2	K->1	L->1	O->1	R->1	S->1	T->1	V->3	Ä->1	
 åra	t->1	
 åre	n->39	t->31	
 årh	u->7	
 årl	i->8	
 års	 ->11	b->2	r->2	t->1	
 årt	a->1	i->1	u->3	
 åsa	m->3	t->1	
 åsi	k->50	
 åsk	å->2	
 åst	a->25	
 åsy	f->5	
 åt 	E->1	F->1	a->8	b->1	d->27	e->6	f->2	g->1	h->1	i->3	j->1	k->4	l->1	m->1	n->2	p->1	r->4	s->6	t->3	u->1	Ö->1	ä->3	å->1	
 åt,	 ->2	
 åt.	K->1	N->1	
 åta	 ->3	g->30	l->18	n->1	r->2	
 åte	r->250	
 åtf	ö->12	
 åtg	ä->218	
 åtm	i->27	
 åtn	j->1	
 åts	k->3	t->2	
 ått	a->5	o->1	
 åvi	l->1	
 öar	 ->1	n->5	
 öbo	 ->1	
 öde	 ->1	,->4	.->1	?->1	l->1	m->1	s->4	
 öga	t->1	
 ögo	n->19	
 öka	 ->29	.->3	d->36	n->3	r->16	s->3	t->16	
 ökn	i->18	
 öl 	o->1	
 öm 	t->1	
 ömm	a->1	
 öms	e->5	
 ömt	å->1	
 ön 	N->1	
 öns	k->63	
 öpp	e->78	n->20	
 öre	 ->1	g->7	
 öro	n->3	
 öst	 ->1	b->1	e->52	l->1	r->2	u->2	
 öva	t->1	
 öve	r->602	
 övn	i->5	
 övr	i->65	
! 19	9->1	
! Al	l->2	
! At	t->1	
! Av	 ->1	f->1	s->1	
! Be	r->1	s->1	t->1	
! Bl	a->1	
! Ce	n->1	
! Da	g->1	
! De	 ->3	n->10	t->39	
! Di	r->1	
! Dä	r->1	
! Dí	e->1	
! EU	 ->1	
! Ef	t->4	
! En	d->1	
! Er	a->1	t->1	
! Et	t->1	
! Eu	r->7	
! Fr	a->1	u->1	å->1	
! Få	r->1	
! Fö	r->16	
! Ge	n->1	
! Go	t->1	
! Gr	u->3	
! He	r->1	
! Hi	t->1	
! I 	b->3	d->9	e->3	l->1	m->1	u->1	
! In	g->1	t->1	
! Ja	,->1	g->109	
! Jo	n->1	
! Jä	m->1	
! Ka	r->1	
! Ko	m->4	n->1	
! Li	k->2	
! Lå	t->9	
! Ma	n->1	
! Me	d->1	
! Mi	n->5	
! Ni	 ->5	
! Nu	 ->1	
! Nä	r->7	
! Nå	g->1	
! Ol	j->1	
! Om	 ->2	
! PP	E->1	
! Pa	r->1	
! Pr	i->1	
! På	 ->2	s->1	
! Re	g->1	
! Ro	t->1	
! Rå	d->2	
! Sc	h->1	
! Se	d->3	
! Sk	u->1	
! So	m->7	
! St	r->1	
! Ta	c->3	
! Th	e->1	
! Ti	l->7	
! To	r->1	
! Tr	o->1	
! Un	d->4	
! Up	p->1	
! Ur	s->1	
! Ut	s->2	
! Va	d->4	r->1	
! Vi	 ->20	d->2	s->1	
! Vå	r->3	
! Än	n->1	
! Äv	e->9	
! Å 	P->1	k->1	s->1	
! År	l->1	
! Ös	t->1	
!".D	e->1	
!"De	t->1	
!"Ja	g->1	
!"Om	 ->1	
!(Pa	r->1	
!. (	F->1	
!.(N	L->1	
!.He	r->1	
!All	t->2	
!Ams	t->1	
!And	r->1	
!Av 	d->1	
!De 	a->1	f->1	s->1	
!Den	 ->2	n->1	
!Det	 ->13	t->1	
!Där	f->1	
!Eft	e->2	
!En 	v->1	
!Eri	k->1	
!Eur	o->1	
!Fru	 ->3	
!För	 ->1	e->1	
!Gen	o->1	
!Han	 ->1	
!Her	r->9	
!Här	 ->1	
!I d	e->1	
!Jag	 ->18	
!Kul	t->1	
!Led	a->1	
!Låt	 ->1	
!Med	 ->1	
!Men	 ->4	
!Min	 ->1	a->1	
!Myc	k->1	
!Män	n->1	
!Ni 	h->1	
!När	 ->3	
!Om 	n->1	v->1	
!Pre	c->1	
!Rös	t->1	
!San	n->1	
!Ska	l->1	
!Tac	k->1	
!Til	l->3	
!Tro	r->1	
!Tvä	r->1	
!Und	e->1	
!Vi 	b->1	f->1	h->1	s->1	ä->1	
!Äve	n->2	
" (s	e->1	
" - 	e->1	
" al	d->1	
" at	t->1	
" av	 ->1	
" bi	l->1	
" et	c->1	
" fr	a->1	
" fö	r->1	
" ge	m->1	
" gö	r->1	
" ha	r->1	
" i 	A->1	
" me	d->2	
" må	s->2	
" oc	h->6	
" på	 ->1	
" sk	a->1	
" so	m->8	
" ti	l->2	
" va	r->1	
" Är	a->1	
" är	 ->1	
"!I 	d->1	
"), 	v->1	
", "	s->1	
", a	l->1	
", b	e->1	
", d	e->2	v->1	ä->1	
", e	f->1	
", f	ö->1	
", i	 ->1	
", m	e->1	
", o	c->4	
", s	o->5	
", v	i->3	
".. 	(->1	
".Ba	r->1	
".Bå	d->1	
".De	 ->2	n->1	s->1	t->6	
".En	 ->1	
".Eu	r->1	
".Hi	s->1	
".I 	n->1	
".Ja	g->4	
".Ju	s->1	
".Ka	n->1	
".Ki	n->1	
".Nä	r->1	
".Om	 ->1	
".Or	d->1	
".Rå	d->1	
".Vi	 ->1	
"; ö	v->1	
"Ams	t->1	
"Att	 ->1	
"Big	 ->1	
"Det	 ->6	
"EU-	k->1	
"Equ	a->1	
"Eur	o->2	
"I d	e->1	
"Ja 	E->1	
"Ja,	 ->1	
"Jag	 ->2	
"Kul	t->4	
"Kvi	n->3	
"Lot	h->1	
"Med	 ->1	
"Min	d->1	
"Mis	t->1	
"Olj	e->1	
"Om 	d->1	e->1	
"Por	t->1	
"Tib	e->2	
"Ty 	h->1	
"Urb	a->1	
"aff	ä->1	
"ald	r->2	
"all	m->1	
"ang	i->3	
"avg	ö->1	
"ban	k->1	
"cou	p->1	
"den	 ->3	
"det	t->1	
"die	 ->1	
"död	a->1	
"ege	n->1	
"eko	l->1	
"en 	e->1	l->1	w->1	
"ent	r->1	
"eur	o->3	
"for	t->1	
"för	"->1	
"gem	e->1	
"gen	d->1	
"hel	l->1	
"her	o->1	
"in 	s->1	
"ind	i->1	
"inl	e->1	
"irr	e->1	
"ja 	t->1	
"kol	l->2	
"kro	n->1	
"kul	t->1	
"län	d->1	
"läs	 ->2	
"mel	l->1	
"nat	u->1	
"ne 	j->1	
"nor	m->1	
"någ	o->1	
"obe	r->1	
"orm	e->1	
"ovi	l->1	
"par	t->1	
"påp	e->1	
"ref	u->1	
"res	t->1	u->3	
"rik	t->1	
"se 	p->1	
"sha	l->1	
"ska	d->1	
"spe	c->1	
"sva	g->1	
"til	l->1	
"utv	e->1	
"utå	t->1	
"val	u->1	
"var	j->1	
"åte	r->1	
"öpp	e->1	
"öve	r->1	
'Vad	 ->1	
'eau	 ->1	
("di	e->1	
(140	9->2	
(199	7->1	8->5	9->7	
(571	3->1	
(809	5->2	
(961	4->1	
(98)	0->1	
(99)	0->2	
(A5-	0->36	
(App	l->5	
(Arb	e->1	
(B5-	0->4	
(Ben	e->1	
(Bry	s->2	
(C5-	0->7	
(CEN	)->2	
(CER	N->1	
(CNS	)->9	
(COD	)->13	
(COS	)->2	
(DA)	 ->2	
(DE)	 ->3	
(EG,	 ->1	
(EIF	)->1	
(EL)	 ->3	
(EN)	 ->34	
(ES)	 ->1	
(EU-	f->1	
(EUG	F->2	
(FI)	 ->1	
(FIP	O->1	
(FPÖ	)->1	
(FR)	 ->18	
(FUF	)->1	
(Gen	o->1	
(H-0	0->1	7->12	8->8	
(How	i->1	
(ICE	S->1	
(IFO	P->1	
(IMO	)->1	
(IT)	 ->3	
(Ihå	l->1	
(Int	e->1	
(KOM	(->8	
(Kul	t->2	
(Liv	l->2	
(NL)	 ->4	
(PPE	-->1	
(PT)	 ->16	
(Par	l->16	
(Pro	t->1	
(SEK	(->1	
(SPÖ	)->1	
(SYN	)->1	
(Sam	m->4	
(Tal	m->8	
(Uts	k->2	
(art	.->1	i->6	
(att	 ->1	
(avs	n->1	
(de 	n->1	
(det	 ->1	
(eft	e->1	
(ell	e->1	
(en 	i->1	m->1	
(fis	k->4	
(for	t->1	
(för	e->3	
(häl	s->1	
(i d	e->1	
(i s	å->1	
(inf	ö->1	
(inr	e->1	
(kod	i->2	
(kom	m->1	
(kon	s->1	
(kri	s->2	
(mai	n->2	
(mer	 ->1	
(och	 ->1	
(rec	o->1	
(råd	e->1	
(se 	a->1	
(sås	o->1	
(t.e	x->1	
(tyv	ä->1	
(ung	.->1	
(ÖVP	)->1	
(Öst	e->4	
(åte	r->1	
) "T	y->1	
) (C	5->1	
) (K	O->2	
) (S	E->1	
) (U	t->2	
) (f	ö->1	
) - 	A->1	H->1	S->1	
) 01	1->1	
) 05	5->1	
) 06	5->1	
) 15	8->1	
) 34	4->1	
) 51	9->1	
) 52	0->1	2->1	
) At	t->1	
) Bo	r->1	
) C5	-->1	
) De	 ->1	n->5	t->2	
) Ef	t->2	
) FP	Ö->1	
) Fr	u->5	å->1	
) Få	r->1	
) Fö	r->1	
) He	r->23	
) I 	S->1	d->2	g->1	s->1	
) Ja	,->1	g->14	
) Jö	r->1	
) Ko	m->1	
) Le	d->1	
) Lå	t->2	
) Mi	t->1	
) Ne	j->1	
) Nä	r->3	
) Om	 ->1	
) Se	d->1	
) Ta	c->3	l->1	
) Th	y->1	
) Ti	d->1	
) Un	d->1	
) Va	d->2	
) Ve	n->1	
) Vi	 ->2	
) ad	 ->1	
) av	 ->32	
) bä	t->1	
) ef	t->1	
) fi	n->1	
) fr	å->3	
) fö	r->5	
) ha	d->1	r->2	
) i 	G->1	e->1	h->1	ä->1	
) in	f->3	n->1	t->1	
) li	k->1	
) mi	n->1	
) oc	h->12	
) om	 ->1	
) på	 ->1	
) sa	m->1	
) si	n->1	
) so	m->2	
) tä	c->1	
) zo	n->1	
) Är	a->1	
) är	 ->2	
)(Ge	n->1	
)(Pa	r->9	
)(Ta	l->1	
)) (	U->2	f->1	
)) i	n->2	
))(G	e->1	
))(P	a->7	
)). 	V->1	
))..	 ->1	(->2	
)).F	r->1	
)).J	a->1	
))Fr	u->1	
))He	r->1	
))oc	h->1	
), b	i->1	
), d	e->1	
), m	e->1	
), o	c->2	
), r	å->1	
), s	o->2	
), t	j->1	v->1	
), v	i->1	
), ä	r->1	
). V	i->1	
).(E	N->1	
).)B	e->1	
).. 	(->1	-->1	
)..(	D->1	E->1	
).De	 ->2	t->3	
).Fr	u->1	å->1	
).Fö	r->1	
).He	r->5	
).Ja	g->3	
).Ka	n->1	
).Ko	m->1	
).Li	k->1	
).Vi	d->1	l->1	
)000	3->2	
)006	6->1	
)059	8->2	
)066	2->1	
):An	g->19	
); a	n->1	
); e	n->1	
)? H	a->1	
)And	r->2	
)Ang	å->2	
)Ans	v->1	
)Bet	ä->8	
)Det	 ->1	
)Fru	 ->8	
)För	f->1	s->1	
)Gem	e->1	
)Hea	t->1	
)Her	r->2	
)Jag	 ->3	
)Jus	t->1	
)Kon	r->1	
)Näs	t->3	
)Olj	e->1	
)Ref	o->1	
)Säk	e->1	
)Tac	k->1	
)Utt	j->1	
)].)	 ->1	
)].H	e->2	
)och	I->1	
)Åte	r->1	
, "a	f->1	
, "e	n->1	
, "n	e->1	
, "o	v->1	
, "s	e->1	
, (B	r->1	
, , 	a->1	
, 1 	p->1	
, 10	,->1	
, 11	 ->1	,->2	
, 12	 ->1	,->3	
, 13	,->1	
, 15	 ->1	,->2	
, 16	 ->1	,->1	6->1	7->1	
, 18	,->1	
, 19	9->3	
, 2 	o->1	
, 20	,->1	
, 22	,->1	
, 24	 ->1	5->1	8->1	
, 27	,->1	
, 28	,->2	
, 30	,->1	
, 31	 ->1	
, 32	,->2	
, 34	,->1	
, 36	,->1	
, 37	,->2	
, 38	,->1	
, 4,	 ->1	
, 40	,->1	
, 42	 ->2	
, 44	 ->1	
, 46	 ->1	
, 50	 ->1	0->1	
, 56	 ->1	
, 6,	 ->1	
, 7,	 ->2	
, 8,	 ->1	
, 88	 ->1	
, 9,	 ->2	
, 95	/->1	
, Al	s->1	
, Am	o->2	
, An	v->1	
, Ar	i->3	
, As	i->1	
, BN	I->1	
, Be	l->2	r->2	
, Br	e->1	o->1	y->1	
, Bu	s->1	
, Co	s->1	
, Cu	x->1	
, Da	g->1	n->1	r->1	v->1	
, Di	m->1	
, Du	b->1	
, EC	H->1	
, ED	D->1	
, EE	G->2	
, EG	-->1	
, Ef	t->1	
, Er	i->1	k->1	
, Eu	r->8	
, Ev	a->2	
, Fi	n->1	
, Fr	a->1	
, Fö	r->1	
, Ga	r->1	
, Gi	l->1	n->1	
, Gr	a->1	
, Ha	g->1	i->1	v->1	
, He	l->1	
, II	 ->1	I->1	
, IV	 ->1	
, Il	e->1	
, In	g->1	
, Ir	l->1	
, It	a->2	
, Ja	p->1	
, Jo	n->2	r->1	
, Ka	n->1	r->1	z->1	
, Ko	c->1	r->1	
, Ku	l->1	
, Kv	ä->1	
, La	 ->1	n->4	
, Le	i->1	
, Li	s->1	
, Lo	m->1	r->1	
, Lu	x->1	
, Ma	r->1	
, Mi	s->1	t->1	
, Ne	d->1	
, No	r->1	
, OL	A->1	
, Ob	e->1	
, Ol	y->1	
, PV	C->1	
, Pa	l->4	
, Pe	i->1	
, Ra	f->1	p->1	
, Re	a->1	d->1	
, Ro	t->1	
, SE	K->2	
, Sa	g->1	m->1	
, Sc	h->2	
, Sh	a->1	
, Sl	o->1	
, So	a->1	
, Sp	a->3	
, St	o->1	
, Sv	e->1	
, Ta	n->1	
, Th	y->1	
, To	m->1	t->1	
, Ty	s->3	
, Uz	b->1	
, V 	-->1	
, Vl	a->1	
, Wa	f->1	
, We	s->1	
, Wi	e->1	
, Wu	l->1	
, Wy	e->1	
, Zi	m->1	
, ac	c->2	
, ad	e->1	m->1	
, ak	t->1	
, al	b->1	d->1	l->23	
, am	b->1	
, an	a->1	d->3	f->1	g->4	n->3	s->17	t->1	v->2	
, ar	b->5	r->1	t->1	
, at	t->174	
, av	 ->23	f->1	s->5	
, ba	n->1	r->5	
, be	d->1	g->3	h->1	k->1	l->1	n->1	r->5	s->6	t->4	v->4	
, bi	d->2	l->3	
, bl	.->16	a->10	i->4	
, bo	r->9	
, br	i->3	o->1	ö->1	
, by	g->1	r->1	
, bä	r->2	s->5	
, bå	d->13	
, bö	r->19	
, ci	v->1	
, co	m->1	
, de	 ->36	c->3	l->8	m->9	n->51	r->3	s->12	t->116	
, di	a->1	f->1	s->2	
, dj	u->4	
, dr	i->1	
, du	 ->1	
, dv	s->43	
, dä	c->1	r->65	
, då	 ->27	l->1	
, dö	d->2	l->1	
, ef	f->2	t->120	
, ek	o->3	
, el	e->1	l->30	
, em	e->1	
, en	 ->81	d->1	e->3	h->1	k->1	l->19	
, er	a->1	b->1	k->1	
, et	a->1	c->2	i->1	n->1	t->37	
, eu	r->3	
, ex	a->2	e->5	i->1	
, fa	c->1	k->3	s->7	
, fi	c->2	n->10	
, fl	y->1	
, fo	l->7	r->8	
, fr	a->27	e->2	i->6	u->55	ä->12	å->20	
, fu	l->1	n->1	
, få	r->10	t->1	
, fö	d->1	r->254	
, ga	m->1	n->1	r->1	v->1	
, ge	 ->1	d->1	m->3	n->22	r->2	
, gi	v->3	
, gj	o->2	
, gl	ö->1	
, go	d->1	
, gr	a->1	u->4	ä->1	
, gu	l->1	
, gy	n->1	
, gä	l->1	
, gå	 ->2	r->4	t->1	
, gö	r->9	
, ha	 ->1	d->2	f->1	m->3	n->12	r->75	
, he	l->7	r->145	t->1	
, hj	ä->2	
, ho	p->2	s->1	t->1	
, hu	m->1	r->13	s->1	v->3	
, hy	g->1	r->1	s->1	
, hä	l->3	n->2	r->4	v->1	
, hå	l->2	
, hö	g->3	j->2	
, i 	A->1	B->1	I->1	P->1	S->1	T->1	a->7	b->5	d->22	e->19	f->9	h->3	i->1	j->2	k->2	l->5	m->4	n->1	p->3	r->4	s->43	t->1	u->1	v->6	ö->2	
, ib	l->2	
, ic	k->1	
, id	r->1	
, ig	å->1	
, in	b->3	d->1	f->9	g->4	k->15	l->2	n->13	o->15	r->1	s->3	t->74	v->2	
, ir	o->1	
, ja	 ->3	g->36	
, jo	r->2	
, ju	 ->3	s->13	
, jä	m->2	r->8	
, ka	d->2	l->3	m->1	n->37	o->1	t->1	
, ki	d->1	
, kl	a->2	
, ko	f->1	l->14	m->58	n->11	o->1	r->3	s->2	
, kr	a->3	i->2	o->2	ä->6	
, ku	l->5	n->2	r->1	
, kv	i->3	
, kä	n->2	r->48	
, la	d->2	n->2	
, le	d->5	g->3	m->1	
, li	d->1	k->33	t->1	v->2	
, lj	u->1	
, lo	k->1	
, lä	g->3	k->1	m->4	n->1	s->1	
, lå	n->7	t->4	
, lö	n->1	
, ma	k->1	n->5	r->2	t->1	
, me	d->92	l->1	n->321	r->7	s->1	
, mi	k->1	l->10	n->35	s->3	
, mo	d->3	n->1	r->2	t->7	
, mu	l->1	s->1	
, my	c->6	n->1	
, mä	n->9	
, må	 ->1	n->1	s->25	
, na	r->1	t->11	z->1	
, ne	d->3	j->1	k->1	p->1	
, ni	 ->4	
, no	g->1	r->1	
, nu	 ->6	
, ny	 ->1	a->3	l->1	
, nä	m->36	r->69	s->1	
, nå	g->29	
, nö	d->1	
, oa	k->1	n->1	v->4	
, ob	e->4	
, oc	h->668	k->8	
, of	f->1	t->1	
, ol	i->1	y->1	
, om	 ->99	d->1	e->1	f->2	v->1	
, op	p->1	
, or	d->4	e->1	g->4	
, os	t->1	v->2	
, ot	y->1	
, pa	r->7	
, pe	n->1	r->3	
, pl	a->1	u->2	
, po	l->2	
, pr	a->1	e->15	i->7	o->4	
, pu	b->1	
, på	 ->53	g->1	m->2	p->1	
, ra	p->1	s->5	
, re	a->1	g->10	k->2	n->1	s->3	v->1	
, ri	k->3	
, ro	m->1	
, rä	d->2	k->2	t->9	
, rå	d->11	
, rö	r->4	s->1	
, sa	d->2	k->2	l->1	m->31	n->1	t->1	
, se	 ->3	d->3	k->1	r->2	t->1	x->2	
, si	n->6	s->1	
, sj	u->3	ä->1	
, sk	a->22	e->2	i->1	j->1	o->1	r->4	u->18	y->1	ä->1	
, sl	u->3	ä->1	
, sm	a->1	å->1	
, sn	a->5	e->2	
, so	c->5	l->2	m->381	
, sp	a->2	e->8	o->1	
, st	a->6	i->1	o->1	r->7	y->1	å->2	ö->4	
, sv	a->2	å->1	
, sy	r->1	
, sä	g->4	k->29	l->1	r->34	
, så	 ->109	d->2	g->1	s->17	v->20	
, sö	k->1	n->1	
, t.	e->8	
, ta	c->9	k->1	l->2	r->4	
, te	o->1	
, ti	l->58	o->1	t->1	
, tj	ä->6	
, to	b->1	g->1	l->1	n->1	r->2	t->1	
, tr	a->16	e->3	o->27	å->1	
, tu	l->1	r->1	
, tv	i->3	ä->1	å->5	
, ty	 ->12	c->1	d->1	v->3	
, tä	c->1	n->1	
, tå	g->1	l->1	
, tö	m->1	
, un	d->20	g->4	i->2	
, up	p->14	
, ur	 ->3	
, ut	a->132	b->5	f->1	g->2	i->2	m->1	n->1	o->3	r->5	s->1	t->5	v->7	ö->1	
, va	d->15	l->2	n->1	r->47	t->2	
, ve	k->1	m->1	r->4	t->4	
, vi	 ->35	a->3	c->2	d->12	k->1	l->188	s->7	
, vo	n->1	r->3	
, vä	c->2	d->2	g->3	l->2	r->4	
, vå	g->1	l->1	r->6	
, yt	t->1	
, Îl	e->1	
, äg	a->2	
, än	 ->3	d->9	
, är	 ->89	a->21	l->1	
, äv	e->60	
, å 	a->1	
, ån	y->1	
, år	 ->1	
, åt	 ->1	a->1	e->17	f->1	g->1	m->7	t->1	
, ök	a->2	
, öp	p->3	
, öv	e->6	
,07 	m->1	
,2 m	i->1	
,2 o	c->1	
,2 p	r->1	
,3 p	r->1	
,4 t	r->1	
,42 	m->1	
,487	 ->1	
,5 m	i->1	
,5 p	r->2	
,6 p	r->1	
,7 p	r->1	
,8 m	i->3	
,8 t	i->1	
,9 p	r->1	
- "d	e->1	
- 'V	a->1	
- (D	E->1	
- (P	T->14	
- , 	v->1	
- 19	9->26	
- 2,	8->1	
- 31	 ->1	
- 6 	m->1	
- 80	 ->1	
- Al	t->2	
- C4	-->6	
- C5	-->14	
- Ca	m->1	
- De	n->1	
- Do	m->1	
- EU	-->1	
- Fr	u->1	
- He	r->3	
- Ka	l->1	
- Ko	m->1	
- Pa	r->1	
- Re	v->1	
- Ri	k->1	
- Rå	d->1	
- Sa	v->2	
- al	l->5	
- an	s->1	v->1	
- ar	b->1	
- at	t->27	
- av	 ->9	
- be	t->1	
- bi	d->1	
- bl	i->1	
- bö	r->1	
- ce	n->1	
- de	 ->10	l->2	n->5	s->1	t->33	
- do	c->1	
- dv	s->2	
- dä	r->2	
- då	 ->2	
- ef	t->2	
- ek	o->1	
- el	l->6	
- en	 ->8	a->1	d->1	h->1	l->1	
- et	t->3	
- ev	e->1	
- ex	e->1	i->1	
- fa	t->1	
- fi	c->1	
- fr	a->1	ä->1	å->1	
- få	 ->1	r->1	t->1	
- fö	r->16	
- ge	n->1	r->1	
- gä	l->1	
- gö	r->2	
- ha	n->1	r->9	
- ho	s->1	
- hu	r->3	
- hä	r->1	
- i 	K->1	a->1	d->1	f->1	m->1	r->1	s->3	u->1	v->1	
- id	a->1	
- in	f->2	n->1	o->2	s->1	t->10	
- ja	 ->1	,->2	g->12	
- ju	s->1	
- ka	n->1	
- kn	a->1	
- ko	m->6	n->1	s->2	
- kr	ä->1	
- li	k->1	n->1	
- ly	s->1	
- lå	t->2	
- ma	n->2	r->1	
- me	d->5	n->8	r->1	
- mi	n->1	s->1	
- mo	n->1	t->1	
- må	n->1	s->1	
- na	t->1	
- ny	 ->1	
- nä	m->3	r->3	
- nå	g->6	
- oc	h->159	k->1	
- of	f->1	
- om	 ->8	r->1	
- or	d->1	
- pa	r->1	
- pr	e->1	i->1	o->1	
- på	 ->4	m->1	
- ra	p->1	
- re	g->1	s->1	
- ri	s->1	
- rå	d->1	
- rö	r->1	
- sa	d->1	m->4	
- se	 ->1	r->2	
- si	t->1	
- sk	a->2	u->1	
- sn	a->1	e->1	
- so	m->26	
- st	a->2	o->1	
- sy	f->1	s->1	
- sä	g->1	r->1	
- så	 ->5	l->1	
- sö	k->1	
- ta	c->1	
- te	k->1	
- ti	l->3	
- tr	o->3	
- tv	e->1	
- tä	n->1	
- un	d->1	
- ut	a->7	g->1	s->1	t->1	
- va	r->2	
- ve	r->1	t->1	
- vi	 ->6	k->1	l->10	s->1	
- vä	l->1	
- Ös	t->2	
- är	 ->7	
- äv	e->10	
- åt	m->2	
- öp	p->1	
- öv	e->4	
-(EN	)->1	
-, S	a->1	
-, a	t->1	
-, d	ä->1	
-, f	ö->1	
-, i	 ->1	n->1	
-, m	e->1	
-, s	k->1	
-, t	r->1	
-, u	t->2	
-, ä	r->1	
-000	1->1	2->1	3->4	4->2	6->4	7->3	9->2	
-001	0->2	1->2	2->2	8->3	
-002	0->1	2->2	
-004	0->1	1->1	5->2	
-005	0->1	
-006	9->1	
-007	3->1	8->1	
-008	7->1	
-009	5->1	
-010	4->2	5->2	6->1	7->2	8->2	
-012	0->1	2->1	
-016	7->1	
-018	0->2	
-020	8->2	
-021	2->1	
-030	5->1	
-032	7->2	
-033	3->2	4->2	
-034	1->2	
-035	0->1	1->1	2->1	
-071	5->1	
-077	8->1	
-078	0->1	1->1	2->1	5->1	6->1	8->1	
-079	1->1	3->1	5->1	6->1	8->1	
-080	1->1	5->1	7->1	8->1	
-081	3->1	7->1	9->1	
-082	9->1	
-199	5->2	7->1	9->1	
-2 d	a->1	
-2-o	m->1	
-200	0->1	2->2	4->2	6->17	
-4 p	r->1	
-98/	0->1	
-Alp	e->1	
-Als	t->2	
-Ard	e->1	
-Atl	a->1	
-Beh	r->7	
-Car	p->1	
-Cla	u->1	
-DE)	.->1	
-DE-	 ->2	g->4	l->1	
-Del	g->1	
-Exu	p->1	
-Fin	a->3	
-Fra	n->2	
-Har	r->1	
-Hei	n->1	
-I);	 ->1	
-II)	 ->1	
-Isr	a->1	
-Jør	g->2	
-Kee	s->1	
-Le 	B->1	
-Loi	r->1	
-Man	n->1	
-Mat	h->2	
-Nor	m->1	
-PM 	s->1	
-Pla	t->4	
-Rob	l->1	
-Rom	a->1	
-SS:	s->1	
-Sha	r->1	
-She	i->5	
-Syr	i->1	
-aff	ä->3	
-alb	a->1	
-ana	l->6	
-anp	a->1	
-avt	a->3	
-avv	i->1	
-bel	o->1	
-ben	e->5	
-bes	t->1	
-bil	a->1	d->1	e->1	
-bis	t->1	
-bri	t->1	
-bud	g->1	
-bug	g->1	
-dam	m->1	
-dan	s->1	
-de-	F->2	L->1	
-dir	e->3	
-dis	k->2	
-dom	s->22	
-eff	e->1	
-el-	S->1	
-enh	e->1	
-er 	r->1	
-fal	l->1	
-fon	d->1	
-fos	s->1	
-fra	n->1	
-fre	e->3	
-frå	g->1	
-för	d->19	e->1	k->2	s->1	
-gem	e->1	
-gen	o->1	
-gru	p->20	
-how	 ->1	
-ini	t->2	
-ins	t->5	
-int	ä->2	
-irl	ä->1	
-isr	a->1	
-kan	a->1	
-kat	a->3	
-kol	i->1	
-kom	m->3	
-kor	t->20	
-kos	t->1	
-kri	s->3	t->1	
-lag	s->1	
-lan	d->1	
-led	a->2	
-lek	s->1	
-lit	e->2	
-lob	b->1	
-län	d->5	
-mai	l->1	
-man	t->1	
-med	b->4	e->1	l->1	
-met	a->1	
-nat	i->1	
-niv	å->1	
-not	i->1	
-nyt	t->1	
-oly	c->1	
-omr	å->8	
-ord	f->1	
-org	a->3	
-pos	i->1	
-pro	g->25	t->2	
-ram	p->1	
-ras	i->1	
-reg	e->1	i->6	
-rät	t->4	
-råd	e->4	
-sho	p->1	
-sit	u->1	
-ska	n->1	
-soc	i->2	
-spr	i->3	
-sta	t->13	
-sti	p->1	
-sto	p->1	
-str	u->1	
-stö	d->2	
-sys	t->1	
-sän	d->3	
-tal	 ->1	e->7	s->1	
-tes	t->1	
-tex	t->1	
-tra	n->1	
-upp	d->1	
-utv	i->1	
-van	 ->1	
-vär	l->1	
-zon	 ->1	e->2	
. (E	L->1	N->23	
. (F	I->1	R->12	
. (P	T->1	
. -(	E->1	
. 11	 ->1	,->1	.->6	
. 12	.->6	0->1	
. 13	.->1	
. 15	.->2	
. 17	.->1	
. 19	.->1	
. 20	.->1	
. 21	.->2	
. 7 	l->1	
. 7)	.->1	
. Al	l->1	
. Av	 ->1	
. De	 ->2	n->9	r->1	s->3	t->39	
. Dä	r->6	
. Då	 ->2	
. Ef	t->2	
. En	 ->5	l->1	
. Eq	u->1	
. Et	t->1	
. Eu	r->4	
. Fo	g->1	
. Fr	a->1	u->2	ä->1	
. Fö	l->1	r->2	
. Gu	t->1	
. Ha	n->1	
. He	r->3	
. Ho	n->1	
. Hu	r->1	
. Hä	r->3	
. Hå	l->1	
. I 	r->1	s->1	
. In	g->1	i->1	t->1	
. Ja	g->10	
. Ko	m->1	s->1	
. Kä	r->1	
. Lå	t->1	
. Ma	n->2	
. Me	n->15	
. Ne	d->1	
. Ni	 ->1	
. Nä	s->1	
. Oc	h->4	
. Of	f->1	
. Om	 ->1	
. Pa	r->1	
. Pr	o->1	
. På	 ->1	
. Rå	d->1	
. Sk	o->1	ä->1	
. So	m->2	
. Sy	r->1	
. Så	 ->2	
. Ta	c->1	
. Ti	l->1	
. US	A->1	
. Va	r->3	
. Vi	 ->10	,->1	l->1	
. Vå	r->2	
. Wa	l->1	
. ai	d->1	
. an	s->1	
. ar	b->1	t->1	
. at	t->12	
. av	 ->1	s->2	
. be	t->1	
. de	 ->1	n->3	s->2	t->2	
. en	 ->1	h->1	
. er	t->1	
. et	t->3	
. fo	r->1	
. få	r->1	
. fö	r->8	
. ge	n->1	
. gr	a->1	
. gö	r->1	
. ho	s->1	
. hu	r->1	
. i 	M->1	d->1	e->1	p->1	
. id	é->1	
. in	f->1	n->1	o->1	t->3	
. ja	g->1	
. kr	i->1	
. ku	n->1	
. kä	n->1	
. ma	n->2	
. me	d->2	n->1	
. mi	n->1	t->2	
. nä	r->5	t->1	
. oc	h->2	
. ol	j->2	
. om	 ->3	
. på	 ->3	
. sk	a->2	o->1	
. so	f->1	
. sp	e->1	
. st	o->1	
. sä	k->1	
. tr	a->1	
. un	d->1	
. ut	f->1	
. va	d->1	r->2	
. vi	 ->1	
. Äm	n->1	
. Än	d->1	n->1	
. Äv	e->1	
. Åt	g->1	
. Ös	t->1	
. än	n->1	
. är	 ->1	
. ös	t->1	
." Ä	r->1	
."De	t->1	
."I 	d->1	
."Ja	g->1	
."Me	d->1	
.(Ap	p->5	
.(Ar	b->1	
.(DA	)->2	
.(DE	)->2	
.(EL	)->2	
.(EN	)->10	
.(ES	)->1	
.(FR	)->6	
.(IT	)->3	
.(Ih	å->1	
.(Li	v->2	
.(NL	)->4	
.(PT	)->1	
.(Pa	r->5	
.(Pr	o->1	
.(Sa	m->4	
.(Ta	l->7	
.) H	e->3	
.) T	a->1	
.).D	e->1	
.).H	e->1	
.)An	d->2	s->1	
.)Be	t->8	
.)Fr	u->5	
.)Fö	r->2	
.)Ge	m->1	
.)He	a->1	r->1	
.)Ju	s->1	
.)Ol	j->1	
.)Re	f->1	
.)Sä	k->1	
.)Åt	e->1	
., d	e->1	
., f	r->1	
., ä	v->1	
.- (	D->1	P->10	
.- D	e->1	
.- F	r->1	
.- H	e->2	
.. (	E->16	F->10	
.. -	(->1	
.. D	e->1	
.. F	r->1	ö->1	
.. H	e->1	
.. P	r->1	
.. T	a->1	
.. V	i->1	
..(D	A->2	E->2	
..(E	L->1	N->5	S->1	
..(F	R->5	
..(I	T->1	
..(N	L->3	
..(T	a->5	
..).	D->1	
...(	T->5	
...)	.->1	
....	(->1	
...F	r->1	
...H	e->1	
...L	å->1	
..Fr	u->1	
..He	r->5	
..Lå	t->1	
..Ta	c->1	
..Vi	 ->1	
.00.	(->2	)->2	D->1	F->2	O->1	S->3	T->2	
.05 	o->1	
.1 d	å->1	
.1 i	 ->3	
.1 o	c->2	
.1 v	i->1	
.1 ö	v->1	
.1) 	e->1	
.1.1	 ->1	
.1.F	ö->1	
.1.V	i->1	
.12.	0->1	
.14 	e->1	
.15 	m->1	
.18 	m->1	
.199	8->1	
.2 i	 ->5	
.2 o	c->1	
.2).	K->1	
.25.	)->1	
.3 E	G->1	
.3 b	l->1	
.3 i	n->1	
.3, 	n->1	
.30,	 ->1	
.3; 	d->1	
.4 i	n->1	
.4.D	e->1	
.4.F	ö->1	
.50 	o->1	
.55)	U->1	
.8 i	 ->1	
.90 	p->1	
.?An	s->1	
.Acc	e->1	
.Ahe	r->1	
.Akt	i->1	
.Ald	r->1	
.All	a->21	d->1	m->4	t->18	
.Alt	e->2	
.Ame	r->1	
.Ams	t->1	
.And	r->4	
.Ang	å->1	
.Anh	å->1	
.Anl	e->1	
.Ann	a->4	
.Ans	e->1	v->3	
.Ant	a->2	
.Anv	ä->1	
.Ara	b->1	
.Arb	e->2	
.Art	i->2	
.Att	 ->22	a->1	
.Av 	4->1	a->5	b->2	d->13	e->1	s->2	v->2	
.Avb	r->1	
.Avg	å->1	
.Avs	a->1	e->1	l->13	
.Bak	o->2	
.Bar	a->4	
.Bed	r->2	ö->2	
.Bef	o->1	
.Bek	v->1	
.Ber	e->2	o->1	
.Bes	l->3	
.Bet	r->6	ä->16	
.Bev	i->1	
.Bil	i->1	l->2	t->2	
.Bis	t->1	
.Bla	n->7	
.Bor	d->2	
.Bos	ä->1	
.Bre	t->1	
.Bri	s->3	t->1	
.Bry	s->1	
.Bud	g->1	
.Byg	g->1	
.Bäs	t->1	
.Båd	a->5	
.CSU	:->1	
.Cen	t->2	
.Cor	p->1	
.Cun	h->1	
.DEB	A->1	
.Dag	e->3	l->2	
.Dal	a->1	
.Dan	m->1	
.De 	1->2	a->7	b->5	d->3	e->2	f->20	g->4	h->10	i->1	k->11	l->2	m->7	n->7	o->2	p->3	r->1	s->22	t->5	u->4	v->3	ä->4	å->2	
.Del	s->1	v->1	
.Den	 ->180	n->48	
.Der	a->1	
.Des	s->56	
.Det	 ->789	,->1	a->1	s->1	t->196	
.Dir	e->7	
.Dis	k->1	
.Doc	k->2	
.Dok	u->1	
.Dom	s->2	
.Där	 ->10	a->2	e->9	f->91	i->3	m->4	u->1	v->1	
.Då 	d->1	f->3	g->1	h->2	k->7	m->1	o->1	s->2	v->2	ä->2	ö->1	
.EG-	d->3	
.EKS	G->1	
.EU 	m->1	ä->1	
.EU-	k->2	o->1	
.Eff	e->5	
.Eft	e->36	
.Eko	n->2	
.Eme	l->8	
.En 	a->15	b->3	d->6	f->4	g->1	k->5	m->2	r->4	s->9	u->1	v->7	ö->2	
.Enb	a->1	
.End	a->9	
.Enk	e->1	
.Enl	i->31	
.Er 	a->1	
.Erf	a->2	
.Eri	k->4	
.Ert	 ->1	
.Ett	 ->43	
.Eur	o->51	
.Eve	n->1	
.Exc	e->1	
.Exe	m->1	
.Exp	e->2	
.FEO	 ->1	
.FPÖ	 ->2	:->2	
.Fac	k->3	
.Fak	t->4	
.Far	l->1	
.Fas	c->1	
.Fel	a->1	
.Fem	 ->1	
.Fin	a->2	n->2	
.Fle	r->4	
.Flo	r->3	
.Fol	k->2	
.For	s->2	
.Fra	m->8	n->2	
.Fre	d->1	
.Fri	h->1	
.Fru	 ->54	t->1	
.Frå	g->34	n->2	
.Fyr	t->1	
.Får	 ->1	
.Föl	j->5	
.För	 ->165	b->2	d->3	e->14	h->3	l->1	m->1	p->1	s->25	t->2	u->7	v->4	ä->1	
.Gem	e->3	
.Gen	e->1	o->25	
.Ger	 ->1	
.Giv	e->2	
.Gol	a->1	
.Gra	t->1	
.Gre	k->2	
.Gru	n->1	p->2	
.Gäl	l->1	
.Gå 	h->1	
.Gör	 ->2	
.Had	e->2	
.Hai	d->1	
.Han	 ->16	d->3	s->2	
.Har	 ->3	
.Hel	a->3	t->2	
.Her	r->268	
.His	t->2	
.Hit	 ->3	t->2	
.Hon	 ->3	
.Hop	p->1	
.Hul	t->1	
.Hur	 ->24	u->1	
.Huv	u->7	
.Hyc	k->1	
.Hän	d->2	
.Här	 ->28	m->1	o->1	
.Hög	e->1	
.I A	m->1	
.I E	u->4	
.I F	r->1	
.I H	e->1	
.I I	r->2	t->1	
.I N	e->1	
.I R	a->1	
.I T	i->1	y->1	
.I a	l->3	n->3	p->1	r->1	v->3	
.I b	e->4	
.I d	a->17	e->51	i->1	
.I e	g->4	n->10	t->2	
.I f	l->1	o->1	r->6	ö->6	
.I g	å->2	
.I j	u->1	
.I k	l->1	o->3	
.I l	i->6	
.I m	i->2	o->4	å->1	
.I n	o->2	ä->2	
.I o	c->4	
.I p	a->1	r->2	
.I r	a->2	e->7	ä->1	å->1	
.I s	a->3	i->2	j->4	l->2	t->10	y->2	å->3	
.I t	j->1	
.I u	p->1	t->1	
.I v	a->2	e->1	i->6	o->1	ä->2	å->6	
.I ä	n->1	
.I ö	v->3	
.Ibl	a->3	
.Idé	n->1	
.Ill	e->1	
.Imm	i->1	
.Ind	u->1	
.Inf	ö->4	
.Ing	a->1	e->11	
.Ini	t->1	
.Inn	e->2	
.Ino	m->10	
.Inr	e->2	ä->1	
.Ins	a->2	
.Int	e->12	
.Irl	a->1	
.Isr	a->1	
.Ita	l->1	
.Ja 	e->1	t->1	
.Ja,	 ->3	
.Jac	k->1	q->1	
.Jag	 ->765	
.Jon	c->1	
.Jor	d->1	
.Ju 	m->1	
.Jus	t->9	
.Jäm	f->1	s->1	
.Kaf	o->1	
.Kan	 ->10	s->6	
.Kar	l->1	
.Kat	a->1	
.Kin	n->3	
.Kna	p->1	
.Koc	h->1	
.Kod	e->1	
.Kom	 ->1	m->102	p->1	
.Kon	k->13	s->5	v->1	
.Kor	t->2	
.Kos	o->1	t->3	
.Kra	v->3	
.Kul	t->7	
.Kva	n->1	
.Kvi	n->1	
.Kär	a->4	n->2	
.La 	R->1	
.Lan	d->1	g->1	
.Led	a->2	n->1	
.Lik	a->3	r->1	s->6	v->1	
.Lit	t->1	
.Liv	s->3	
.Lyc	k->2	
.Lyn	n->1	
.Läg	g->2	
.Län	d->1	
.Lån	 ->1	g->1	
.Låt	 ->48	
.Maj	o->1	
.Mal	t->2	
.Man	 ->52	n->1	
.Mar	g->1	k->4	
.Max	i->2	
.Med	 ->29	a->4	b->3	g->1	l->9	
.Mel	l->3	
.Men	 ->189	,->2	t->1	
.Mer	 ->3	
.Mil	j->1	
.Min	 ->27	a->16	n->1	s->1	
.Mit	t->2	
.Mor	a->1	
.Mot	 ->8	
.Myl	l->1	
.Myn	d->3	
.Män	n->4	
.Mär	k->1	
.Måh	ä->1	
.Mål	e->2	
.Mån	g->10	
.Möj	l->2	
.Nat	i->3	u->14	
.Nej	,->1	
.Ni 	a->1	b->3	f->3	h->7	k->7	l->1	m->4	s->5	t->2	v->2	
.Nie	l->1	
.Niv	å->1	
.Nor	m->1	
.Nu 	a->2	b->1	f->2	h->7	k->2	m->1	t->1	v->2	ä->7	å->1	
.Num	e->1	
.Nuv	a->1	
.Nya	 ->1	
.Nyl	i->1	
.När	 ->64	
.Näs	t->1	
.Någ	o->2	r->2	
.Nåj	a->1	
.Nöd	v->1	
.OK,	 ->1	
.OLA	F->2	
.OMR	Ö->2	
.Oav	s->2	
.Obe	r->2	
.Och	 ->60	
.Ock	s->2	
.Off	e->2	
.Oft	a->1	
.Om 	5->1	E->1	S->2	a->3	b->1	d->22	e->4	f->1	g->2	i->1	j->2	k->5	l->1	m->10	n->6	p->2	r->2	s->2	t->2	u->1	v->22	
.Omr	ö->15	
.Onö	d->1	
.Ord	 ->1	e->3	f->7	
.Ork	a->2	
.Oro	n->1	v->1	
.Ors	a->2	
.Oz 	h->1	
.PPE	-->2	
.Par	a->1	l->21	
.Per	s->4	
.Pla	n->1	s->2	
.Plä	d->1	
.Por	t->2	
.Pre	c->5	s->1	
.Pro	b->8	c->2	d->5	g->1	j->2	
.Pun	k->2	
.På 	a->1	d->19	e->1	g->1	l->1	m->3	o->2	p->1	s->10	u->1	v->2	
.Rap	p->3	
.Ras	i->1	
.Rea	k->1	
.Red	a->3	
.Ref	o->6	
.Reg	e->4	i->1	
.Ren	t->2	
.Res	t->2	u->5	
.Ret	r->1	
.Rev	i->2	
.Rik	a->1	t->3	
.Ris	k->1	
.Rop	e->1	
.Rot	h->2	
.Rum	ä->1	
.Räk	n->1	
.Rät	t->2	
.Råd	e->16	
.Sam	h->2	m->7	o->1	t->14	
.San	n->5	
.Sav	e->2	
.Sch	r->1	u->1	ü->1	
.Sed	a->15	
.Set	t->1	
.Sis	t->2	
.Sit	u->3	
.Sju	 ->1	
.Sjä	l->2	
.Ska	d->1	l->3	
.Sko	t->1	
.Sku	l->4	
.Sky	d->1	
.Slu	t->38	
.Små	 ->1	f->1	
.Sna	b->1	r->1	
.Soc	i->3	
.Som	 ->42	l->3	
.Sta	b->1	t->8	
.Sto	r->4	
.Str	a->1	u->1	ä->1	
.Stä	m->1	
.Stå	l->1	
.Stö	d->6	r->4	
.Sub	v->2	
.Sve	p->1	
.Syf	t->6	
.Syr	i->1	
.Säg	 ->1	
.Säk	e->1	
.Sär	s->2	
.Så 	b->1	d->3	e->2	f->1	h->1	j->3	k->2	l->4	n->1	s->4	t->1	v->6	ä->3	
.Såd	a->2	
.Sål	e->4	
.Sån	g->1	
.Sås	o->2	
.Såv	ä->1	
.TV-	b->1	
.Ta 	d->1	
.Tac	k->28	
.Tad	z->1	
.Tal	a->1	
.Tan	k->3	
.Ter	r->1	
.The	a->2	
.Thy	s->1	
.Tid	i->1	
.Til	l->37	
.Tit	t->1	
.Ton	g->1	
.Top	p->2	
.Tor	v->2	
.Tra	n->2	
.Tre	 ->1	
.Tro	r->1	t->16	v->1	
.Trä	d->1	
.Tus	e->1	
.Tvä	r->3	
.Två	 ->2	
.Ty 	e->1	i->1	s->1	u->1	v->3	
.Tyd	l->1	
.Tyv	ä->9	
.Tän	k->1	
.Und	a->3	e->27	
.Ung	d->1	e->2	
.Uni	o->5	
.Upp	e->1	f->1	g->3	r->1	
.Ur 	d->2	e->1	p->1	
.Uta	n->3	
.Utb	i->2	
.Utd	e->1	
.Ute	s->1	
.Utf	o->2	ö->1	
.Utg	i->1	
.Uti	f->1	
.Utm	a->2	
.Utn	ä->1	
.Uts	k->2	
.Utv	e->1	i->1	
.Vad	 ->58	a->1	
.Val	e->3	
.Van	 ->1	l->1	
.Var	 ->7	e->2	f->11	j->5	
.Vem	 ->2	s->2	
.Ver	k->1	
.Vet	e->2	
.Vi 	a->25	b->36	d->8	e->2	f->26	g->8	h->90	i->13	j->1	k->56	l->4	m->78	o->1	p->2	r->6	s->39	t->17	u->8	v->53	ä->29	ö->1	
.Via	 ->1	
.Vid	 ->12	a->7	
.Vik	t->1	
.Vil	j->1	k->10	l->5	
.Vin	d->1	
.Vis	s->13	
.Vit	b->3	
.Von	 ->1	
.Vär	d->1	
.Väs	t->2	
.Vår	 ->14	a->7	t->5	
.Wor	l->1	
.Ytt	e->3	
.a. 	a->2	b->1	d->1	e->2	f->5	g->2	i->2	k->1	m->1	n->3	o->2	p->1	s->3	u->1	v->1	
.d. 	Ö->1	ö->1	
.d.,	 ->1	
.ex.	 ->20	
.g.a	.->1	
.k. 	a->1	i->1	s->2	
.kom	m->1	
.m. 	a->2	d->1	i->1	ä->2	
.m.,	 ->1	
.m.O	c->1	
.o.m	.->7	
.Än 	e->3	
.Änd	a->1	r->14	å->4	
.Änn	u->1	
.Änt	l->1	
.Är 	I->1	d->11	k->1	r->1	s->1	
.Ära	d->3	
.Äve	n->31	
.Å E	D->1	
.Å a	n->10	
.Å e	n->2	
.År 	1->4	2->1	
.Åre	t->1	
.Åta	g->1	
.Åte	r->2	
.Åtg	ä->2	
.ÖVP	 ->1	
.Ögo	n->2	
.Öka	d->1	
.Öst	e->2	
.Öve	r->2	
.Övr	i->1	
/00 	-->1	
/00)	 ->1	:->1	
/001	2->1	3->1	
/008	3->1	
/009	0->1	
/010	6->2	
/016	9->2	
/019	4->2	
/022	8->1	
/024	0->2	
/031	8->1	
/035	2->1	
/037	0->2	1->2	
/080	3->1	5->1	
/082	5->2	
/1/1	9->2	
/199	8->2	9->39	
/200	0->26	
/212	3->1	7->1	
/3 a	v->1	
/35/	E->4	
/409	 ->1	
/43.	T->1	
/55/	E->2	
/591	/->2	
/60/	9->1	
/71 	a->1	
/71/	E->1	
/728	/->1	
/75 	o->1	
/92 	o->1	
/95.	F->1	
/98 	-->1	
/98-	9->1	
/99 	(->1	-->1	b->1	o->2	
/99)	 ->2	:->18	A->2	
/99.	J->1	
/EG 	a->1	o->2	s->1	u->1	
/EG,	 ->3	
/EKS	G->2	
/Eur	o->1	
/NGL	-->2	
/Nor	d->2	
/Oil	-->1	
/den	 ->1	
/ell	e->1	
/hal	v->1	
/int	ä->1	
/rik	e->1	
/sam	m->1	
/år)	?->1	
/år,	 ->1	
0 - 	1->3	C->2	d->1	
0 00	0->11	
0 En	l->1	
0 an	s->1	
0 ar	b->2	r->1	
0 at	t->1	
0 ba	r->1	
0 bi	l->1	
0 de	t->1	
0 do	l->1	m->1	
0 dö	d->1	
0 el	l->2	
0 en	s->1	
0 eu	r->1	
0 fr	a->1	å->4	
0 få	g->2	
0 fö	r->1	
0 gu	l->1	
0 gå	n->1	
0 ha	n->1	r->2	
0 he	k->1	
0 i 	a->3	f->4	
0 in	n->3	
0 ja	n->1	
0 ju	n->1	r->1	
0 ka	n->1	
0 ki	l->4	
0 km	 ->2	,->1	.->1	
0 lä	g->1	
0 me	d->2	
0 mi	l->17	n->2	
0 mo	t->1	
0 ny	a->1	
0 nä	r->1	
0 oc	h->7	
0 ol	i->1	
0 pr	o->37	
0 på	 ->1	
0 ri	m->1	
0 sk	a->1	u->1	
0 so	m->2	
0 st	å->1	
0 ti	b->1	
0 to	n->10	
0 ut	a->2	
0 va	r->1	
0 º 	C->1	
0 än	d->7	
0 är	 ->5	
0 år	 ->7	.->2	s->1	
0 åt	g->1	
0" s	o->1	
0" t	i->2	
0".D	e->1	
0".V	i->1	
0(CN	S->2	
0(CO	D->3	
0) a	v->20	
0) f	r->1	ö->1	
0) o	c->1	
0).F	r->1	
0).J	a->1	
0):A	n->1	
0, 1	2->1	
0, 2	2->1	
0, 3	2->1	
0, 4	6->1	
0, d	ä->1	
0, f	ö->1	
0, i	 ->1	
0, m	o->1	å->1	
0, o	c->1	
0, s	k->1	å->1	
0, ä	v->1	
0- o	c->1	
0-20	0->17	
0-bu	g->1	
0-pr	o->4	
0-ta	l->9	
0.(S	a->2	
0.)A	n->1	
0.)O	l->1	
0.25	.->1	
0.4.	F->1	
0.De	n->1	t->5	
0.Fa	s->1	
0.Fr	u->1	
0.Fö	r->2	
0.Ja	g->2	
0.Ko	m->1	
0.Ma	n->1	
0.Me	n->1	
0.OM	R->1	
0.Sa	m->1	
0.St	o->1	r->1	
0.Ti	l->1	
0.Tr	a->1	
0.Vi	 ->1	
0/19	9->4	
0/20	0->3	
0/92	 ->1	
0/99	 ->2	)->2	
00 -	 ->4	
00 0	0->6	
00 E	n->1	
00 a	r->3	t->1	
00 b	a->1	i->1	
00 d	o->1	
00 f	å->2	ö->1	
00 h	a->3	e->1	
00 i	n->2	
00 k	i->4	m->4	
00 l	ä->1	
00 m	e->1	i->4	o->1	
00 n	ä->1	
00 o	c->4	l->1	
00 p	r->1	å->1	
00 s	k->2	o->1	t->1	
00 t	i->1	o->10	
00 u	t->1	
00 v	a->1	
00 ä	n->4	r->4	
00 å	r->1	
00" 	s->1	t->2	
00".	D->1	V->1	
00) 	a->20	f->2	o->1	
00).	F->1	J->1	
00):	A->1	
00, 	d->1	f->1	i->1	m->2	s->1	ä->1	
00-2	0->17	
00-b	u->1	
00-p	r->4	
00-t	a->4	
00.(	S->2	
00.)	A->1	O->1	
00.D	e->5	
00.F	a->1	r->1	ö->2	
00.J	a->2	
00.M	a->1	e->1	
00.O	M->1	
00.S	a->1	t->2	
00.T	i->1	r->1	
00.V	i->1	
000 	-->3	E->1	a->3	b->1	f->3	h->3	i->2	k->4	l->1	m->3	n->1	o->2	p->1	s->3	t->11	u->1	v->1	ä->4	
000"	 ->3	.->2	
000)	 ->22	.->2	
000,	 ->7	
000-	2->17	b->1	p->4	t->4	
000.	D->4	F->2	J->2	M->2	V->1	
0001	/->1	
0002	/->1	
0003	 ->2	/->4	
0004	/->2	
0006	/->4	
0007	/->3	
0009	/->2	
000N	ä->1	
001 	ä->1	
001,	 ->1	
001/	2->1	
0010	/->2	
0011	/->2	
0012	(->1	/->2	
0013	(->1	
0018	/->3	
002 	(->1	f->1	
002)	 ->2	
002,	 ->2	
002.	 ->1	H->1	M->1	P->1	V->1	
002/	2->1	
0020	/->1	
0022	/->2	
003 	-->2	
003/	2->4	
003?	H->1	
004 	i->1	
004.	D->1	K->1	
004/	1->1	2->1	
0040	/->1	
0041	/->1	
0045	/->2	
0050	/->1	
006 	[->1	f->2	g->1	k->1	l->1	o->1	s->1	t->2	å->1	
006,	 ->5	
006.	D->2	E->1	F->1	H->1	J->2	M->1	T->1	
006/	0->2	2->2	
0066	 ->1	
0069	/->1	
007,	 ->1	
007/	2->3	
0073	/->1	
0078	/->1	
008 	t->2	
0083	 ->1	
0087	/->1	
009/	2->2	
0090	(->1	
0095	/->1	
00Nä	s->1	
01 ä	n->1	
01, 	m->1	
01/2	0->1	
01/9	9->1	
010 	e->1	
010/	2->2	
0104	/->2	
0105	/->2	
0106	(->2	/->1	
0107	/->2	
0108	/->2	
011/	2->2	
0113	 ->1	
012 	e->1	
012(	C->1	
012/	2->2	
0120	/->1	
0122	/->1	
013(	C->1	
0167	/->1	
0169	(->2	
018/	2->2	9->1	
0180	/->2	
0194	(->2	
02 (	K->1	
02 f	a->1	
02) 	-->2	
02, 	k->1	s->1	
02. 	J->1	
02.H	e->1	
02.M	i->1	
02.P	å->1	
02.V	i->1	
02/2	0->1	
020/	1->1	
0208	/->2	
0212	/->1	
022/	2->2	
0228	(->1	
0240	(->2	
03 -	 ->2	
03(C	N->1	
03/2	0->4	
0305	/->1	
0318	(->1	
0327	/->2	
0333	/->2	
0334	/->2	
0341	/->2	
0350	/->1	
0351	/->1	
0352	(->1	/->1	
0370	(->2	
0371	(->2	
03?H	e->1	
04 i	n->1	
04.D	e->1	
04.K	o->1	
04/1	9->3	
04/2	0->1	
040/	9->1	
041/	9->1	
045/	0->1	2->1	
05 i	 ->1	
05 o	c->1	
05 t	i->1	
05(C	N->1	
05/1	9->3	
05/9	9->1	
050/	2->1	
0550	 ->1	
0598	 ->2	
06 [	K->1	
06 f	ö->2	
06 g	ä->1	
06 k	o->1	
06 l	i->1	
06 o	c->1	
06 s	å->1	
06 t	a->1	o->1	
06 å	t->1	
06(C	O->2	
06, 	f->1	m->1	n->1	s->2	
06.D	e->2	
06.E	n->1	
06.F	r->1	
06.H	e->1	
06.J	a->2	
06.M	a->1	
06.T	a->1	
06/0	0->2	
06/1	9->1	
06/2	0->2	
0652	 ->1	
066 	-->1	
0662	 ->1	
069/	1->1	
07 m	i->1	
07, 	r->1	
07/1	9->2	
07/2	0->3	
07/9	9->1	
0715	/->1	
073/	1->1	
0778	/->1	
078/	1->1	
0780	/->1	
0781	/->1	
0782	/->1	
0785	/->1	
0786	/->1	
0788	/->1	
0791	/->1	
0793	/->1	
0795	/->1	
0796	/->1	
0798	/->1	
08 t	o->2	
08/1	9->4	
08/9	9->1	
0801	/->1	
0803	(->1	
0805	(->1	/->1	
0807	/->1	
0808	/->1	
0813	/->1	
0817	/->1	
0819	/->1	
0825	(->2	
0829	/->1	
083 	(->1	
087/	1->1	
09 o	c->1	
09/2	0->2	
090(	C->1	
094/	1->2	
095/	1->3	
0Näs	t->1	
1 00	0->2	
1 40	0->1	
1 an	g->1	
1 då	 ->1	
1 ef	t->1	
1 fr	å->3	
1 ge	r->1	
1 i 	A->1	E->1	a->1	k->1	r->1	
1 ja	n->9	
1 ju	l->1	n->1	
1 ma	j->1	r->3	
1 me	n->1	
1 mi	l->1	
1 oc	h->18	k->1	
1 om	 ->1	
1 pr	o->7	
1 ri	s->1	
1 se	p->1	
1 st	a->2	
1 ur	 ->1	v->1	
1 ut	a->1	
1 vi	l->1	
1 än	t->1	
1 är	 ->1	
1 år	 ->1	
1 öv	e->1	
1(CO	D->2	
1) e	f->1	
1, 1	2->2	
1, 2	 ->1	
1, 4	,->1	
1, a	t->1	
1, f	ö->1	
1, m	å->1	
1, o	c->1	
1, s	k->1	
1,2 	o->1	p->1	
1,3 	p->1	
1,4 	t->1	
1-2 	d->1	
1-om	r->4	
1-re	g->5	
1-st	a->2	
1.00	.->4	
1.1 	d->1	o->2	ö->1	
1.1.	F->1	V->1	
1.3 	E->1	b->1	i->1	
1.3,	 ->1	
1.3;	 ->1	
1.55	)->1	
1.Al	t->1	
1.Ex	c->1	
1.Fö	r->1	
1.Ja	g->1	
1.Ku	l->1	
1.Vi	 ->1	
1/19	9->5	
1/20	0->3	
1/3 	a->1	
1/99	)->4	
1/EG	 ->1	
1/EK	S->2	
10 0	0->2	
10 e	l->2	
10 f	r->1	
10 i	 ->1	
10 j	a->1	
10 k	a->1	
10 m	i->2	
10 p	r->4	
10 r	i->1	
10 s	o->1	
10 ä	n->1	r->1	
10 å	r->1	
10, 	1->1	
10.K	o->1	
10/2	0->2	
100 	d->1	k->1	m->1	o->1	p->1	ä->4	
104/	1->2	
105 	i->1	t->1	
105/	1->2	
106(	C->2	
106/	1->1	
107/	1->2	
108/	1->2	
11 i	 ->1	
11 j	a->2	
11 m	i->1	
11 o	c->1	
11 s	t->1	
11, 	1->2	f->1	
11,3	 ->1	
11.0	0->3	
11.A	l->1	
11.E	x->1	
11.K	u->1	
11/2	0->2	
110 	i->1	
113 	-->1	
115 	m->1	
12 e	n->1	
12 f	r->1	
12 i	n->1	
12 j	a->1	
12 m	i->1	å->1	
12 o	c->1	
12 p	r->1	
12 s	t->1	
12(C	O->1	
12, 	1->2	d->1	t->1	
12.0	0->7	
12/1	9->1	
12/2	0->2	
12/9	9->3	
120 	m->1	
120/	9->1	
122/	1->1	
123 	p->1	
123(	C->1	
1244	 ->1	.->2	
125 	m->1	
1260	/->1	
127(	C->1	
13 (	E->1	
13 -	 ->1	
13 0	0->1	
13 A	m->1	
13 f	e->1	
13 i	 ->2	
13 j	a->1	
13 n	y->1	
13 o	k->1	
13 p	r->2	
13 s	a->1	
13 ä	r->1	
13(C	N->1	
13, 	2->2	
13.0	5->1	
13.F	ö->1	
13/1	9->1	
13/9	9->1	
130 	d->1	
133.	2->1	
138.	4->1	
14 e	u->1	
14 f	e->5	
14 l	e->1	
14 m	e->5	
14 o	c->1	
14 s	e->1	
14 t	i->1	
14, 	e->1	
14/1	9->1	
140 	j->1	
1409	4->2	
143 	o->1	
15 a	v->1	
15 m	a->2	i->1	
15 o	l->2	m->1	
15 p	r->3	
15 r	ä->1	
15 s	e->1	t->1	
15 å	r->1	
15, 	1->2	
15.0	0->2	
15/9	8->1	
150 	g->1	o->1	
158 	-->1	i->1	
158)	.->1	
158.	1->1	
16 0	0->1	
16 o	c->3	
16 p	e->1	r->1	
16 r	a->1	
16) 	s->1	
16, 	2->1	
164 	r->1	
166 	e->1	
167 	m->3	
167/	1->1	
169(	C->2	
17 d	e->2	
17 m	i->1	
17 o	c->1	k->1	
17 s	å->1	
17, 	1->1	s->1	
17.3	0->1	
17.S	l->1	
17/9	9->1	
170 	m->1	
174 	t->1	
1762	 ->1	.->1	
18 d	e->1	
18 h	ä->1	
18 i	 ->1	
18 m	i->2	å->1	
18 n	o->3	
18(S	Y->1	
18, 	2->1	
18/2	0->2	
18/9	8->1	
180 	m->1	
180/	1->2	
19 -	 ->1	
19 d	e->1	
19 m	a->1	
19 p	r->1	
19 s	o->1	
19 ä	r->1	
19.5	0->1	
19/9	9->1	
1917	 ->1	
1923	,->1	
193 	o->1	
1930	-->1	
194(	C->2	
194.	D->1	
1945	.->1	
1948	.->1	
195 	m->1	
1957	 ->1	.->1	
1967	 ->5	,->1	
1969	 ->1	
1976	 ->1	
1977	 ->1	
1982	,->1	.->1	
1986	 ->2	.->1	
1989	,->1	
1990	 ->1	.->1	
1991	 ->3	
1992	 ->3	,->1	
1993	 ->3	,->1	-->2	.->1	?->1	
1994	 ->4	,->1	-->1	
1995	 ->6	,->2	-->1	
1996	 ->11	,->2	.->5	
1997	 ->20	)->1	,->2	.->10	/->7	?->1	N->1	
1998	 ->18	)->3	,->3	-->2	.->3	/->4	
1999	 ->67	"->1	)->21	,->7	-->2	.->14	/->13	:->1	
1:a 	å->1	
2 (K	O->1	
2 - 	C->3	v->1	
2 00	0->1	
2 40	0->1	
2 av	 ->1	
2 bl	a->1	i->1	
2 da	g->1	
2 de	c->1	
2 el	l->1	
2 en	l->1	
2 eu	r->1	
2 fa	k->1	
2 fr	å->2	
2 ha	r->1	
2 i 	A->2	S->1	a->3	f->3	r->1	s->1	t->1	
2 in	n->2	
2 ja	n->1	
2 mi	l->5	
2 må	n->1	
2 oc	h->9	
2 pr	o->4	
2 pu	n->1	
2 ri	k->1	
2 sk	r->1	
2 so	m->2	
2 st	a->1	
2 un	d->1	
2 up	p->1	
2 år	s->1	
2(CN	S->1	
2(CO	D->1	
2) -	 ->2	
2) f	ö->1	
2).K	a->1	
2, 1	1->1	3->1	5->1	
2, 2	4->2	
2, 3	7->2	
2, d	e->1	v->1	
2, e	l->1	n->1	
2, f	r->1	
2, i	 ->2	
2, k	o->1	
2, l	ä->1	
2, s	k->1	o->2	
2, t	i->1	r->1	
2, v	i->2	
2,48	7->1	
2,5 	m->1	
2,6 	p->1	
2,8 	m->1	
2-om	r->3	
2-st	ö->1	
2. J	a->1	
2.00	.->7	
2.1 	i->1	
2.2 	i->1	
2.De	t->1	
2.He	r->1	
2.I 	e->1	
2.Is	r->1	
2.Ja	g->1	
2.Ma	n->1	
2.Me	n->1	
2.Mi	n->1	
2.På	 ->1	
2.Vi	 ->1	
2.Äv	e->1	
2/19	9->3	
2/20	0->5	
2/43	.->1	
2/99	 ->2	)->1	.->1	
20 -	 ->1	
20 0	0->1	
20 e	u->1	
20 f	r->1	
20 g	å->1	
20 m	i->3	
20 n	y->1	
20 p	r->3	
20 º	 ->1	
20 ä	n->1	
20 å	r->5	
20, 	2->1	
20.2	5->1	
20/1	9->1	
20/9	9->1	
200 	0->4	å->1	
2000	 ->24	"->5	)->24	,->7	-->26	.->10	N->1	
2001	 ->1	,->1	
2002	 ->2	)->2	,->2	.->5	
2003	?->1	
2004	 ->1	.->2	
2006	 ->11	,->5	.->9	
2007	,->1	
2010	 ->1	
2012	 ->1	
208/	1->2	
21 j	a->1	u->1	
21 o	c->1	m->1	
21 s	t->1	
21 ä	r->1	
21 å	r->1	
21.0	0->1	
21.5	5->1	
212/	1->1	
2123	(->1	
2127	(->1	
21:a	 ->1	
22 -	 ->1	
22 a	v->1	
22 r	i->1	
22, 	2->1	i->1	v->1	
22,5	 ->1	
22.Ä	v->1	
22/1	9->1	
22/2	0->2	
226 	i->1	
228(	C->1	
23 d	e->1	
23 i	n->1	
23 p	e->1	
23(C	O->1	
23, 	e->1	
23,7	 ->1	
24 n	y->2	
24 o	c->1	k->1	
24 p	r->1	
240(	C->2	
244 	o->1	
244.	I->1	J->1	
245 	o->1	
248,	 ->1	
25 g	r->1	
25 m	e->1	i->2	
25 o	m->1	
25 p	r->7	
25 t	i->1	
25(C	N->2	
25.)	J->1	
25.D	e->1	
250 	m->1	
255 	i->4	
26 "	p->1	
26 i	 ->1	n->1	
26 m	e->1	
26 n	o->1	
26 o	c->1	
26 p	r->1	
260/	9->1	
262 	e->1	
27 d	e->1	
27 f	a->1	
27 l	ä->1	
27 o	c->1	
27 p	r->2	
27(C	O->1	
27, 	3->1	
27/1	9->2	
28 f	r->1	
28 j	u->1	
28 n	y->1	
28 p	r->1	
28(C	N->1	
28, 	3->2	
28/E	G->1	
280 	i->4	
280.	4->1	
28:e	 ->1	
29 d	ö->1	
29 f	r->1	
29 l	ä->1	
29 m	i->1	
29, 	3->1	
29/9	9->1	
299.	2->2	
3 (C	O->1	
3 (E	U->1	
3 - 	C->3	
3 00	0->5	
3 Am	s->1	
3 EG	-->1	
3 av	 ->2	
3 bl	i->1	
3 de	c->1	
3 fe	b->2	
3 fr	å->1	
3 fö	r->1	
3 ha	r->1	
3 hö	r->1	
3 i 	E->1	d->1	f->1	
3 in	n->1	t->1	
3 ja	n->2	
3 ma	j->1	
3 ny	a->1	
3 oc	h->4	
3 ok	t->2	
3 om	 ->1	
3 pe	r->2	
3 pr	o->6	
3 pu	n->1	
3 sa	m->1	
3 ut	e->1	
3 är	 ->1	
3(CN	S->2	
3(CO	S->1	
3, 1	9->1	
3, 2	8->2	
3, 7	,->1	
3, e	f->1	
3, n	å->1	
3,7 	p->1	
3,8 	m->1	t->1	
3,9 	p->1	
3-19	9->2	
3-4 	p->1	
3-li	t->2	
3.05	 ->1	
3.1)	 ->1	
3.2 	o->1	
3.8 	i->1	
3.Fr	å->1	
3.Fö	r->1	
3.I 	ö->1	
3.Om	 ->1	
3.Ty	d->1	
3/19	9->4	
3/20	0->4	
3/75	 ->1	
3/99	)->2	
30 d	o->1	
30 f	r->1	
30 i	 ->1	n->1	
30 j	u->1	
30 m	e->1	i->1	
30 o	c->1	
30 p	r->3	
30, 	3->1	o->1	
30-t	a->1	
300 	s->1	
305/	1->1	
31 f	r->1	
31 j	a->1	
31 m	a->2	
31 o	c->2	
314 	l->1	
318(	S->1	
32 m	i->1	
32, 	2->1	3->2	
32.J	a->1	
327/	1->2	
33 0	0->2	
33 a	v->1	
33 f	r->1	ö->1	
33 i	 ->1	
33 o	c->1	
33.2	 ->1	
33/1	9->2	
332,	 ->1	
333/	1->2	
334/	1->2	
34 i	 ->1	
34 s	k->1	
34 t	i->1	
34 å	r->1	
34, 	3->1	
34.1	.->1	
34/1	9->2	
341/	1->2	
344 	-->1	
35 f	r->1	
35 m	i->5	
35.S	å->1	
35/E	G->4	
350 	m->1	
350/	1->1	
351/	1->1	
352(	C->1	
352/	1->1	
36 f	r->1	
36, 	3->1	
367 	0->1	
37 f	r->1	
37 i	 ->1	
37 p	r->1	
37, 	4->2	
37.2	 ->1	
37/6	0->1	
370 	m->1	
370(	C->2	
371(	C->2	
38 f	r->1	ö->1	
38 o	c->2	
38, 	4->1	
38.4	.->1	
38: 	f->1	
39 f	r->1	
39 i	 ->1	
39 p	r->1	
39, 	4->1	
3: f	ö->1	
3; d	e->1	
3?Fr	å->1	
3?He	r->1	
4 - 	C->1	
4 00	0->1	
4 c 	i->1	
4 en	 ->1	
4 et	t->1	
4 eu	r->1	
4 fe	b->5	
4 fr	å->1	
4 ha	r->1	
4 i 	E->2	a->1	d->3	
4 in	l->1	t->1	
4 ju	n->2	
4 le	d->1	
4 li	k->1	
4 me	d->5	
4 ny	a->2	
4 nä	r->1	
4 oc	h->8	
4 ok	t->1	
4 pr	o->5	
4 rö	s->1	
4 se	p->1	
4 sk	a->1	
4 ti	l->2	
4 tr	i->1	
4 tu	s->1	
4 år	 ->1	
4(CO	D->2	
4, 1	1->2	
4, 3	6->1	
4, 6	,->1	
4, e	l->1	
4, f	ö->1	
4, k	o->1	
4, o	c->1	
4-00	1->1	
4-02	1->1	
4-03	5->3	
4-07	1->1	
4-19	9->1	
4.1.	1->1	
4.2)	.->1	
4.De	 ->1	t->2	
4.Fö	r->1	
4.I 	d->3	
4.Ja	g->2	
4.Ko	m->1	
4/19	9->8	
4/20	0->1	
4/55	/->2	
4/72	8->1	
40 f	r->1	
40 j	u->1	
40 m	i->2	
40 p	r->6	
40 å	r->3	
40(C	N->2	
40, 	4->1	
40/9	9->1	
400 	0->1	k->3	m->2	
409 	o->1	
4094	/->2	
41 f	r->1	
41 p	r->1	
41 r	i->1	
41 u	r->1	
41/1	9->2	
41/9	9->1	
410 	f->1	
42 f	r->1	
42 i	 ->1	
42 m	i->1	
42 o	c->2	
43 h	ö->1	
43 o	m->1	
43.F	r->1	
43.T	y->1	
44 -	 ->1	
44 f	r->1	
44 o	c->3	
44.I	 ->1	
44.J	a->1	
45 a	v->1	
45 c	e->1	
45 f	r->1	
45 g	ä->1	
45 o	c->1	
45, 	d->1	
45. 	D->1	
45."	I->1	
45.F	r->1	
45.H	e->1	
45.V	i->1	
45/0	0->1	
45/2	0->1	
46 o	c->2	
462 	u->1	
47 g	ä->1	
48 g	ä->1	
48 i	 ->2	n->1	
48 ä	n->1	
48, 	2->1	
48.D	e->1	
487 	m->1	
5 (e	n->1	
5 - 	8->1	
5 00	0->3	8->2	
5 av	 ->2	
5 ce	n->1	
5 fr	å->3	
5 gr	a->1	
5 gä	l->2	
5 ha	r->1	
5 i 	A->1	E->1	f->3	
5 in	t->1	
5 ko	m->1	
5 ma	r->2	
5 me	s->1	
5 mi	l->16	n->1	
5 mo	r->1	
5 oc	h->4	
5 ok	t->1	
5 ol	i->2	
5 om	 ->2	r->1	
5 pr	o->14	
5 ri	k->1	
5 rä	c->1	
5 se	p->1	
5 sl	u->1	
5 st	a->1	
5 ti	l->4	
5 vi	s->1	
5 år	.->2	s->1	
5(CN	S->3	
5)Ut	t->1	
5, 1	6->2	
5, d	e->1	ä->1	
5, n	å->1	
5, o	c->2	
5, u	t->1	
5,5 	p->1	
5,8 	m->1	
5-00	0->16	1->8	2->3	4->4	5->1	6->1	7->2	8->1	9->1	
5-01	0->9	2->2	6->1	8->2	
5-02	0->2	
5-03	0->1	2->2	3->4	4->2	
5-19	9->1	
5. D	ä->1	
5."I	 ->1	
5.)J	u->1	
5.00	.->2	
5.4 	i->1	
5.De	s->1	
5.Em	e->1	
5.Fr	u->1	å->1	
5.He	r->1	
5.Så	d->1	
5.Vi	 ->1	
5/00	 ->1	
5/1/	1->2	
5/19	9->4	
5/20	0->1	
5/35	/->1	
5/95	.->1	
5/98	-->1	
5/99	)->3	
5/EG	 ->4	,->2	
50 -	 ->1	
50 0	0->1	
50 g	u->1	
50 i	 ->1	
50 m	i->4	
50 o	c->2	
50 p	r->3	
50, 	s->1	
50- 	o->1	
50-t	a->2	
50/1	9->1	
50/2	0->1	
500 	0->1	
51/1	9->1	
519 	-->1	
52 -	 ->1	
52 i	 ->1	
52(C	N->1	
52/1	9->1	
520 	-->1	f->1	
522 	-->1	
53 p	r->1	
540 	m->1	
55 i	 ->3	n->1	
55 m	o->1	
55 p	r->1	
55)U	t->1	
55/E	G->2	
550 	-->1	
56 p	r->1	
56, 	s->1	
57 (	m->1	
57,5	 ->1	
57.E	u->1	
5713	/->1	
58 -	 ->1	
58 i	 ->1	
58).	D->1	
58.1	 ->1	
591/	E->2	
598 	-->2	
5b k	a->1	
5b-o	m->1	
5b.D	e->1	
6 "p	å->1	
6 - 	C->1	s->1	
6 00	0->1	
6 [K	O->1	
6 de	c->1	
6 ef	t->1	
6 el	l->1	
6 em	o->1	
6 fr	å->2	
6 fö	r->2	
6 gä	l->1	
6 ha	d->1	r->1	
6 i 	E->1	a->1	f->6	h->1	u->1	
6 in	d->1	
6 ko	m->1	
6 li	g->1	
6 lå	g->1	
6 me	d->1	
6 mi	l->1	
6 no	v->1	
6 oc	h->15	
6 om	 ->1	
6 pe	r->1	
6 pr	o->6	
6 ra	d->1	
6 så	 ->1	
6 ta	s->1	
6 to	t->1	
6 va	r->1	
6 vi	l->1	
6 är	 ->1	
6 år	s->2	
6 åt	e->1	
6(CO	D->2	
6) s	a->1	
6, 2	0->1	
6, 3	8->1	
6, 7	,->1	
6, f	ö->1	
6, h	a->1	
6, m	e->1	
6, n	ä->1	
6, s	o->3	
6, t	a->1	
6, v	i->1	
6,07	 ->1	
6.De	t->3	
6.En	l->2	
6.Fr	å->1	
6.He	r->1	
6.Ja	g->3	
6.Ma	n->1	
6.Me	n->1	
6.Oc	h->1	
6.Så	 ->1	
6.Ta	c->1	
6.År	 ->1	
6/00	)->2	
6/19	9->1	
6/20	0->2	
6/35	/->3	
6/71	 ->1	/->1	
6/99	)->2	
60 0	0->1	
60 f	r->1	
60-t	a->1	
60/9	2->1	9->1	
600 	b->1	
614/	1->1	
62 -	 ->1	
62 e	u->1	
62 i	 ->1	
62 u	n->1	p->1	
62.M	a->1	
64 r	ö->1	
652 	-->1	
66 -	 ->1	
66 e	m->1	
662 	-->1	
67 0	0->1	
67 h	a->1	
67 i	 ->2	
67 m	e->1	i->3	
67 o	c->2	
67, 	o->1	
67/1	9->1	
68 a	t->1	
685/	9->1	
69 o	c->1	
69(C	O->2	
69/1	9->1	
7 (a	v->1	
7 (m	e->1	
7 - 	d->1	i->2	
7 00	0->1	
7 de	c->4	
7 dä	r->1	
7 fa	l->1	
7 fr	å->1	
7 fö	r->2	
7 gr	a->1	
7 gä	l->1	
7 ha	r->2	
7 hä	r->1	
7 i 	A->3	a->2	b->1	d->1	f->3	u->1	v->1	
7 le	d->1	
7 ly	d->1	
7 lä	n->1	
7 me	d->1	
7 mi	l->7	
7 nä	m->1	
7 oc	h->11	
7 ok	t->1	
7 om	 ->1	
7 pr	o->5	
7 på	 ->2	
7 så	 ->1	
7 tr	o->2	
7 up	p->1	
7 är	 ->1	
7 år	s->1	
7(CO	S->1	
7) 0	6->1	
7)..	 ->1	
7, 1	8->1	
7, 3	4->1	
7, 4	2->2	
7, 8	8->1	
7, 9	,->1	
7, d	v->1	
7, m	e->1	
7, o	c->2	m->1	
7, r	e->1	
7, s	o->1	å->1	
7, v	a->1	
7,2 	m->1	
7,42	 ->1	
7,5 	p->1	
7.- 	D->1	
7.. 	(->1	
7.1 	i->1	
7.2 	i->2	
7.30	,->1	
7.Be	t->1	
7.De	t->2	
7.Eu	r->1	
7.Fr	å->1	
7.I 	v->1	
7.Ma	n->1	
7.Nu	 ->1	
7.Se	d->1	
7.Sl	u->1	
7.Vi	 ->2	
7/01	9->2	
7/03	5->1	7->4	
7/19	9->6	
7/20	0->3	
7/60	/->1	
7/99	 ->1	)->2	
70 a	n->1	
70 m	i->2	
70 p	r->1	
70(C	O->2	
700 	a->1	h->1	o->2	
71 a	n->1	
71(C	O->2	
71/E	G->1	
713/	1->1	
715/	9->1	
728/	E->1	
73,9	 ->1	
73/1	9->1	
74 t	u->1	
75 -	 ->1	
75 m	i->2	
75 o	m->1	
76 e	l->1	
76 p	r->1	
762 	u->1	
762.	M->1	
77 -	 ->1	
77 m	i->1	
778/	9->1	
78/1	9->1	
78/9	9->1	
780/	9->1	
781/	9->1	
782/	9->1	
785/	9->1	
786/	9->1	
788/	9->1	
79/4	0->1	
791/	9->1	
793/	9->1	
795/	9->1	
796/	9->1	
798/	9->1	
7?De	 ->1	
7Näs	t->1	
8 - 	1->1	C->3	
8 46	2->1	
8 at	t->1	
8 be	h->1	
8 de	c->1	
8 fr	å->3	
8 fö	r->1	
8 go	d->1	
8 gä	l->1	
8 ha	d->1	
8 hä	n->1	
8 i 	E->2	b->1	d->1	f->2	
8 in	n->1	
8 ju	l->1	
8 ko	s->1	
8 mi	l->6	
8 må	n->1	
8 no	v->3	
8 ny	a->1	
8 oc	h->12	
8 pr	o->1	
8 re	g->1	s->1	
8 sk	a->1	
8 ti	l->2	
8 to	n->2	
8 un	d->1	
8 ut	b->1	g->1	
8 va	r->2	
8 än	d->1	
8 är	 ->4	
8(CN	S->1	
8(SY	N->1	
8) 5	1->1	2->2	
8).D	e->1	
8)06	6->1	
8, 2	4->1	7->1	
8, 3	0->1	2->1	
8, 4	4->1	
8, 9	,->1	
8, S	E->2	
8, d	ä->1	
8, s	å->1	
8-20	0->2	
8-98	/->1	
8. D	e->1	
8.1 	i->1	
8.4.	D->1	
8.De	t->1	
8.Pr	e->1	
8.St	o->1	
8/01	0->2	6->2	
8/03	1->1	
8/19	9->5	
8/20	0->2	
8/59	1->2	
8/98	 ->1	
8/99	)->4	
8/EG	,->1	
80 e	n->1	
80 i	 ->4	
80 m	i->1	
80 p	r->11	
80 ä	n->1	
80 å	t->1	
80.4	.->1	
80/1	9->2	
80/9	9->1	
801/	9->1	
803(	C->1	
805(	C->1	
805/	9->1	
807/	9->1	
808/	9->1	
8095	/->2	
81 o	c->5	
81 p	r->1	
81.1	 ->3	.->2	
81.3	 ->3	,->1	;->1	
81/9	9->1	
813/	9->1	
817/	9->1	
819/	9->1	
82 h	a->1	
82 i	n->1	
82) 	f->1	
82, 	d->1	e->1	f->1	l->1	t->1	
82.I	 ->1	s->1	
82/9	9->1	
825(	C->2	
829/	9->1	
83 (	C->1	
83 p	r->1	
85 o	c->2	
85 p	r->1	
85 t	i->1	
85/9	5->1	9->1	
86 h	a->1	
86 i	 ->2	
86 o	c->1	
86 p	r->1	
86.Å	r->1	
86/9	9->1	
87 m	i->1	
87, 	8->1	
87.1	 ->1	
87.2	 ->1	
87/1	9->1	
88 i	 ->1	
88 o	c->1	
88 ä	r->1	
88/5	9->2	
88/9	9->1	
89 i	 ->1	
89 t	i->1	
89, 	1->1	
8: f	o->1	
8:e 	å->1	
9 (H	o->1	
9 - 	1->20	3->1	C->7	
9 an	t->3	
9 av	s->1	
9 be	t->1	
9 de	c->1	p->1	
9 dä	r->1	
9 dö	d->1	
9 er	h->1	
9 fa	l->1	
9 fe	b->1	
9 fr	a->2	å->3	
9 go	d->1	
9 ha	d->1	m->1	r->3	
9 i 	M->1	f->1	h->1	s->1	v->1	
9 in	n->1	t->1	
9 jä	m->1	
9 ka	n->1	
9 ko	m->2	
9 ku	n->1	
9 lä	n->1	
9 ma	r->1	
9 mi	l->3	n->1	
9 nä	r->1	
9 oc	h->6	k->1	
9 om	 ->1	
9 pr	o->3	ä->1	
9 ra	s->1	
9 sk	a->1	
9 so	m->1	
9 ti	l->2	
9 up	p->2	
9 ut	 ->1	
9 va	r->2	
9 vi	s->1	
9 är	 ->1	
9 äv	e->1	
9 år	s->1	
9 öv	e->1	
9".B	å->1	
9(CO	D->2	
9) 0	1->1	5->1	
9) 1	5->1	
9) 3	4->1	
9) a	v->12	
9) f	r->2	
9) o	c->1	
9).K	o->1	
9)00	0->2	6->1	
9)05	9->2	
9):A	n->18	
9)An	g->2	
9, 1	9->1	
9, 3	1->1	
9, 4	0->1	
9, a	n->1	v->1	
9, b	e->1	
9, d	v->1	
9, f	ö->1	
9, h	a->1	
9, n	ä->1	
9, o	c->2	
9-20	0->2	
9. V	i->1	
9..(	F->1	
9.1 	v->1	
9.2 	i->2	
9.50	 ->1	
9.De	 ->1	s->1	t->1	
9.En	 ->1	
9.Eu	r->1	
9.Fr	å->1	
9.Fö	r->2	
9.Ja	g->2	
9.Ko	m->1	
9.Un	d->1	
9.Vi	 ->1	
9/00	1->2	8->1	9->1	
9/02	2->1	4->2	
9/08	0->2	2->2	
9/19	9->1	
9/20	0->2	
9/21	2->2	
9/40	9->1	
9/99	)->2	
90 d	e->1	ö->1	
90 p	r->4	
90 u	t->1	
90(C	O->1	
90-t	a->1	
90.D	e->1	
91 e	f->1	
91 g	e->1	
91 o	c->1	
91 p	r->1	
91/9	9->1	
91/E	K->2	
917 	o->1	
92 o	c->1	
92 s	k->1	o->1	
92 å	r->1	
92, 	e->1	
92/4	3->1	
923,	 ->1	
93 h	a->1	
93 o	c->2	
93 p	e->1	
93 u	t->1	
93, 	1->1	
93-1	9->2	
93.O	m->1	
93/7	5->1	
93/9	9->1	
930-	t->1	
93?F	r->1	
94 e	t->1	
94 h	a->1	
94 n	ä->1	
94 o	c->2	
94 p	r->2	
94(C	O->2	
94, 	f->1	k->1	
94-1	9->1	
94.D	e->1	
94/1	9->2	
94/5	5->2	
94/7	2->1	
945.	F->1	
948.	D->1	
95 (	e->1	
95 h	a->1	
95 i	 ->1	
95 k	o->1	
95 m	i->3	
95 r	i->1	
95 s	l->1	
95 t	i->1	
95 å	r->1	
95, 	n->1	o->1	
95-1	9->1	
95.F	r->1	
95/1	/->2	9->1	
95/3	5->1	
95/9	9->1	
957 	(->1	
957.	E->1	
96 -	 ->1	
96 e	f->1	
96 h	a->1	
96 i	 ->1	
96 l	å->1	
96 o	c->1	
96 v	a->1	i->1	
96 ä	r->1	
96 å	r->2	
96, 	h->1	v->1	
96.D	e->1	
96.E	n->1	
96.J	a->1	
96.M	e->1	
96.O	c->1	
96/3	5->3	
96/7	1->2	
96/9	9->1	
9614	/->1	
967 	h->1	i->1	m->1	o->2	
967,	 ->1	
969 	o->1	
97 (	a->1	
97 -	 ->1	
97 d	ä->1	
97 f	ö->1	
97 h	a->1	ä->1	
97 i	 ->1	
97 l	y->1	
97 o	c->5	m->1	
97 p	å->1	
97 t	r->2	
97 u	p->1	
97 ä	r->1	
97 å	r->1	
97) 	0->1	
97, 	m->1	v->1	
97.-	 ->1	
97..	 ->1	
97.B	e->1	
97.D	e->2	
97.I	 ->1	
97.M	a->1	
97.N	u->1	
97.S	e->1	
97.V	i->2	
97/0	1->2	3->5	
97/9	9->1	
976 	e->1	
977 	-->1	
97?D	e->1	
97Nä	s->1	
98 -	 ->3	
98 g	o->1	
98 h	a->1	
98 k	o->1	
98 m	i->1	
98 o	c->6	
98 r	e->1	
98 s	k->1	
98 u	n->1	t->2	
98 v	a->2	
98 ä	r->2	
98) 	5->3	
98)0	6->1	
98, 	S->2	d->1	
98-2	0->2	
98-9	8->1	
98. 	D->1	
98.P	r->1	
98.S	t->1	
98/0	1->4	3->1	
98/9	9->1	
982,	 ->1	
982.	I->1	
986 	h->1	o->1	
986.	Å->1	
989,	 ->1	
99 (	H->1	
99 -	 ->27	
99 a	n->3	v->1	
99 b	e->1	
99 d	ä->1	
99 e	r->1	
99 f	r->2	
99 g	o->1	
99 h	a->5	
99 i	 ->3	n->1	
99 j	ä->1	
99 k	a->1	o->2	u->1	
99 n	ä->1	
99 o	c->5	m->1	
99 p	r->1	
99 r	a->1	
99 s	k->1	
99 t	i->1	
99 u	p->2	t->1	
99 v	a->2	i->1	
99 ä	v->1	
99 å	r->1	
99 ö	v->1	
99".	B->1	
99) 	0->2	1->1	3->1	a->12	f->2	o->1	
99).	K->1	
99)0	0->3	5->2	
99):	A->18	
99)A	n->2	
99, 	a->1	b->1	d->1	h->1	n->1	o->2	
99-2	0->2	
99. 	V->1	
99..	(->1	
99.2	 ->2	
99.D	e->3	
99.E	n->1	u->1	
99.F	r->1	ö->2	
99.J	a->2	
99.K	o->1	
99.U	n->1	
99.V	i->1	
99/0	0->4	2->3	8->4	
99/2	1->2	
990 	u->1	
990.	D->1	
991 	e->1	g->1	o->1	
992 	s->2	å->1	
992,	 ->1	
993 	h->1	o->1	u->1	
993,	 ->1	
993-	1->2	
993.	O->1	
993?	F->1	
994 	e->1	h->1	o->2	
994,	 ->1	
994-	1->1	
995 	(->1	h->1	k->1	r->1	s->1	å->1	
995,	 ->2	
995-	1->1	
996 	-->1	e->1	h->1	i->1	l->1	o->1	v->2	ä->1	å->2	
996,	 ->2	
996.	D->1	E->1	J->1	M->1	O->1	
997 	(->1	-->1	d->1	f->1	h->2	i->1	l->1	o->6	p->1	t->2	u->1	ä->1	å->1	
997)	 ->1	
997,	 ->2	
997.	-->1	.->1	B->1	D->2	I->1	M->1	N->1	V->2	
997/	0->7	
997?	D->1	
997N	ä->1	
998 	g->1	h->1	k->1	o->6	r->1	s->1	u->3	v->2	ä->2	
998)	 ->3	
998,	 ->3	
998-	2->2	
998.	 ->1	P->1	S->1	
998/	0->4	
999 	-->26	a->4	d->1	e->1	f->2	g->1	h->5	i->4	j->1	k->4	n->1	o->4	p->1	r->1	s->1	t->1	u->3	v->3	ä->1	å->1	ö->1	
999"	.->1	
999)	 ->17	.->1	0->3	
999,	 ->7	
999-	2->2	
999.	 ->1	.->1	D->3	E->2	F->3	J->1	K->1	U->1	V->1	
999/	0->11	2->2	
999:	 ->1	
99: 	"->1	
9: "	j->1	
: "A	t->1	
: "D	e->4	
: "J	a->1	
: "M	i->1	
: "O	m->1	
: "a	l->1	
: "d	e->1	
: "h	e->1	
: "i	n->1	
: "j	a->1	
: "v	a->1	
: An	l->1	m->1	
: Ar	b->1	t->1	
: As	t->1	
: At	t->1	
: De	 ->3	s->1	t->5	
: Ef	t->1	
: Er	i->1	
: Eu	r->1	
: Fi	n->1	r->1	
: Fl	o->1	
: Fr	i->2	ä->1	
: Fö	r->5	
: Ge	m->1	n->1	
: Gr	e->1	
: Ha	m->1	n->1	
: Ho	l->1	
: I 	b->1	m->1	s->1	
: In	g->1	
: Ja	g->7	
: Jo	r->1	
: Ko	c->1	m->4	n->1	
: Kä	n->1	r->1	
: Ma	i->1	
: Na	r->1	
: Ny	t->1	
: Nä	r->3	
: Om	 ->1	
: Os	l->1	
: Pa	r->1	
: Po	r->1	
: På	 ->1	
: Re	v->1	
: St	a->1	ö->1	
: Tu	r->1	
: Tå	g->1	
: Un	d->1	i->1	
: Ut	n->1	v->1	
: Va	d->3	p->1	
: Ve	m->3	
: Vi	 ->7	
: an	g->1	t->3	
: at	t->8	
: ba	l->1	
: be	s->1	
: de	 ->2	f->1	l->1	n->8	t->13	
: di	r->1	
: du	b->1	
: dä	r->1	
: en	 ->8	
: et	t->2	
: fo	r->2	
: fr	å->2	
: fö	r->12	
: ge	m->1	n->1	
: gö	r->1	
: ha	n->2	
: hu	r->4	
: hö	g->1	
: i 	F->1	l->1	r->1	
: in	o->1	s->2	
: ja	,->1	g->4	
: ka	n->1	
: ko	m->3	
: ma	n->1	
: me	d->2	
: mi	n->1	
: nu	 ->1	
: nä	r->2	
: om	 ->4	
: op	e->1	
: pa	r->1	
: pr	o->1	
: rä	t->1	
: sk	a->1	
: sy	s->1	
: ta	n->1	
: ti	l->1	
: to	l->1	
: un	d->1	
: up	p->1	
: ut	b->2	n->1	v->1	
: va	d->2	r->3	
: ve	m->3	
: vi	 ->10	l->2	
: vå	g->1	r->1	
: Är	 ->1	
: Äv	e->1	
: Åt	g->2	
: Öp	p->1	
: å 	e->1	
: ön	s->1	
:Ang	å->19	
:Den	 ->1	
:Det	 ->1	
:För	 ->1	o->1	
:a å	r->1	
:e r	a->2	
:e å	r->1	
:s (	f->1	
:s B	a->1	
:s E	u->1	
:s a	n->1	r->3	
:s b	e->3	i->2	u->2	y->1	
:s d	e->1	i->1	o->1	
:s e	g->1	k->1	u->1	
:s f	r->2	ö->2	
:s g	a->1	e->1	i->1	
:s h	a->1	e->1	
:s i	n->6	
:s k	o->1	u->1	
:s l	a->1	i->2	
:s m	e->3	i->2	
:s n	u->1	ä->1	
:s o	c->3	m->1	r->2	
:s p	a->1	o->3	
:s r	e->2	
:s s	a->1	i->1	t->5	ä->1	
:s t	e->1	j->1	
:s u	p->1	r->1	t->1	
:s v	e->1	
:s.L	e->1	
; Da	n->1	
; Ja	v->1	
; al	l->1	
; an	n->1	t->1	
; ar	t->1	
; at	t->3	
; av	 ->1	
; b)	 ->1	
; de	 ->1	n->4	s->4	t->22	
; dä	r->1	
; då	 ->1	
; en	 ->5	d->1	l->1	
; fi	s->1	
; fo	r->1	
; fr	i->1	
; fö	r->7	
; hä	r->1	
; i 	F->1	d->1	e->1	
; in	f->1	l->1	s->1	t->1	
; ja	g->4	
; ko	m->1	
; lo	j->1	
; ma	n->1	
; me	n->2	
; mi	n->2	
; oc	h->5	
; pu	n->3	
; sa	m->1	
; sk	o->1	
; sl	u->1	
; un	d->1	
; vi	 ->5	d->1	
; än	n->1	
; å 	e->1	
; öv	e->1	
? 21	 ->1	
? De	n->2	
? Ha	r->2	
? In	t->1	
? Me	d->1	
? Oc	h->1	
? Rå	d->1	
?"Ja	 ->1	
?, r	å->2	
?- (	P->3	
?. (	E->8	F->1	
?.(E	N->2	
?.He	r->2	
?Ans	e->3	l->1	
?Att	 ->2	
?Av 	t->1	
?Avs	l->1	
?Bor	d->1	
?Dag	e->1	
?De 	h->1	p->1	t->1	
?Den	 ->8	
?Des	s->1	
?Det	 ->18	t->1	
?Där	 ->1	f->2	
?Eft	e->1	
?Ell	e->1	
?End	a->1	
?Enl	i->1	
?Ett	 ->3	
?Eur	o->2	
?Fin	n->1	
?Fol	k->1	
?Fru	 ->6	
?Frå	g->3	
?För	 ->7	s->1	
?Har	 ->4	
?Hem	l->1	
?Her	r->15	
?Hur	 ->10	
?Här	 ->1	m->1	
?I F	r->1	
?I d	a->2	
?I e	r->1	
?I f	j->1	
?I m	e->1	
?I s	å->1	
?I v	i->1	
?Ini	t->1	
?Int	e->1	
?Ja,	 ->2	
?Jag	 ->21	
?Jo 	d->1	
?Jo,	 ->3	
?Kan	 ->2	s->3	
?Kol	l->1	
?Kom	m->6	
?Kär	a->1	
?Man	 ->1	
?Men	 ->2	a->1	
?Nat	u->1	
?Nej	,->5	.->1	
?Ni 	k->2	n->1	
?När	 ->3	
?Näs	t->1	
?Och	 ->3	
?Oli	k->1	
?Om 	i->2	
?Par	l->1	
?Pro	b->1	
?På 	d->1	v->1	
?RIN	A->1	
?Reg	e->1	
?Sed	a->1	
?Ser	i->1	
?Sku	l->3	
?Som	 ->2	
?Sva	r->1	
?Tac	k->1	
?Til	l->1	
?Tyc	k->1	
?Tän	k->1	
?Utg	i->1	
?Vad	 ->7	
?Vem	 ->2	
?Vet	s->1	
?Vi 	b->2	f->1	h->1	m->2	s->2	t->1	ä->2	
?Vil	k->13	
?Vis	s->2	
?Är 	d->8	h->1	i->1	v->1	
?Äve	n->2	
A - 	o->1	
A OC	H->1	
A at	t->1	
A el	l->1	
A ha	r->3	
A på	 ->1	
A va	r->1	
A) D	e->1	
A) V	e->1	
A, K	a->1	
A, e	f->1	
A, s	o->1	
A-in	s->1	
A-st	ö->1	
A. G	u->1	
A.Ja	g->1	
A.Vi	 ->1	
A5-0	0->27	1->9	
A:s.	L->1	
ABB 	A->1	
ABB-	A->2	
ABC 	d->1	
ADR)	 ->1	
AF g	ö->1	
AF i	 ->2	
AF k	a->1	o->1	
AF s	k->1	
AF, 	E->1	d->1	e->1	k->1	s->2	v->1	ö->1	
AF.A	l->1	
AF.F	ö->1	
AF.H	e->1	
AF.M	e->1	
AF:s	 ->2	
AKTU	E->1	
ANDE	 ->1	
ARPO	L->1	
AS (	I->1	
ASP 	m->1	
ATT 	O->1	
Acce	p->1	
Act.	 ->1	
Adan	a->1	
Aden	a->1	
Adol	f->2	
Adri	a->1	
Afri	k->4	
Agri	f->1	
Agus	t->1	
Aher	n->8	
Aids	,->1	
Akku	y->2	
Akkö	y->1	
Akti	v->1	
Alav	a->2	
Alba	c->1	n->1	
Albe	r->1	
Albr	i->1	
Aldr	i->1	
Alex	a->2	
Alge	r->1	
Alic	a->1	
Alla	 ->25	
Alld	e->1	
Allm	ä->4	
Allt	 ->16	f->1	s->4	
Alpe	r->1	s->1	
Alsa	c->3	
Alst	h->3	
Alte	n->18	
Amer	i->2	
Amoc	o->1	
Amok	o->5	
Amos	 ->1	
Amst	e->39	
Andr	a->7	
Ange	l->1	
Angå	e->22	
Anhå	l->1	
Anka	r->1	
Anle	d->1	
Anlä	g->1	
Anmä	l->1	
Anna	 ->1	r->4	
Anse	r->4	
Ansl	a->1	
Ansv	a->4	
Anta	l->2	
Antó	n->1	
Anve	r->1	
Anvä	n->1	
Apar	i->1	
Appl	å->5	
Arab	r->1	v->1	
Araf	a->1	
Arbe	t->4	
Arde	n->1	
Ari 	V->1	
Aria	n->3	
Arti	k->3	
Asie	n->2	
Assa	d->2	
Astu	r->1	
Atat	u->1	ü->1	
Atla	n->4	
Att 	F->1	a->1	b->1	d->4	f->1	g->3	h->2	i->2	k->1	l->2	m->2	r->1	s->1	t->2	u->3	v->1	
Atta	c->1	
Ausc	h->1	
Auto	/->1	
Auve	r->1	
Av 4	1->1	
Av a	l->4	v->1	
Av b	e->2	
Av d	e->15	
Av e	n->1	
Av o	m->1	
Av s	a->2	
Av t	r->1	
Av v	i->2	
Avbr	o->1	
Avfa	l->1	
Avgå	n->1	
Avia	n->1	
Avsa	t->1	
Avse	r->1	v->1	
Avsl	u->14	
Azor	e->2	
B Al	s->1	
B oc	h->1	
B ta	 ->1	
B-Al	s->2	
B5-0	0->4	
BATT	 ->1	
BB A	l->1	
BB-A	l->2	
BC d	e->1	
BI -	 ->1	
BNI 	b->1	i->1	o->2	p->2	
BNI,	 ->1	
BNP 	j->1	m->1	p->4	å->1	
BNP,	 ->2	
BP, 	e->1	
BRÅD	S->1	
BSE 	o->2	
BSE-	k->3	t->1	
Bako	m->2	
Balf	o->1	
Balk	a->7	
Bank	 ->1	
Bara	 ->4	k->9	
Barc	e->2	
Bare	n->1	
Barn	h->1	i->14	
Baró	n->2	
Bask	i->2	
Bass	e->1	
Bedr	ä->2	
Bedö	m->2	
Befo	r->1	
Behr	e->7	
Bekv	ä->1	
Belg	i->9	
Bene	l->1	
Bere	n->14	
Berg	 ->1	e->12	
Berl	i->7	
Bern	a->1	d->3	i->1	
Bero	e->1	
Bert	h->1	i->1	
Besl	u->4	
Besq	u->1	
Betr	ä->7	
Betä	n->25	
Bevi	s->1	
Big 	b->1	
Bili	n->1	
Bill	o->2	
Bilt	i->2	
Bisc	a->6	
Bist	å->1	
Blak	 ->1	
Blan	d->8	
Blok	 ->1	
Boet	t->1	
Bolk	e->1	
Bond	e->1	
Bord	e->4	
Bort	o->1	
Bosä	t->1	
Bour	l->6	
Bowe	.->2	
Bowi	s->2	
Bran	d->2	
Bras	i->1	
Brav	e->1	
Brem	e->1	
Bret	a->8	
Bris	t->3	
Brit	i->1	t->1	
Brok	 ->6	,->3	
Brun	o->1	
Brys	s->19	
Buda	p->1	
Budg	e->1	
Bulg	a->1	
Bush	,->1	
Busq	u->1	
Bygg	e->1	
Byrn	e->2	
Byrå	n->1	
Bäst	a->1	
Båda	 ->5	
C de	n->1	
C, a	t->1	
C-le	k->1	
C. D	e->1	
C. E	f->1	
C.Vi	 ->1	
C4-0	0->1	2->1	3->3	7->1	
C5-0	0->6	1->5	2->2	3->9	
CAF:	s->1	
CECA	F->1	
CEN 	e->1	h->1	k->1	o->1	
CEN)	 ->2	
CEN,	 ->2	
CEN:	s->4	
CERN	)->1	
CES)	 ->1	
CES-	z->3	
CH B	R->1	
CHO 	i->1	
CHO,	 ->1	
CHO.	D->1	
CK n	u->1	
CLAF	 ->1	
CM.A	t->1	
CNS)	)->9	
COD)	)->12	]->1	
COS)	]->2	
CSU-	g->1	
CSU:	s->2	
Cadi	z->5	
Cado	u->1	
Camr	e->1	
Camu	s->1	
Cana	d->1	
Cand	u->1	
Cany	o->3	
Carp	e->1	
Cart	h->1	
Casa	b->1	c->1	
Caud	r->1	
Cava	l->1	
Cent	r->13	
Cerm	i->1	
Ceyh	u->1	
Cham	p->1	
Chiq	u->1	
Clau	d->1	
Clin	t->1	
Coca	 ->1	
Coci	l->1	
Cola	,->1	
Cona	k->1	
Cons	t->1	
Corb	e->1	
Corp	u->1	
Cost	a->9	
Coun	c->1	
Cox 	o->1	s->1	
Cox!	J->1	
Cox,	 ->1	
Cres	p->2	
Cunh	a->1	
Curi	e->1	
Cusí	 ->1	
Cuxh	a->1	
Cype	r->1	
D bö	r->1	
D fö	r->1	
D kr	ä->1	
D)) 	(->2	i->2	
D))(	P->4	
D)).	.->2	F->1	
D))H	e->1	
D)].	)->1	
D, o	c->1	
D-gr	u->2	
DA) 	D->1	V->1	
DD, 	o->1	
DD-g	r->2	
DDR.	S->1	
DE F	R->1	
DE) 	H->1	J->1	Ä->1	
DE).	(->1	
DE- 	o->2	
DE-g	r->4	
DE-l	e->1	
DEBA	T->1	
DR a	n->1	
DR) 	o->1	
DR-g	r->1	
DR.S	e->1	
DR:s	 ->1	
DSKA	N->1	
Da C	o->3	
Dage	n->5	
Dagl	i->2	
Dagm	a->1	
Dala	i->7	
Dam 	b->1	s->1	
Dama	s->1	
Danm	a->26	
Darm	s->1	
Davi	d->3	
De 1	4->1	5->1	
De G	r->1	
De P	a->1	
De R	o->1	
De a	k->1	l->2	n->4	v->1	
De b	e->4	i->1	
De d	a->2	i->2	r->1	
De e	u->2	
De f	a->2	i->2	l->5	r->3	å->1	ö->9	
De g	j->1	r->8	ä->1	
De h	a->11	å->1	
De i	n->1	
De k	a->6	o->4	r->2	
De l	a->1	ö->1	
De m	i->1	y->1	å->5	
De n	o->2	u->1	y->4	ä->1	
De o	l->3	
De p	e->1	o->2	r->1	
De r	e->1	
De s	e->5	i->2	k->5	l->1	o->5	t->8	
De t	o->2	u->2	v->2	y->1	
De u	p->2	t->2	
De v	a->2	i->1	
De ä	r->4	
De å	t->2	
Delg	a->1	
Delo	r->3	
Dels	 ->1	
Delv	i->1	
Demi	n->1	
Demo	k->1	
Den 	1->2	2->2	a->22	b->4	c->1	e->15	f->24	g->10	h->17	i->5	k->14	l->2	m->10	n->7	o->7	p->3	r->7	s->25	t->11	u->2	v->8	ä->9	å->3	ö->1	
Denn	a->56	e->1	
Dera	s->2	
Dess	 ->2	a->34	u->25	
Det 	a->11	b->35	c->2	d->6	e->11	f->112	g->38	h->56	i->12	j->1	k->49	l->5	m->32	n->2	o->1	p->10	r->24	s->76	t->6	u->2	v->44	ä->361	å->4	ö->3	
Det,	 ->1	
Deta	l->1	
Dets	a->1	
Dett	a->211	
Deut	s->1	
Dimi	t->5	
Dire	k->9	
Disk	u->1	
Dock	 ->2	
Doku	m->1	
Doms	t->3	
Dori	s->1	
Dubl	i->7	
Duha	m->1	
Duis	e->3	
Dutr	o->1	
Där 	b->1	d->1	f->2	h->5	j->1	k->1	l->1	m->1	v->1	ä->1	
Dära	v->2	
Däre	f->4	m->6	
Därf	ö->96	
Däri	 ->1	g->2	
Därm	e->4	
Däru	t->1	
Därv	i->1	
Då b	ö->1	
Då d	e->1	
Då f	i->1	r->1	å->1	
Då g	i->1	
Då h	a->2	
Då k	a->3	o->4	
Då m	å->1	
Då o	c->1	
Då s	k->1	y->1	
Då t	a->1	
Då v	a->1	i->1	
Då ä	r->2	
Då ö	v->1	
Díez	 ->1	
Dühr	k->1	
E FR	Å->1	
E ha	r->2	
E oc	h->2	
E ti	l->1	
E är	 ->1	
E) H	e->1	
E) J	a->1	
E) Ä	r->1	
E).(	E->1	
E)Ja	g->1	
E- o	c->2	
E-DE	)->1	-->7	
E-gr	u->12	
E-ko	l->1	
E-kr	i->3	
E-le	d->1	
E-te	s->1	
E/NG	L->2	
EBAT	T->1	
ECAF	:->1	
ECHO	 ->1	,->1	.->1	
EDD,	 ->1	
EDD-	g->2	
EEG 	t->1	
EEG,	 ->2	
EG a	t->1	
EG o	m->2	
EG s	k->1	
EG t	i->2	
EG u	p->1	
EG, 	E->4	f->1	o->1	v->1	
EG-d	i->2	o->22	
EG-f	ö->8	
EG-i	n->1	
EG-k	o->16	
EG-r	ä->3	
EG.V	i->1	
EG:s	 ->3	
EG?,	 ->1	
EIF 	h->1	
EIF)	,->1	
EK (	d->1	
EK(1	9->3	
EK(9	9->1	
EKSG	,->2	-->6	
EL) 	F->1	H->1	J->1	
ELDR	 ->1	-->1	:->1	
ELLA	 ->1	
EM-2	0->1	
EMU,	 ->1	
EMU-	a->1	k->1	
EMU:	s->3	
EN e	l->1	
EN h	a->1	
EN k	o->1	
EN o	c->1	
EN) 	D->2	F->6	H->4	I->3	J->7	K->1	L->2	M->1	S->1	T->4	U->1	V->2	i->1	s->1	
EN, 	a->1	s->1	
EN-g	r->1	
EN:s	 ->4	
EO b	e->2	
EO ä	r->1	
EP (	"->1	
EP r	e->1	
ERN)	 ->1	
ERRE	G->3	
ES) 	-->1	ä->1	
ES-z	o->3	
EU "	c->1	
EU I	 ->1	
EU a	g->1	t->2	
EU b	l->1	ö->1	
EU d	ä->1	
EU f	r->1	
EU g	e->1	ö->1	
EU h	a->2	
EU i	 ->1	n->3	
EU k	a->3	
EU m	e->1	y->1	å->1	
EU o	c->4	
EU p	å->1	
EU r	e->1	
EU s	k->1	o->4	y->1	
EU u	t->2	
EU ä	r->2	
EU, 	f->1	l->1	m->1	p->1	v->1	
EU-b	i->1	u->1	
EU-e	n->1	
EU-f	o->1	ö->5	
EU-g	e->1	
EU-i	n->5	
EU-k	o->6	
EU-l	a->2	ä->3	
EU-m	a->1	e->5	
EU-n	i->1	
EU-o	r->1	
EU-p	r->2	
EU-r	e->1	ä->1	
EU-s	t->1	ä->2	
EU-t	e->1	
EU-u	t->1	
EU-v	ä->1	
EU..	 ->1	
EU.A	l->1	
EU.D	a->1	e->2	
EU.F	r->1	
EU.N	u->1	
EU.R	o->1	
EU.V	i->3	
EU:s	 ->44	
EU?H	e->1	
EUGF	J->3	
Ecem	i->1	
Edin	b->1	
Effe	k->5	
Efta	r->2	
Efte	r->48	
Egyp	t->2	
Ehud	 ->2	
Eiec	k->1	
Ekof	i->2	
Ekon	o->3	
Elis	a->1	
Elle	r->1	s->3	
Elma	r->2	
Elst	.->1	
Emel	l->8	
Emil	i->1	
En a	l->3	n->6	s->1	v->6	
En b	e->1	o->2	ä->1	
En d	e->7	
En f	r->2	ö->2	
En g	e->1	
En k	a->1	n->1	o->3	
En m	a->1	e->1	
En p	e->1	r->1	
En r	a->2	e->2	
En s	a->1	i->1	u->1	y->1	ä->1	å->4	
En u	p->1	
En v	a->1	e->1	i->4	ä->4	
En ö	k->1	v->1	
Enba	r->1	
Enda	s->11	
Enke	l->1	
Enli	g->37	
Equa	l->8	
Equq	a->2	
Er a	n->1	
Era 	t->1	
Erfa	r->2	
Erik	a->29	
Erit	r->1	
Erkk	i->2	
Ert 	b->1	p->1	
Etio	p->3	
Ett 	E->1	a->11	d->2	e->5	f->4	h->1	l->1	m->1	n->3	o->2	p->1	s->10	t->2	v->3	å->1	
Eura	t->4	
Euro	-->1	d->5	j->6	n->1	p->832	s->2	
Evan	s->7	
Even	t->1	
Exce	p->1	
Exem	p->1	
Expe	r->2	
Exup	é->1	
Exxo	n->3	
F gö	r->1	
F ha	r->1	
F i 	e->1	r->1	
F ka	n->1	
F ko	n->1	
F sk	a->1	
F) ä	r->1	
F), 	b->1	
F, E	u->1	
F, d	e->1	
F, e	n->1	
F, k	o->1	
F, s	å->2	
F, v	i->1	
F, ö	v->1	
F.Al	l->1	
F.Fö	r->1	
F.He	r->1	
F.Me	n->1	
F:s 	(->1	u->1	
FAF,	 ->1	
FBI 	-->1	
FEO 	b->2	ä->1	
FI) 	J->1	
FIL,	 ->1	
FIPO	L->1	
FJ) 	f->1	
FJ),	 ->1	
FJ:s	 ->1	
FMI 	d->1	
FN, 	s->1	
FN-u	p->1	
FN.H	e->1	
FN:s	 ->8	
FOP)	.->1	
FPÖ 	(->2	f->1	h->1	i->1	m->1	o->3	s->1	v->1	ä->1	
FPÖ)	.->1	
FPÖ-	l->1	m->1	
FPÖ:	s->4	
FR) 	"->1	D->4	E->1	F->1	H->1	I->2	J->4	N->3	T->1	
FRÅG	O->1	
FSR 	-->1	
FUF)	 ->1	
Fack	f->3	
Fact	o->1	
Fakt	u->4	
Farl	i->1	
Faro	u->1	
Fasc	i->1	
Feir	a->2	
Fela	k->1	
Fem 	l->1	
Fina	 ->3	.->1	n->2	
Finl	a->6	
Finn	s->4	
Firm	a->1	
Fisc	h->4	
Flau	t->2	
Fler	a->3	t->1	
Flor	e->19	
Fléc	h->1	
FoU,	 ->1	
FoU-	r->1	
Fog 	f->1	
Folk	 ->3	f->1	r->2	
Font	a->1	
Ford	,->1	
Fore	s->1	
Fors	k->2	
Frag	a->1	
Fram	 ->1	f->2	l->1	s->2	t->2	å->1	
Fran	c->3	k->39	o->1	s->2	z->3	ç->1	
Fras	s->1	
Fred	s->1	
Frih	e->3	
Fru 	A->1	B->1	L->1	M->1	P->1	S->1	k->4	l->2	t->70	
Frut	e->3	
Främ	j->1	s->1	
Fråg	a->37	e->2	o->3	
Från	 ->2	
Fund	 ->1	
Fyrt	i->1	
Fäst	n->1	
Får 	j->3	
Följ	a->5	d->1	
För 	1->2	a->31	b->1	d->100	e->4	f->2	i->1	k->1	l->1	m->9	n->8	o->6	p->1	s->3	t->4	u->1	v->7	å->1	ö->3	
Förb	u->5	
Förd	e->1	r->2	
Före	b->1	d->8	n->44	t->2	
Förf	a->1	
Förh	i->1	o->3	
Föri	n->2	
Förl	u->1	
Förm	o->1	
Föro	r->1	
Förp	a->1	
Förs	i->1	l->8	t->28	ä->1	ö->1	
Fört	j->1	r->1	
Föru	t->7	
Förv	a->1	i->2	ä->1	
Förä	n->1	
G at	t->1	
G om	 ->2	
G sk	u->1	
G ti	l->2	
G up	p->1	
G(Pa	r->1	
G, E	E->2	u->4	
G, f	ö->1	
G, o	m->1	
G, v	i->1	
G-di	r->2	
G-do	m->22	
G-fö	r->14	
G-in	i->1	
G-ko	r->16	
G-rä	t->3	
G.(E	N->1	
G.Vi	 ->1	
G:s 	d->1	l->1	m->1	
G?, 	r->1	
GA-s	t->1	
GASP	 ->1	
GFJ)	 ->1	,->1	
GFJ:	s->1	
GL-g	r->2	
GORN	ä->1	
GUE/	N->2	
GUSP	 ->1	
Gale	o->1	
Gali	c->2	
Gama	 ->3	
Garg	a->5	
Gaza	 ->1	,->1	.->2	r->2	
Geme	l->1	n->5	
Gene	r->10	
Geno	m->28	
Genè	v->3	
Ger 	d->1	
Gil-	D->1	R->1	
Gino	,->1	
Give	t->2	
Goeb	b->1	
Gola	n->9	
Golf	s->3	
Goll	n->1	
Gome	s->1	
Gonz	á->1	
Good	w->1	
Gors	e->1	
Gott	 ->1	
Grac	a->3	o->1	
Grat	u->1	
Graç	a->5	
Grek	l->14	
Gros	s->3	
Grun	d->1	
Grup	p->10	
Grön	a->1	i->1	
Guat	e->1	
Guig	o->1	
Gulf	k->1	
Gusp	"->1	
Gute	r->2	
Gäll	a->1	
Gå h	e->1	
Gör 	v->2	
Göte	b->1	
H BR	Å->1	
H-00	0->1	
H-07	7->1	8->6	9->5	
H-08	0->4	1->3	2->1	
HO i	 ->1	
HO, 	a->1	
HO.D	e->1	
Haar	d->1	
Hade	 ->2	r->1	
Hagu	e->1	
Haid	e->37	
Hamb	u->1	
Han 	a->1	b->1	h->7	k->1	n->1	s->3	t->1	ä->3	
Hand	e->1	i->1	l->2	
Hans	 ->3	
Har 	k->3	m->2	o->1	r->2	v->3	
Harr	i->1	
Hatz	i->2	
Have	n->1	
Heat	o->1	
Hebr	o->1	
Hedg	e->1	
Hedk	v->1	
Hein	z->2	
Hela	 ->3	
Heli	g->1	
Hels	i->20	
Helt	 ->2	
Heml	i->1	
Henr	y->1	
Herr	 ->329	
Hick	s->1	
Hilt	o->1	
Hima	l->1	
Hist	o->2	
Hit 	h->3	
Hitl	e->6	
Hitt	i->3	
Holl	y->1	
Holz	m->2	
Hon 	h->2	l->1	s->1	
Hopp	e->1	
Howi	t->1	
Huhn	e->1	
Hult	e->19	h->6	
Hur 	b->1	f->2	g->1	h->1	k->3	l->2	m->4	s->19	t->1	ä->1	
Huru	v->1	
Huvu	d->7	
Hyck	l->1	
Händ	e->2	
Häns	c->2	
Här 	b->5	f->3	g->1	h->4	i->1	k->5	m->2	n->1	r->2	s->1	t->3	v->3	ä->2	
Härm	e->2	
Häro	m->1	
Håll	e->1	
Höge	r->1	
I - 	K->1	P->1	R->1	d->1	
I Am	s->1	
I Eu	r->4	
I Fr	a->2	
I He	l->1	
I Ir	l->2	
I It	a->1	
I Ne	d->1	
I Ra	p->1	
I Sc	h->1	
I Ti	b->1	
I Tu	r->1	
I Ty	s->1	
I al	l->3	
I an	d->1	n->2	
I ap	r->1	
I ar	t->1	
I av	s->1	v->2	
I be	t->6	
I bu	d->1	
I bö	r->2	
I da	g->24	
I de	 ->2	n->23	t->35	
I di	r->1	
I dä	r->1	
I eg	e->7	
I en	 ->7	l->4	
I er	a->1	
I et	t->2	
I fj	o->1	
I fl	e->1	
I fo	r->1	
I fr	a->1	å->5	
I fö	r->6	
I gå	r->3	
I ha	r->2	
I i 	E->1	a->1	f->1	
I ju	n->1	
I kl	a->1	
I ko	m->2	n->1	
I kr	i->1	
I li	k->7	
I me	d->1	
I mi	n->1	t->1	
I mo	r->3	t->3	
I må	l->1	
I no	v->2	
I nä	s->2	
I oc	h->8	
I ok	t->1	
I pa	r->1	
I pe	r->2	
I pr	i->1	o->1	
I ra	p->2	
I re	a->1	g->1	s->5	v->1	
I rä	t->1	
I rå	d->1	
I sa	m->3	
I si	n->1	t->2	
I sj	ä->4	
I sk	a->1	
I sl	u->3	
I st	i->1	r->1	ä->9	
I sy	n->1	s->1	
I så	 ->3	d->1	
I tj	u->1	
I up	p->1	
I ut	b->1	s->1	
I va	r->2	
I ve	r->1	
I vi	l->3	s->2	t->2	
I vo	n->1	
I vä	n->2	
I vå	r->6	
I än	d->1	
I öv	r->3	
I) J	a->1	
I) o	c->1	
I); 	e->1	
I, e	t->1	
I, h	a->1	
I-pr	o->3	
I. f	ö->2	
I:e 	r->2	
ICES	)->1	-->3	
IF h	a->1	
IF),	 ->1	
IFIL	,->1	
IFOP	)->1	
II -	 ->2	
II h	a->2	
II i	 ->1	
II k	r->1	
II s	k->1	
II) 	o->1	
II, 	h->1	
II-p	r->2	
II. 	f->1	
II:e	 ->2	
III 	-->1	h->1	k->1	s->1	
III:	e->1	
IK, 	v->1	
IK.D	e->2	
IL, 	f->1	
IMO)	.->1	
IMO.	D->1	
IMO:	s->1	
INA 	h->1	v->1	
INA,	 ->1	
ING(	P->1	
ING.	(->1	
INTE	 ->1	R->3	
IPOL	)->1	
IRA 	h->1	
ISPA	-->1	
IT) 	D->1	H->1	O->1	
IV -	 ->1	
IV i	 ->2	
IX o	c->1	
IX, 	f->1	
Ibla	n->3	
Idén	 ->1	
Ihål	l->1	
Ile-	d->1	
Ille	g->1	
Imbe	n->3	
Immi	g->1	
Indi	e->5	
Indu	s->1	
Infö	r->4	
Inga	 ->2	
Inge	n->10	r->1	t->3	
Ingl	e->2	
Init	i->3	
Inne	b->1	h->1	
Inom	 ->10	
Inre	 ->1	s->1	
Inrä	t->1	
Insa	t->2	
Inte	 ->15	r->21	
Irla	n->22	
Isab	e->2	
Isla	n->1	
Isra	e->38	
Ista	n->1	
Ital	i->18	
Izqu	i->1	
J) f	i->1	
J), 	ä->1	
J:s 	g->1	
Ja E	r->1	
Ja e	l->1	
Ja t	i->1	
Ja, 	d->1	f->1	h->2	j->1	n->1	s->1	v->1	
Jack	s->2	
Jaco	b->2	
Jacq	u->3	
Jag 	a->64	b->34	d->8	e->1	f->48	g->13	h->98	i->9	j->1	k->50	l->3	m->26	n->4	o->1	p->5	r->14	s->131	t->133	u->31	v->212	ä->56	ö->11	
Jan-	K->1	
Japa	n->3	
Jave	t->1	
Jean	-->1	
Jeru	s->2	
Jo d	å->1	
Jo, 	d->1	i->1	s->1	
Jona	s->2	
Jonc	k->14	
Jord	a->2	b->2	
Josp	i->1	
Ju m	i->1	
Jugo	s->1	
Junk	e->1	
Just	 ->8	e->2	
Jämf	ö->2	
Jäms	t->1	
Jörg	 ->14	
Jørg	e->2	
K (d	e->1	
K nu	 ->1	
K(19	9->3	
K(99	)->1	
K, d	e->1	
K, v	i->1	
K.De	t->2	
KAND	E->1	
KOM(	1->8	9->2	
KSG,	 ->2	
KSG-	f->6	
KTUE	L->1	
Kafo	r->1	
Kale	i->2	j->1	
Kan 	k->5	m->1	n->4	r->1	u->1	v->1	
Kana	d->1	
Kans	k->9	
Kant	a->3	
Kara	s->3	
Karl	 ->4	-->1	s->2	
Kart	e->2	
Kasp	i->1	
Kata	s->1	
Kauf	m->1	
Kauk	a->3	
Kaza	k->1	
Kees	 ->1	
Kfor	 ->1	
Kina	 ->7	,->1	.->1	s->1	
Kinn	o->24	
Kirg	i->5	
Knap	p->1	
Koch	 ->6	)->1	,->5	.->1	I->1	s->1	
Kode	n->1	
Koll	e->1	
Kom 	i->1	
Komm	e->12	i->107	u->1	
Komp	r->1	
Konk	r->1	u->13	
Konr	a->1	
Kons	e->1	t->1	u->3	
Konv	e->2	
Kore	a->2	
Kort	 ->2	
Koso	v->60	
Kost	n->4	
Kouc	h->12	
Krav	 ->1	e->2	
Kult	u->25	
Kuma	r->1	
Kung	l->1	
Kvan	t->1	
Kvin	n->5	
Kväk	a->1	
Kyot	o->7	
Känn	e->1	
Kära	 ->6	
Kärn	a->1	k->2	t->1	
Köln	 ->2	
Köpe	n->1	
L (e	n->1	
L) A	t->1	
L) F	P->1	
L) H	e->4	
L) J	a->1	
L), 	m->1	
L, f	i->1	
L-gr	u->2	
LA O	C->1	
LAF 	g->1	i->2	k->2	s->1	
LAF,	 ->7	
LAF.	A->1	F->1	H->1	M->1	
LAF:	s->1	
LAS 	(->1	
LDR 	a->1	
LDR-	g->1	
LDR:	s->1	
LFAF	,->1	
LLA 	O->1	
LTCM	.->1	
La R	é->2	
Laan	 ->1	.->1	s->5	
Lama	 ->3	.->2	s->2	
Land	i->1	s->1	
Lang	e->30	
Lank	a->3	
Lapp	l->2	
Le B	e->1	
Lead	e->5	
Leda	m->4	
Ledn	i->1	
Lein	e->6	s->2	
Leon	i->1	
Liba	n->5	
Libe	r->2	
Liby	e->1	
Liik	a->3	
Lika	 ->1	s->2	
Likr	i->1	
Liks	o->8	
Likv	ä->1	
Lill	e->1	
Liss	a->8	
Lita	u->1	
Litt	e->1	
Livl	i->2	
Livs	m->3	
Lloy	d->1	
Loir	e->3	
Lomé	a->1	k->1	
Lond	o->4	
Lord	 ->2	
Lorr	a->2	
Loth	a->3	
Lous	e->1	
Loyo	l->2	
Lutt	e->1	
Luxe	m->6	
Lyck	a->1	l->1	
Lynn	e->4	
Lägg	 ->2	
Länd	e->1	
Lån 	a->1	
Lång	r->1	
Låt 	e->1	i->1	m->40	o->18	v->1	
Lööw	 ->1	
M AK	T->1	
M so	m->1	
M(19	9->8	
M(98	)->1	
M(99	)->1	
M-20	0->1	
M.At	t->1	
MARP	O->1	
MI d	ä->1	
MIK,	 ->1	
MIK.	D->2	
MO).	F->1	
MO.D	e->1	
MO:s	 ->1	
MRÖS	T->2	
MU, 	t->1	
MU-a	n->1	
MU-k	r->1	
MU:s	 ->3	
Maas	t->6	
Maca	o->1	
Mada	g->1	
Made	i->2	
Madr	i->3	
Main	s->1	
Majo	r->1	
Malt	a->7	
Man 	b->8	f->3	g->2	h->4	i->1	j->1	k->12	l->1	m->14	r->1	s->3	t->2	u->3	v->1	
Mann	e->2	
Marg	a->1	o->1	
Mari	a->1	e->1	n->6	
Mark	n->4	o->1	
Marp	o->1	
Mars	e->1	
Mart	i->1	
Math	i->2	
Maxi	m->2	
McCa	r->1	
McNa	l->5	
Med 	a->3	d->12	e->2	f->1	h->6	o->2	s->2	t->7	
Meda	n->4	
Medb	e->1	o->2	
Mede	l->3	
Medg	e->1	
Medl	e->9	
Mell	a->20	
Men 	-->2	C->1	E->1	F->1	a->5	b->2	d->55	e->6	f->7	g->1	h->7	i->9	j->33	k->5	m->4	n->5	o->4	p->5	s->13	t->3	u->4	v->32	ä->3	å->1	
Men,	 ->3	
Mena	r->1	
Ment	a->1	
Mer 	s->1	v->1	ä->1	
Mexi	k->1	
Mich	i->1	
Midd	e->1	
Midl	a->1	
Milj	ö->1	
Min 	a->6	d->1	f->5	g->9	k->1	p->1	s->4	t->2	u->1	å->1	ö->1	
Mina	 ->18	
Mind	r->1	
Mini	s->1	
Minn	s->1	
Mins	k->1	
Minu	c->1	
Mist	e->2	
Mitr	o->1	
Mitt	 ->3	e->2	
Mont	i->17	r->2	
Mora	l->1	t->4	
Morb	i->1	
Morg	a->4	
Mosk	v->1	
Mot 	b->4	d->4	
Mour	a->8	
Mous	k->1	
Muld	e->1	
Myck	e->1	
Myll	e->1	
Mynd	i->3	
Männ	i->5	
Märk	l->1	
Måhä	n->1	
Måle	t->2	
Mång	a->10	
Möjl	i->2	
Münc	h->1	
N el	l->1	
N ha	r->1	
N ko	m->1	
N oc	h->1	
N) D	e->2	
N) F	r->4	å->1	ö->1	
N) H	e->4	
N) I	 ->3	
N) J	a->7	
N) K	o->1	
N) L	å->2	
N) M	i->1	
N) S	e->1	
N) T	a->3	i->1	
N) U	n->1	
N) V	a->2	
N) i	 ->1	n->1	
N) s	o->1	
N)).	 ->1	
N, a	l->1	
N, s	o->2	
N-gr	u->1	
N-up	p->1	
N.He	r->1	
N:s 	a->3	b->2	e->1	g->1	r->1	s->3	v->1	
NA h	a->1	
NA v	a->1	
NA, 	e->1	
NDE 	F->1	
NG(P	a->1	
NG.(	E->1	
NGL-	g->2	
NI b	e->1	
NI i	 ->1	
NI o	c->2	
NI p	e->2	
NI, 	e->1	
NIFI	L->1	
NING	(->1	.->1	
NL) 	A->1	H->3	
NMIK	,->1	.->2	
NP j	ä->1	
NP m	i->1	
NP p	e->3	å->1	
NP å	r->1	
NP, 	i->1	m->1	
NS))	 ->1	(->4	.->2	F->1	o->1	
NTE 	h->1	
NTER	R->3	
Nall	y->5	
Nana	 ->1	
Napo	l->1	
Nark	o->1	
Nati	o->7	
Nato	 ->1	a->1	b->1	s->2	
Natu	r->15	
Nede	r->9	
Nej,	 ->7	
Nej.	I->1	
New 	Y->1	
Ni a	g->1	
Ni b	e->3	o->1	
Ni f	r->1	ö->2	
Ni h	a->11	
Ni k	a->2	o->5	ä->2	
Ni l	ä->1	
Ni m	å->4	
Ni n	ä->1	
Ni s	a->3	k->2	ä->1	
Ni t	a->2	
Ni v	e->2	i->1	
Niel	s->6	
Niki	t->2	
Nivå	n->1	
Nogu	e->1	
Noir	m->1	
Nord	i->3	
Norg	e->2	
Norm	a->1	e->1	
Nu a	n->2	
Nu b	e->1	
Nu f	i->1	å->1	ö->1	
Nu h	a->6	o->1	
Nu k	a->2	
Nu m	å->1	
Nu t	i->1	
Nu v	e->1	ä->1	
Nu ä	r->7	
Nu å	t->1	
Nume	r->1	
Nuva	r->1	
Nya 	Z->2	r->1	
Nyli	g->1	
Nytt	 ->1	
När 	a->3	b->2	d->35	e->1	f->1	j->7	k->6	m->7	n->1	p->1	s->1	t->2	v->16	
Näst	a->26	
Någo	n->2	t->1	
Någr	a->2	
Nåja	,->1	
Nödv	ä->1	
O be	f->1	s->1	
O i 	b->1	
O är	 ->1	
O).F	ö->1	
O, a	k->1	
O.De	t->2	
O:s 	n->1	
O?En	d->1	
OCH 	B->1	
OD))	 ->4	(->4	.->3	H->1	
OD)]	.->1	
OFSR	 ->1	
OK, 	d->1	
OL (	e->1	
OL),	 ->1	
OLAF	 ->5	,->7	.->4	:->1	
OLAS	 ->1	
OLFA	F->1	
OM A	K->1	
OM(1	9->8	
OM(9	8->1	9->1	
OMRÖ	S->2	
OP).	V->1	
ORNä	s->1	
OS)]	.->2	
OSSE	 ->1	
Oavs	e->2	
Ober	b->1	o->2	
Och 	E->1	S->1	a->2	d->21	e->2	g->1	h->1	i->2	j->10	k->1	m->1	n->5	o->2	s->7	t->1	v->8	ä->1	
Och:	 ->1	
Ocks	å->2	
Offe	n->3	
Offi	c->1	
Ofta	 ->1	
Oil 	P->1	
Oil-	p->1	
Olik	a->1	
Oliv	i->1	
Olje	b->2	t->1	
Olym	p->1	
Om 5	0->1	
Om E	U->1	u->1	
Om S	c->1	y->1	
Om a	l->3	
Om b	e->1	
Om d	e->21	o->1	u->1	
Om e	n->2	r->1	t->2	
Om f	o->1	
Om g	e->1	i->1	
Om i	n->4	
Om j	a->2	
Om k	a->1	o->4	
Om l	a->1	
Om m	a->11	
Om n	i->7	å->1	
Om o	m->1	
Om p	a->2	
Om r	e->1	å->1	
Om s	l->1	y->1	
Om t	r->1	v->1	
Om u	p->1	
Om v	i->23	
Omag	h->1	
Omrö	s->15	
Ones	t->1	
Onöd	i->1	
Oran	i->1	
Ord 	s->1	
Orde	n->1	r->1	t->1	
Ordf	ö->7	
Orka	n->2	
Oron	 ->1	
Orov	ä->1	
Orsa	k->2	
Oslo	 ->1	,->2	
Osma	n->1	
Ouvr	i->1	
Oz d	y->1	
Oz h	a->1	
Oz, 	b->1	
P ("	d->1	
P (Ö	s->2	
P at	t->2	
P jä	m->1	
P mi	n->1	s->1	
P må	s->1	
P oc	h->1	
P pe	r->3	
P på	 ->1	
P re	p->1	
P år	 ->1	
P) o	c->1	
P).V	i->1	
P, e	f->1	
P, i	 ->1	
P, m	e->1	
PA-i	n->1	
PE h	a->1	
PE ä	r->1	
PE-D	E->8	
PE-g	r->5	
PM s	o->1	
POL 	(->1	
POL)	,->1	
PPE 	h->1	ä->1	
PPE-	D->8	g->5	
PR-e	f->1	
PSE)	J->1	
PSE-	g->3	
PT) 	E->1	F->1	H->9	J->2	L->1	N->1	V->1	
PVC,	 ->1	
PVC-	l->1	
PVC.	V->1	
Pack	 ->2	s->1	
Padd	i->2	
Paki	s->5	
Pala	c->15	
Pale	r->1	s->10	
Papa	y->2	
Para	g->1	
Pari	s->3	
Parl	a->42	
Patt	e->23	
Pays	 ->1	-->1	
Peak	e->1	
Peij	s->2	
Peki	n->1	
Pers	o->4	
Pete	r->1	
Petr	o->1	
Plan	e->1	t->1	
Plas	t->2	
Plat	h->4	o->1	
Ploo	i->1	
Pläd	e->1	
Poet	t->5	
Pohj	a->1	
Pole	n->1	
Poll	u->1	
Pomé	s->1	
Ponn	a->1	
Poos	 ->1	
Port	u->27	
Powe	r->3	
Prec	i->6	
Pres	e->1	
Preu	s->1	
Prio	r->1	
Prob	l->9	
Proc	e->3	
Prod	i->28	u->2	
Prog	r->1	
Proj	e->2	
Prot	o->2	
Prov	a->3	
Prín	c->1	
Punk	t->2	
Purv	i->1	
PÖ (	Ö->2	
PÖ f	ö->1	
PÖ h	ä->1	
PÖ i	n->1	
PÖ m	i->1	
PÖ o	c->3	m->1	
PÖ s	o->1	
PÖ v	i->1	
PÖ ä	r->1	
PÖ) 	s->1	
PÖ).	J->1	
PÖ-l	e->1	
PÖ-m	e->1	
PÖ:s	 ->4	
På a	l->1	
På d	e->22	
På e	t->1	
På g	r->2	
På l	a->1	
På m	a->1	i->1	å->1	
På o	m->2	
På p	a->1	
På s	a->4	i->3	å->4	
På u	p->1	
På v	i->3	
Påst	å->1	
Péta	i->1	
Quec	e->1	
R - 	o->1	
R an	s->1	
R) "	T->1	
R) D	e->4	
R) E	f->1	
R) F	r->1	
R) H	e->1	
R) I	 ->2	
R) J	a->3	ö->1	
R) N	e->1	ä->2	
R) T	h->1	
R) o	c->1	
R-ef	f->1	
R-gr	u->1	
R.Se	d->1	
R:s 	u->1	
RA h	a->1	
REG,	 ->1	
REG-	i->1	
REG?	,->1	
REP 	(->1	r->1	
RINA	 ->2	,->1	
RN) 	i->1	
RNäs	t->1	
RPOL	 ->1	
RREG	,->1	-->1	?->1	
Rack	 ->1	,->1	
Rafa	e->3	
Rand	z->4	
Rapk	a->11	
Rapp	o->3	
Rasc	h->1	
Rasi	s->1	
Read	i->1	
Reak	t->1	
Reda	n->3	
Redi	n->8	
Refo	r->7	
Rege	r->6	
Regi	o->1	
Rent	 ->2	
Repu	b->1	
Rest	e->2	
Resu	l->5	
Retr	o->1	
Revi	d->1	s->3	
Rhôn	e->1	
Rich	a->1	t->2	
Riis	-->2	
Rika	 ->1	
Rikt	l->4	
Riof	ö->1	
Risk	e->1	
Robe	r->1	
Robl	e->1	
Rois	s->1	
Rojo	s->1	
Rom-	 ->1	
Roma	g->1	n->2	
Romá	n->1	
Roo 	f->1	
Rope	t->1	
Roth	-->7	
Rott	e->2	
Rove	r->2	
Roya	l->1	
Ruiz	 ->1	
Rumä	n->1	
Rush	 ->1	
Ryss	l->4	
RÅDS	K->1	
RÅGO	R->1	
RÖST	N->2	
Räkn	a->1	
Rätt	s->2	
Råde	r->1	t->20	
Råds	o->1	
Réun	i->2	
Röst	a->1	
S (I	n->1	
S oc	h->1	
S) -	 ->1	
S) ä	r->1	
S)) 	(->1	
S))(	G->1	P->3	
S)).	.->1	J->1	
S))F	r->1	
S))o	c->1	
S)].	H->2	
S-zo	n->3	
S:s 	p->1	
SA -	 ->1	
SA a	t->1	
SA e	l->1	
SA h	a->1	
SA p	å->1	
SA, 	K->1	s->1	
SA.J	a->1	
SA.V	i->1	
SA:s	.->1	
SD f	ö->1	
SE o	c->2	
SE t	i->1	
SE)J	a->1	
SE-g	r->3	
SE-k	r->3	
SE-t	e->1	
SEK 	(->1	
SEK(	1->3	9->1	
SEM-	2->1	
SG, 	E->2	
SG-f	ö->6	
SKAN	D->1	
SOLA	S->1	
SP m	å->1	
SP o	c->1	
SPA-	i->1	
SPÖ 	o->1	
SPÖ)	 ->1	
SR -	 ->1	
SS o	c->1	
SS:s	 ->1	
SSE 	t->1	
STNI	N->2	
SU-g	r->1	
SU:s	 ->2	
SYN)	)->1	
Sage	s->1	
Sain	t->1	
Sala	f->1	
Samh	ä->2	
Samm	a->26	
Samo	r->1	
Samt	i->14	
San 	S->1	
Sann	i->5	o->1	
Sant	a->1	e->2	
Save	 ->4	,->1	-->3	N->1	
Sche	n->10	
Schr	e->3	o->14	ö->1	
Schu	l->3	
Schw	a->1	e->1	
Schö	r->1	
Schü	s->4	
Seat	t->4	
Seba	s->1	
Seda	n->20	
Segn	i->1	
Segu	r->1	
Seix	a->5	
Seri	ö->1	
Sett	 ->1	
Shar	a->1	m->5	
Shei	k->5	
Shel	l->2	
Shep	h->3	
Simp	s->1	
Sist	 ->2	
Situ	a->3	
Sju 	ä->1	
Sjuk	h->1	
Själ	v->2	
Sjät	t->1	
Sjös	t->4	
Skad	o->1	
Skal	l->4	
Skog	s->1	
Skot	t->5	
Skul	l->8	
Skyd	d->1	
Skäl	e->1	
Slov	a->1	
Slut	l->34	r->1	s->3	
Små 	o->1	
Småf	ö->1	
Snab	b->1	
Snar	a->1	
Soar	e->1	
Soci	a->4	
Sokr	a->1	
Sola	n->4	
Solb	e->2	
Som 	E->1	T->1	a->2	b->1	e->9	f->3	h->1	j->8	k->3	l->2	m->1	n->9	p->3	s->4	t->1	u->1	v->3	
Soml	i->3	
Soul	a->1	
Span	i->7	
Spen	c->1	
Sper	o->1	
Sri 	L->3	
St.V	a->1	
Stab	i->1	
Stad	g->1	
Stat	e->6	i->1	l->2	
Stoc	k->3	
Stor	a->2	b->14	m->2	
Stra	f->1	s->5	x->1	
Stru	k->1	
Strä	v->1	
Stäm	m->1	
Stål	s->1	
Stöd	 ->3	e->3	s->1	
Stör	r->2	s->2	
Suan	z->1	
Subv	e->2	
Sudr	e->2	
Svar	e->1	
Svep	e->1	
Sver	i->7	
Swob	o->3	
Syda	f->2	
Sydk	o->1	
Sydo	s->2	
Syft	e->6	
Syri	e->24	
Sánc	h->1	
São 	T->2	
Säg 	m->1	
Säke	r->2	
Särs	k->2	
Så b	l->1	
Så d	e->3	
Så e	n->1	r->1	
Så f	r->1	
Så h	ä->1	
Så j	a->3	
Så k	a->1	o->1	
Så l	ä->3	å->2	
Så n	å->1	
Så r	i->1	
Så s	e->1	o->2	ä->1	
Så t	i->1	
Så v	a->1	i->4	å->1	
Så ä	r->1	v->2	
Såda	n->2	
Såle	d->4	
Sång	e->1	
Såso	m->2	
Såvä	l->1	
Söde	r->2	
T OM	 ->1	
T) D	e->1	
T) E	f->1	
T) F	r->1	
T) H	e->10	
T) J	a->2	
T) L	e->1	
T) N	ä->1	
T) O	m->1	
T) V	i->1	
TCM.	A->1	
TE h	a->1	
TERR	E->3	
TNIN	G->2	
TO?E	n->1	
TT O	M->1	
TUEL	L->1	
TV a	n->1	
TV-b	i->1	
TV-k	a->1	
TV-p	r->1	
TV-s	ä->1	
Ta d	ä->1	
Taci	s->2	
Tack	 ->24	,->13	.->1	
Tadz	j->5	
Taiw	a->1	
Tala	r->1	
Talm	a->9	
Tamm	e->22	
Tang	 ->1	
Tani	o->1	
Tank	e->3	
Taue	r->1	
Terr	o->1	ó->3	
Tesa	u->1	
Texa	s->2	
Thea	t->21	
Thys	s->5	
Tibe	t->21	
Tidi	g->1	
Tidn	i->1	
Till	 ->31	s->2	v->3	ä->3	å->10	
Titt	a->1	
Todi	n->1	
Tom 	S->1	
Tomé	 ->2	
Tong	i->1	
Topp	m->2	
Torr	e->3	
Torv	 ->1	e->1	
Tota	l->6	
Tran	s->3	
Tre 	ä->1	
Tred	j->1	
Trit	t->1	
Tror	 ->2	
Trot	s->17	
Trov	ä->1	
Träd	 ->1	
Tsat	s->3	
Turk	i->35	m->2	
Tuse	n->1	
Tvär	t->4	
Två 	v->1	ä->1	
Ty e	n->1	
Ty h	a->1	
Ty i	n->1	
Ty s	o->1	
Ty u	n->1	
Ty v	a->1	i->2	
Tyck	e->1	
Tydl	i->1	
Tysk	l->20	
Tyvä	r->9	
Tänk	 ->2	
Tågk	r->1	
U "c	o->1	
U I 	e->1	
U ag	e->1	
U at	t->2	
U bl	a->1	
U bö	r->1	
U dä	r->1	
U fr	a->1	
U ge	r->1	
U gö	r->1	
U ha	r->2	
U i 	d->1	
U in	f->2	t->1	
U ka	n->3	
U me	r->1	
U my	c->1	
U må	s->1	
U oc	h->4	
U på	 ->1	
U re	d->1	
U sk	a->1	
U so	m->4	
U sy	s->1	
U ut	s->1	v->1	
U är	 ->2	
U, f	ö->1	
U, l	å->1	
U, m	e->1	
U, n	ä->1	
U, p	å->1	
U, t	y->1	
U, v	i->1	
U-an	p->1	
U-bi	s->1	
U-bu	d->1	
U-en	h->1	
U-fo	n->1	
U-fö	r->5	
U-ge	n->1	
U-gr	u->1	
U-in	i->1	s->4	
U-ko	m->2	r->4	
U-kr	i->1	
U-la	g->1	n->1	
U-lä	n->3	
U-ma	n->1	
U-me	d->5	
U-ni	v->1	
U-or	d->1	
U-pr	o->2	
U-ra	m->1	
U-re	g->1	
U-rä	t->1	
U-st	r->1	
U-sä	n->2	
U-te	x->1	
U-ut	v->1	
U-vä	r->1	
U.. 	(->1	
U.Al	l->1	
U.Da	g->1	
U.De	 ->1	t->1	
U.Fr	å->1	
U.Nu	 ->1	
U.Ro	p->1	
U.Vi	 ->3	
U:s 	B->1	E->1	b->6	d->1	e->2	f->3	g->1	h->2	i->6	k->2	l->2	m->4	n->1	o->6	p->3	r->1	s->4	t->2	u->1	
U?He	r->1	
UCK 	n->1	
UCLA	F->1	
UE/N	G->2	
UELL	A->1	
UEN-	g->1	
UF) 	ä->1	
UGFJ	)->2	:->1	
UNIF	I->1	
UNMI	K->3	
USA 	-->1	a->1	e->1	h->1	p->1	
USA,	 ->2	
USA.	J->1	V->1	
USA:	s->1	
USD 	f->1	
USP 	o->1	
Ulst	e->1	
Unda	n->3	
Unde	r->34	
Ungd	o->1	
Unge	f->2	
Unio	n->8	
Uppd	a->1	
Uppe	n->1	
Uppf	ö->1	
Uppg	i->3	
Uppr	ä->1	
Ur d	e->2	
Ur e	n->1	
Ur p	a->1	
Urba	-->1	n->1	
Urqu	i->1	
Ursä	k->1	
Utan	 ->3	
Utbi	l->2	
Utde	l->1	
Utes	t->1	
Utfo	r->2	
Utfö	r->1	
Utgi	f->2	
Utif	r->1	
Utma	n->2	
Utnä	m->2	
Utsk	o->6	
Uttj	ä->1	
Utve	c->1	
Utvi	d->1	
Utvä	r->1	
Uzbe	k->2	
V - 	D->1	R->1	
V an	k->1	
V i 	E->1	f->1	
V-bi	l->1	
V-ka	n->1	
V-pr	o->1	
V-sä	n->1	
VC, 	a->1	
VC-l	e->1	
VC.V	i->1	
VD b	ö->1	
VI i	 ->1	
VII:	e->1	
VIII	 ->2	:->1	
VP (	Ö->2	
VP a	t->2	
VP m	i->1	
VP) 	o->1	
Vad 	a->2	b->13	d->1	e->1	f->2	g->16	h->1	j->5	k->7	m->1	s->9	t->3	u->1	v->7	ä->6	
Vada	n->1	
Vald	e->3	
Vale	n->2	t->1	
Vall	e->3	
Van 	H->3	
Vand	a->1	
Vanl	i->1	
Vape	n->1	
Var 	d->1	f->2	h->1	o->2	s->1	
Vare	 ->2	l->1	
Varf	ö->12	
Varj	e->7	
Vark	e->1	
Vata	n->3	
Velz	e->1	
Vem 	b->2	d->1	k->1	s->2	v->1	
Vems	 ->2	
Vend	é->1	
Vene	z->1	
Vens	t->2	
Verh	e->2	
Verk	s->1	
Vers	a->1	
Vete	n->1	r->1	
Vets	k->1	
Vi a	c->1	l->1	n->17	r->1	v->5	
Vi b	e->27	i->1	o->1	ö->11	
Vi d	e->2	i->5	r->1	
Vi e	r->1	u->1	
Vi f	a->1	i->3	o->2	ä->1	å->14	ö->13	
Vi g	e->1	j->1	o->2	r->1	ö->3	
Vi h	a->91	o->6	y->1	ä->2	å->2	
Vi i	 ->6	n->7	
Vi j	a->1	
Vi k	a->26	o->21	r->8	u->1	ä->4	
Vi l	a->2	i->1	ö->1	
Vi m	e->4	i->1	o->1	å->77	
Vi o	r->1	
Vi p	a->1	l->1	
Vi r	a->1	e->1	i->1	ä->2	ö->1	
Vi s	a->1	e->6	i->1	k->22	o->1	t->9	v->3	ä->3	
Vi t	a->5	i->2	r->3	v->2	y->4	ä->2	
Vi u	n->1	p->6	t->2	
Vi v	a->5	e->15	i->31	ä->9	
Vi ä	n->1	r->34	
Vi ö	n->1	
Vi, 	d->1	
Via 	s->1	
Vich	y->1	
Vid 	E->1	b->1	d->4	e->3	l->1	m->2	s->2	
Vida	r->7	
Vikt	e->1	
Vilj	a->1	
Vilk	a->16	e->8	
Vill	 ->4	k->1	
Vind	e->1	
Viss	a->13	e->2	t->1	
Vitb	o->3	
Vito	r->7	
Vivi	e->1	
Vlaa	m->1	
Voda	f->1	
Volk	s->1	
Von 	W->1	
Värd	e->1	
Värl	d->3	
Väst	b->4	m->1	r->1	
Vår 	d->1	e->1	g->5	i->2	o->1	r->2	u->3	ö->1	
Våra	 ->8	
Vårt	 ->7	
WTO?	E->1	
Waff	e->2	
Wale	s->11	
Wall	s->4	
Wash	i->3	
Web,	 ->1	
West	 ->1	
Wide	 ->1	
Wieb	e->1	
Wiel	a->4	
Wien	 ->3	,->1	
Wilh	e->1	
Woga	u->18	
Worl	d->1	
Wulf	-->2	
Wurt	z->3	
Wye 	P->1	
Wye-	a->2	
Wynn	,->1	
X oc	h->2	
X, f	a->1	
XVII	:->1	I->1	
XXVI	I->2	
YN))	.->1	
Yass	e->1	
York	 ->1	
Ytte	r->3	
Zeel	a->2	
Zime	r->1	
[KOM	(->2	
[SEK	(->1	
].) 	H->1	
].He	r->2	
a "A	m->1	
a "b	a->1	
a "i	r->1	
a "l	ä->1	
a "s	h->1	
a "u	t->1	
a (K	O->1	
a (a	r->1	
a - 	a->3	b->1	d->7	e->1	f->7	g->1	h->2	i->3	j->3	k->2	l->2	m->6	o->7	p->3	r->4	s->5	t->1	u->1	v->1	ä->2	
a -,	 ->1	
a 1 	o->2	p->1	
a 10	 ->2	0->1	
a 12	3->1	5->1	
a 13	3->1	
a 15	 ->1	
a 16	 ->2	7->1	
a 17	0->1	
a 2 	p->2	
a 20	0->1	
a 25	 ->4	0->1	
a 30	 ->1	
a 33	 ->1	
a 35	 ->1	
a 37	0->1	
a 40	 ->1	
a 5 	m->1	
a 55	 ->1	
a 6 	o->1	
a 60	 ->1	
a 70	 ->1	
a 81	 ->4	.->1	
a 85	 ->3	
a 87	,->1	
a 90	-->1	
a Ah	e->1	
a Al	e->1	i->1	t->1	
a Am	s->1	
a At	l->1	
a Az	o->1	
a B 	o->1	
a Ba	l->1	r->2	
a Be	r->2	
a Bo	w->1	
a Br	y->2	
a Co	l->1	s->8	
a Da	l->1	n->1	
a EE	G->1	
a EG	-->5	
a EU	 ->4	-->7	:->4	
a El	i->1	l->1	
a Er	i->2	
a Eu	r->56	
a Ev	a->1	
a FN	:->2	
a FP	Ö->2	
a Fe	i->1	
a Fi	s->1	
a Fl	a->1	o->2	é->1	
a Fr	a->4	
a Fö	r->1	
a Go	l->1	
a Gr	a->1	o->1	
a Ha	i->5	n->1	
a Hi	c->1	
a Hu	l->1	
a IX	 ->1	
a In	t->1	
a Is	r->2	
a Iz	q->1	
a Ja	n->1	
a Je	a->1	r->1	
a Jo	n->1	
a Jö	r->2	
a Ka	r->1	
a Ko	c->2	s->1	u->1	
a Ku	n->1	
a La	n->1	
a Li	b->3	i->1	
a Lo	i->1	u->1	
a Ma	a->1	l->1	r->1	
a Me	l->1	
a Mo	u->9	
a Mu	l->1	
a Na	n->1	t->1	
a Ni	e->1	
a OL	A->1	
a PP	E->1	
a PV	C->1	
a Pa	k->1	l->3	
a Po	e->2	
a Pr	o->1	
a Ra	c->1	
a Ri	i->1	
a Ro	b->1	m->1	t->1	
a Ry	s->1	
a Ré	u->2	
a Sa	l->1	v->1	
a Sc	h->1	
a Sh	e->1	
a St	a->1	
a Su	a->1	
a Sv	e->1	
a TV	-->1	
a Te	r->1	x->1	
a Tu	r->2	
a Ty	s->2	
a UC	K->1	
a Wa	l->1	
a Ze	e->2	
a ab	s->3	
a ad	j->1	m->4	
a af	f->3	
a ag	e->5	g->1	
a ak	t->13	
a al	d->1	k->1	l->66	t->5	
a am	b->8	
a an	 ->1	a->3	b->1	d->36	f->2	g->6	h->2	k->1	l->3	m->4	n->2	o->2	p->1	s->74	t->10	v->28	
a ap	p->2	
a ar	a->1	b->75	g->7	m->2	r->3	t->11	v->3	
a as	p->17	y->2	
a at	l->1	o->4	t->476	
a au	k->1	t->1	
a av	 ->176	,->2	.->1	a->1	d->2	f->1	g->2	l->1	s->40	t->15	v->1	
a ba	k->10	l->2	n->4	r->9	s->5	
a be	 ->6	a->1	b->1	d->14	f->25	g->21	h->31	k->14	l->8	m->3	r->9	s->102	t->112	u->1	v->18	
a bi	b->3	d->18	e->2	l->64	n->2	s->2	t->1	
a bj	u->1	
a bl	.->1	a->3	i->25	
a bo	 ->1	l->3	m->1	r->18	s->2	t->2	
a br	a->5	i->9	o->10	u->2	ä->3	å->2	
a bu	d->24	
a by	g->7	r->4	
a bä	r->4	s->2	t->7	
a bå	d->6	t->3	
a bö	r->26	
a ca	n->1	
a ce	n->10	r->4	
a ch	a->5	
a ci	t->1	v->1	
a da	 ->1	g->20	m->38	n->1	t->4	
a de	 ->184	b->42	c->2	f->3	l->73	m->82	n->209	p->1	r->8	s->68	t->237	
a di	a->9	e->1	f->3	g->2	k->2	l->1	m->9	p->4	r->48	s->20	
a dj	u->7	
a do	g->1	k->16	m->15	
a dr	a->12	i->5	o->1	u->1	ö->1	
a du	b->2	m->2	
a dy	n->1	r->3	
a dä	r->20	
a då	 ->5	l->1	
a dö	d->2	m->1	r->2	t->1	
a ef	f->26	t->23	
a eg	e->1	n->26	o->1	
a ek	o->34	v->1	
a el	e->4	i->1	l->48	v->1	
a em	e->5	o->12	
a en	 ->349	,->1	a->2	b->1	d->4	e->44	g->2	h->12	i->1	k->3	l->7	o->2	s->4	v->2	
a er	 ->39	,->4	a->5	b->4	f->12	i->2	k->2	s->2	t->1	
a et	a->3	c->2	n->3	t->178	
a eu	r->35	
a ev	e->3	
a ex	a->2	e->10	i->2	p->4	t->7	
a fa	k->11	l->54	m->4	n->3	r->32	s->14	t->8	
a fe	l->3	m->7	n->1	
a fi	l->2	n->21	s->8	
a fl	a->1	e->14	i->1	o->1	y->2	ö->1	
a fo	g->1	l->32	n->10	r->74	s->1	t->1	
a fr	a->117	e->5	i->18	o->1	u->7	ä->2	å->287	
a fu	l->7	n->11	s->2	
a fy	r->1	
a fä	r->1	s->1	
a få	 ->15	g->3	n->2	r->18	
a fö	d->3	l->30	r->866	
a ga	l->2	m->5	n->2	r->11	v->1	
a ge	 ->9	m->65	n->53	o->1	r->2	s->1	
a gi	c->1	f->1	g->1	l->4	v->11	
a gj	o->6	
a gl	a->1	ä->3	ö->2	
a gn	ä->1	
a go	d->15	
a gr	a->20	e->2	o->1	u->91	y->1	ä->17	ö->1	
a gä	c->1	l->27	r->2	
a gå	 ->2	n->40	r->5	
a gö	r->35	
a ha	 ->10	d->8	f->1	l->2	m->8	n->72	p->1	r->111	t->1	v->4	
a he	l->28	m->4	n->7	r->6	t->1	
a hi	n->14	s->7	t->5	
a hj	ä->6	
a ho	m->1	n->12	p->4	r->1	s->6	t->3	
a hu	m->1	n->2	r->34	s->2	v->5	
a hy	l->1	p->1	s->1	
a hä	f->1	l->4	n->52	r->11	v->3	
a hå	l->19	r->3	v->1	
a hö	g->19	j->1	l->1	r->7	
a i 	A->2	B->1	C->4	D->3	E->50	F->3	G->1	I->2	K->5	L->4	M->1	P->3	R->2	S->1	T->5	U->1	W->1	a->12	b->5	d->90	e->34	f->30	g->9	h->7	i->3	j->1	k->18	l->6	m->19	n->3	o->7	p->7	r->5	s->26	t->5	u->10	v->20	y->2	Ö->6	ä->1	å->1	ö->3	
a i.	D->1	N->1	S->1	
a ia	k->2	
a ib	l->1	
a ic	k->2	
a id	e->6	é->10	
a if	a->1	r->4	
a ig	e->9	n->1	å->3	
a ih	j->1	o->3	å->14	
a ik	a->1	
a il	l->2	
a im	a->1	m->1	p->3	
a in	 ->33	,->1	b->3	c->3	d->15	f->27	g->2	h->1	i->24	k->5	l->13	n->26	o->25	r->6	s->97	t->132	v->15	
a ir	r->1	
a is	o->1	ä->2	
a it	u->14	
a iv	e->1	
a ja	,->1	g->5	
a jo	b->3	r->14	
a ju	l->1	r->6	s->2	
a jä	m->8	r->1	
a ka	l->1	m->31	n->56	p->4	r->8	t->18	
a ke	d->2	
a ki	l->1	n->1	
a kl	.->1	a->21	i->7	o->1	y->3	
a kn	a->1	o->1	u->1	y->2	
a ko	a->1	d->3	k->1	l->102	m->230	n->189	p->1	r->15	s->24	
a kr	a->34	e->5	i->29	o->1	ä->7	å->1	
a ku	l->14	n->13	r->1	s->14	
a kv	a->19	i->14	o->3	ä->1	
a ky	l->1	
a kä	l->3	n->13	r->17	
a kö	l->1	p->1	
a la	b->2	d->1	g->27	n->20	r->2	
a le	d->32	g->1	k->1	v->5	
a li	b->9	g->9	k->15	n->3	s->2	t->8	v->27	
a lj	u->2	
a lo	b->1	k->10	v->1	
a lu	c->2	g->1	
a ly	c->1	f->1	s->3	
a lä	g->11	k->1	m->12	n->70	r->5	s->1	t->3	
a lå	n->4	t->1	
a lö	f->6	n->3	p->1	s->20	
a ma	j->6	k->5	n->12	r->28	s->4	t->8	x->1	
a me	d->430	g->1	k->3	l->21	n->16	r->18	s->3	t->8	
a mi	g->23	k->1	l->30	n->56	s->14	t->23	
a mo	b->2	d->14	m->1	n->8	r->1	t->32	
a mu	n->2	r->1	s->1	
a my	c->46	g->1	n->55	
a mä	k->1	n->26	r->2	t->1	
a må	l->55	n->24	s->62	t->2	
a mö	d->1	j->57	r->1	t->7	
a na	i->1	m->2	r->1	t->43	
a ne	d->8	g->2	j->1	o->1	r->1	
a ni	 ->4	m->1	o->2	v->14	
a no	g->4	n->2	r->8	t->1	
a nr	 ->26	
a nu	 ->1	?->1	l->1	n->1	v->1	
a ny	 ->1	a->30	c->3	h->5	l->1	t->5	å->1	
a nä	m->13	r->35	s->4	t->10	
a nå	 ->2	g->78	t->1	
a nö	d->9	j->3	t->1	
a oa	v->1	
a ob	a->4	e->7	l->3	
a oc	h->539	k->20	
a od	d->1	u->1	
a oe	g->2	n->1	
a of	e->1	f->13	r->1	t->2	ö->2	
a og	e->1	
a oi	n->1	
a oj	ä->2	
a ok	l->3	o->1	
a ol	i->15	j->8	y->10	ö->1	
a om	 ->274	,->6	.->4	b->5	e->2	f->9	g->2	r->93	s->31	v->3	ö->1	
a on	d->1	ö->2	
a op	a->1	e->4	i->1	p->1	t->2	
a or	d->121	e->1	g->32	i->3	o->9	s->8	t->1	ä->1	
a os	s->64	ä->1	
a ot	i->1	
a pa	k->1	l->1	r->130	s->1	t->1	
a pe	d->1	k->1	l->2	n->22	r->23	s->1	
a ph	t->1	
a pi	r->1	
a pl	a->27	e->1	ä->1	
a po	l->82	p->1	r->1	s->6	
a pr	a->9	e->18	i->46	o->179	ö->1	
a pu	b->1	m->1	n->78	
a på	 ->197	,->4	.->3	:->1	f->1	g->2	m->5	p->9	s->4	t->1	v->1	
a ra	d->5	m->13	n->12	p->38	
a re	a->11	d->15	f->33	g->191	k->8	l->6	n->7	p->8	s->92	t->1	v->5	
a ri	g->1	k->40	m->1	s->18	
a ro	,->1	l->6	m->1	
a ru	b->1	m->19	n->3	t->4	
a ry	g->1	
a rä	c->1	d->6	k->4	t->87	
a rå	d->44	o->1	t->1	
a rö	r->20	s->11	t->2	
a s.	k->1	
a sa	d->4	g->1	k->32	m->122	n->5	t->4	
a sc	e->4	
a se	 ->7	d->6	g->1	i->1	k->35	n->5	r->4	s->2	t->4	x->2	
a si	d->41	f->8	g->120	m->1	n->75	t->59	
a sj	u->4	ä->14	ö->8	
a sk	a->88	e->10	i->30	j->1	o->9	r->11	u->32	y->10	ä->21	ö->2	
a sl	a->17	u->25	ä->1	å->3	
a sm	u->2	å->11	
a sn	a->10	e->2	ä->1	
a so	c->37	l->4	m->219	r->1	
a sp	a->1	e->31	o->1	r->2	ä->4	å->1	ö->2	
a st	a->70	e->10	i->4	o->33	r->55	u->10	y->6	ä->26	å->71	ö->101	
a su	b->7	m->7	t->1	v->1	
a sv	a->10	å->21	
a sy	d->1	f->8	m->3	n->21	s->49	
a sä	g->34	k->18	m->1	n->4	r->8	s->1	t->65	
a så	 ->34	.->2	d->11	g->1	n->2	s->2	v->1	
a sö	n->1	r->1	
a t.	o->2	
a ta	 ->18	c->15	g->5	k->1	l->19	n->13	r->6	s->4	x->1	
a te	a->1	c->3	k->9	l->1	m->2	n->6	r->11	x->18	
a ti	d->32	g->1	l->328	m->2	n->1	o->1	t->1	
a tj	ä->27	
a to	g->6	l->5	m->1	n->4	r->3	t->4	x->1	
a tr	a->26	e->17	i->1	o->7	u->3	y->3	ä->6	å->2	ö->1	
a tu	n->3	r->1	s->2	
a tv	i->8	å->26	
a ty	c->6	d->9	n->4	p->18	s->2	
a tä	c->1	n->4	v->1	
a tå	g->1	l->1	
a ul	t->1	
a um	g->1	
a un	d->64	g->4	i->270	
a up	p->198	
a ur	 ->9	a->1	h->1	s->4	v->1	
a ut	 ->24	.->2	:->1	a->20	b->9	e->2	f->10	g->13	h->1	i->1	k->13	l->3	m->10	n->4	r->4	s->20	t->19	v->71	ö->1	
a va	c->2	d->28	g->1	k->2	l->23	n->7	p->8	r->70	t->1	
a ve	c->21	d->1	l->1	m->1	n->1	r->69	t->13	
a vi	 ->10	c->3	d->28	k->38	l->73	n->6	r->1	s->34	t->5	
a vo	n->2	r->2	t->2	
a vr	a->2	
a vä	d->3	g->15	k->1	l->17	n->5	r->42	s->5	v->3	x->5	
a vå	g->2	l->4	r->46	
a yr	k->3	
a yt	l->1	t->15	
a Ös	t->6	
a äg	a->6	d->1	e->1	n->1	t->1	
a äm	b->3	n->17	
a än	 ->4	d->95	n->7	t->3	
a är	 ->292	,->3	.->3	:->2	a->1	e->4	l->2	
a äv	e->10	
a å 	m->2	
a åk	l->8	
a år	 ->16	,->7	.->5	e->24	h->2	l->2	s->3	t->1	
a ås	a->1	i->5	k->1	t->2	
a åt	 ->2	.->1	a->22	e->22	f->1	g->99	
a öa	r->3	
a öd	e->2	
a ög	a->1	o->5	
a ök	a->8	n->2	
a ön	s->7	
a öp	p->6	
a ör	e->1	o->1	
a ös	t->6	
a öv	e->80	r->2	
a! D	e->1	
a! V	i->1	
a!Av	 ->1	
a!De	n->1	t->3	
a!Fr	u->3	
a!Fö	r->1	
a!He	r->2	
a!Ja	g->1	
a!Lå	t->1	
a!Mä	n->1	
a!Om	 ->1	
a!Äv	e->1	
a" b	i->1	
a" s	o->1	
a" v	a->1	
a", 	v->1	
a"..	 ->1	
a".B	a->1	
a".D	e->2	
a".H	i->1	
a".J	u->1	
a".K	i->1	
a"; 	ö->1	
a"in	d->1	
a) a	d->1	
a) b	ä->1	
a, 1	6->1	
a, 5	0->1	
a, B	r->1	
a, E	v->1	
a, J	a->1	
a, K	v->1	
a, S	a->1	c->1	
a, a	d->1	l->3	n->2	r->2	t->24	v->4	
a, b	a->1	e->1	i->2	l->5	o->1	å->1	
a, c	o->1	
a, d	e->36	j->2	v->6	ä->6	å->3	ö->1	
a, e	f->12	k->1	l->4	n->11	r->1	t->5	u->1	x->1	
a, f	o->1	r->13	u->1	å->2	ö->38	
a, g	a->1	e->3	ö->1	
a, h	a->14	e->14	j->1	u->5	ö->2	
a, i	 ->23	b->1	n->15	
a, j	a->3	o->1	u->2	
a, k	a->7	o->9	
a, l	e->1	i->6	ä->1	å->3	
a, m	e->48	i->4	o->1	å->4	
a, n	a->2	e->2	u->1	y->1	ä->8	å->4	
a, o	a->1	b->1	c->87	m->16	r->1	
a, p	a->1	e->1	r->4	å->4	
a, r	a->2	e->7	i->1	ä->2	
a, s	a->5	e->2	k->3	l->1	n->1	o->46	t->5	v->1	ä->4	å->20	ö->1	
a, t	.->1	a->1	e->1	i->10	j->1	o->1	r->5	u->1	y->1	ö->1	
a, u	n->3	p->1	t->22	
a, v	a->8	e->2	i->35	o->1	ä->1	
a, ä	g->1	r->8	v->4	
a, å	t->4	
a, ö	p->1	v->1	
a-, 	S->1	
a-Is	r->1	
a-Ro	m->1	
a-ol	y->1	
a. 1	2->1	
a. D	e->2	ä->1	å->1	
a. E	n->1	
a. F	ö->1	
a. H	å->1	
a. J	a->1	
a. K	o->1	ä->1	
a. M	e->3	
a. S	o->1	
a. V	a->2	
a. a	r->1	t->1	
a. b	e->1	
a. d	e->1	
a. e	n->1	t->1	
a. f	å->1	ö->4	
a. g	e->1	ö->1	
a. i	 ->2	
a. k	r->1	
a. m	e->1	
a. n	ä->3	
a. o	l->1	m->1	
a. p	å->1	
a. s	k->2	t->1	
a. u	n->1	
a. v	a->1	
a. Å	t->1	
a.(I	h->1	
a.(P	a->1	
a.(T	a->2	
a.)B	e->1	
a.)F	r->1	
a.- 	(->4	
a.. 	H->1	T->1	
a..(	E->1	I->1	N->1	
a...	(->1	L->1	
a.18	 ->1	
a.Al	l->10	
a.Am	s->1	
a.An	n->2	s->1	
a.Av	 ->5	
a.Ba	k->2	
a.Be	r->2	s->2	t->1	
a.Bi	l->1	
a.Bl	a->1	
a.Bo	r->1	
a.Co	r->1	
a.De	 ->8	n->24	s->9	t->114	
a.Do	c->1	
a.Dä	r->14	
a.Då	 ->2	
a.EG	-->1	
a.Ef	t->8	
a.Em	e->3	
a.En	 ->9	k->1	l->3	
a.Et	t->8	
a.Eu	r->4	
a.Fa	c->2	
a.Fr	a->1	u->4	å->3	
a.Fö	l->1	r->25	
a.Ge	m->1	r->1	
a.Gi	v->1	
a.Ha	n->2	
a.He	l->1	r->33	
a.Hu	l->1	r->3	
a.Hä	r->4	
a.I 	E->1	a->1	b->1	d->7	e->2	f->5	l->4	m->1	p->3	r->2	s->2	t->1	v->2	ö->1	
a.Ib	l->2	
a.In	g->1	o->3	t->3	
a.Ja	g->98	
a.Ju	s->2	
a.Ka	f->1	n->1	
a.Ko	m->10	n->2	
a.Kä	r->2	
a.Li	k->1	v->1	
a.Lä	g->1	
a.Lå	t->6	
a.Ma	j->1	n->3	
a.Me	d->11	n->27	
a.Mi	n->10	
a.Må	n->2	
a.Na	t->2	
a.Ni	 ->6	
a.Nu	 ->3	
a.Nä	r->10	
a.Oc	h->9	
a.Om	 ->11	
a.Or	d->1	s->1	
a.Pa	r->1	
a.Pe	r->1	
a.Pr	e->2	o->2	
a.På	 ->11	
a.Re	g->1	s->1	
a.Ru	m->1	
a.Rå	d->2	
a.Sa	m->1	
a.Se	d->2	
a.Si	t->2	
a.Sj	u->1	
a.Sk	y->1	
a.Sl	u->3	
a.Sm	å->1	
a.So	m->6	
a.St	a->1	ö->2	
a.Sy	f->1	
a.Sä	g->1	
a.Så	 ->3	n->1	
a.Ta	c->2	d->1	
a.Ti	l->2	
a.To	p->1	
a.Tr	o->5	
a.Ty	 ->1	
a.Un	d->3	g->1	
a.Up	p->2	
a.Ur	 ->1	
a.Ut	a->1	b->1	d->1	f->1	n->1	
a.Va	d->10	r->3	
a.Ve	m->1	r->1	
a.Vi	 ->72	a->1	d->4	k->1	l->1	s->2	
a.Vä	r->1	s->1	
a.Vå	r->3	
a.Än	 ->1	d->1	t->1	
a.Är	 ->3	
a.Äv	e->5	
a.Å 	a->2	
a.År	 ->1	
a.Öv	e->1	
a/Eu	r->1	
a/ha	l->1	
a/sa	m->1	
a: "	D->1	i->1	
a: D	e->1	
a: F	ö->2	
a: I	 ->2	
a: J	a->2	
a: N	ä->1	
a: V	a->1	e->1	
a: a	n->1	t->1	
a: d	e->1	
a: g	e->1	
a: h	u->2	
a: m	a->1	
a: o	m->1	
a: r	ä->1	
a: s	k->1	
a: u	n->1	p->1	t->1	
a: v	e->2	i->3	
a: Ä	v->1	
a:Fö	r->1	
a; d	e->1	
a; e	n->1	
a; f	ö->2	
a; j	a->2	
a; k	o->1	
a; l	o->1	
a; o	c->1	
a; p	u->1	
a; v	i->2	
a?"J	a->1	
a?. 	(->1	
a?An	s->1	
a?Av	s->1	
a?De	 ->1	n->1	t->6	
a?Et	t->1	
a?Fr	u->1	
a?Fö	r->1	
a?Ha	r->1	
a?He	r->1	
a?Hu	r->1	
a?I 	F->1	d->1	
a?In	i->1	
a?Ja	g->3	
a?Jo	,->1	
a?Ma	n->1	
a?Ne	j->1	
a?Nä	r->1	
a?Pr	o->1	
a?På	 ->1	
a?Sv	a->1	
a?Va	d->3	
a?Vi	 ->2	l->1	s->1	
a?Är	 ->1	
aHer	r->1	
aNäs	t->2	
aaff	ä->1	
aams	 ->1	
aan 	f->1	
aan.	V->1	
aans	 ->5	
aard	e->1	
aast	r->6	
ab s	k->1	
abar	é->1	
abas	e->1	
abb 	h->1	o->2	v->1	
abba	 ->11	d->27	r->14	s->10	t->12	
abbt	 ->34	,->3	.->6	
abbv	a->1	
abeh	a->7	
abek	ä->1	
abel	 ->5	!->1	,->3	.->4	l->6	t->21	
aber	g->1	
abet	e->1	h->1	
abil	 ->2	a->2	i->19	t->2	
abin	e->3	
abis	e->1	k->6	
abla	 ->9	"->1	,->1	.->3	n->1	
able	r->13	
ablo	n->1	
aboc	k->2	
abon	 ->4	,->1	.->1	m->2	
abor	a->3	
abre	p->1	
abri	e->3	k->1	
abso	l->40	r->1	
abst	a->2	r->1	
absu	r->3	
abu 	i->1	
abuk	t->2	
abul	a->1	
abvä	r->1	
ac b	l->1	ö->1	
ac o	s->1	
ac",	 ->1	
ac-s	y->1	
aca 	M->3	s->1	
acao	 ->1	
acce	p->88	
ace 	o->1	
ace.	D->1	J->1	
acer	a->15	i->2	
aceu	t->1	
acil	l->1	
acio	 ->7	,->3	.->2	:->1	s->2	
acis	 ->1	-->1	
acit	e->5	
ack 	a->1	f->11	g->2	h->1	m->1	o->4	p->1	s->17	t->11	v->7	
ack,	 ->15	
ack-	p->1	
ack.	F->1	H->1	J->1	
acka	 ->84	r->21	t->3	
ackd	e->8	
acke	n->1	r->2	
ackf	ö->7	
ackl	a->2	
ackn	i->6	
acko	r->1	
ackr	a->6	
acks	 ->1	a->9	o->2	
aco-	a->1	
acob	 ->2	
acqu	e->3	i->1	
acto	r->1	
acèt	e->1	
ad -	 ->1	
ad A	d->1	
ad B	N->1	
ad E	u->1	
ad F	P->1	
ad G	u->1	
ad K	u->2	
ad S	y->1	
ad a	l->1	n->10	r->1	t->16	v->19	
ad b	e->31	i->2	l->2	o->1	y->1	
ad d	a->4	e->31	o->3	å->1	
ad e	f->2	l->5	n->6	r->1	t->1	u->2	
ad f	e->1	i->1	l->1	o->2	r->5	ö->23	
ad g	e->2	i->1	r->2	ä->60	ö->1	
ad h	a->5	o->2	ä->3	
ad i	 ->14	d->1	m->1	n->12	
ad j	a->12	u->1	ä->1	
ad k	a->5	o->27	r->1	v->1	
ad l	e->1	
ad m	a->17	e->9	i->2	o->1	å->3	
ad n	a->2	i->4	å->1	
ad o	c->11	l->2	m->22	r->1	
ad p	a->1	e->1	o->4	r->3	u->1	å->9	
ad r	e->3	i->1	o->2	ä->4	å->1	
ad s	a->3	e->3	i->3	k->6	m->2	n->1	o->67	t->5	u->1	y->8	ä->4	
ad t	a->1	i->13	j->1	r->2	ä->2	
ad u	n->1	p->1	r->1	t->4	
ad v	a->1	e->7	i->26	o->1	å->3	
ad y	r->1	
ad ä	n->1	r->12	v->1	
ad ö	p->1	v->18	
ad, 	"->1	a->2	e->2	f->1	h->1	i->2	m->3	o->1	s->2	t->2	u->1	v->1	ä->1	
ad-k	o->1	
ad."	M->1	
ad.(	S->1	
ad.D	e->7	
ad.E	u->1	
ad.F	r->1	
ad.H	e->6	
ad.J	a->4	
ad.K	o->2	
ad.M	e->4	ä->1	å->1	
ad.O	m->14	
ad.P	a->1	
ad.R	e->1	
ad.S	u->1	
ad.U	t->1	
ad.V	e->1	i->2	
ad: 	e->1	
ad; 	d->1	
ad?D	ä->1	
ad?H	e->1	
ad?V	i->1	
ada 	E->1	d->4	e->1	f->1	k->1	o->1	r->1	s->1	ö->2	
ada!	D->1	
ada,	 ->3	
ada.	M->1	
adad	e->2	
adag	a->1	
adak	i->1	
adan	 ->1	.->1	a->2	
adar	 ->6	
adat	.->1	s->3	
adda	d->1	
adde	 ->2	r->1	
addi	n->2	t->1	
ade 	"->3	-->3	1->2	2->1	4->1	E->4	F->1	H->3	I->1	N->1	O->1	T->1	V->1	a->62	b->25	d->37	e->22	f->51	g->12	h->16	i->53	j->14	k->61	l->7	m->49	n->13	o->70	p->36	r->28	s->59	t->32	u->16	v->40	y->1	Ö->1	ä->6	å->7	ö->6	
ade,	 ->27	
ade.	 ->2	A->2	D->7	E->2	F->2	H->3	J->2	M->1	P->1	S->5	T->3	V->2	
ade:	 ->1	
ade?	J->1	
adee	r->2	
adef	o->1	
adei	r->2	
adek	v->5	
adel	s->2	
adem	i->2	o->2	
aden	 ->85	)->3	,->29	.->31	s->19	
ader	 ->64	,->12	-->1	.->18	;->1	a->4	n->81	s->3	
ades	 ->107	,->5	.->6	t->1	
adet	 ->2	.->1	
adga	 ->14	,->1	d->1	n->10	r->2	
adgo	r->1	
adie	t->4	
adik	a->16	
adin	g->1	s->1	
adio	l->2	
adit	i->19	
adiu	m->4	
adiz	 ->3	,->1	-->1	
adje	k->2	
adko	m->24	
adli	g->10	n->1	
admi	n->25	u->3	
ado,	 ->1	
ador	 ->12	,->4	.->2	n->8	
adou	 ->1	
adox	,->1	a->5	
adra	g->3	
adri	a->1	d->3	
ads 	b->1	
ads-	 ->1	i->2	n->1	
ads/	i->1	
adsa	k->1	n->3	r->1	
adsb	e->5	
adsc	e->1	
adsd	o->1	
adse	f->4	k->14	
adsf	r->4	ö->1	
adsi	n->3	
adsk	r->1	
adsl	i->1	å->1	
adsm	y->1	ö->1	
adsn	i->1	
adso	m->1	r->1	
adsp	r->6	
adss	t->3	
adst	i->1	
adsu	p->1	
adsv	e->1	i->2	
adt,	 ->1	
advi	s->3	
advo	k->5	
adzj	i->5	
adör	 ->1	
ael 	-->1	a->4	b->1	d->1	f->2	h->1	i->1	l->1	m->1	o->10	v->1	
ael,	 ->4	
ael-	S->1	
ael.	D->2	N->1	S->1	
ael?	E->1	
aele	r->5	
aeli	s->15	
aelk	r->1	
aels	 ->6	
af o	m->1	
afae	l->3	
afat	s->1	
afet	y->1	
aff 	o->2	
aff,	 ->1	
aff-	 ->2	
affa	 ->20	d->3	n->1	r->1	s->3	t->1	
affb	e->1	
affe	n->3	
affl	a->1	
affp	r->2	
affr	ä->28	
affä	r->12	
afi 	p->1	
afi.	D->1	V->1	
afik	 ->2	-->1	.->2	e->3	l->1	
afin	.->1	
afis	k->10	
afly	k->1	
afon	e->1	
afor	 ->1	
afra	n->1	
afri	k->2	
afry	t->2	
afrå	g->12	
aft 	2->1	a->6	b->2	d->4	e->4	f->9	h->1	i->4	k->1	m->5	n->4	o->4	p->4	s->13	t->4	u->2	v->3	ä->1	
aft,	 ->11	
aft.	D->2	H->1	M->1	V->2	
aft?	 ->1	N->1	
afte	n->17	r->9	
aftf	u->12	
afti	g->34	
afto	n->1	
afts	a->4	o->1	p->2	r->1	s->1	v->1	
aftt	a->1	r->4	
aftv	e->8	
ag -	 ->11	
ag 1	 ->2	,->2	0->5	1->1	2->1	3->1	5->1	7->1	8->2	9->3	
ag 2	,->2	2->3	3->1	6->1	
ag 3	 ->1	4->1	8->3	
ag 4	 ->1	.->2	3->1	4->1	5->3	
ag 5	,->2	
ag 6	 ->2	
ag G	a->1	
ag I	N->1	
ag a	b->1	c->2	l->3	n->94	t->87	v->22	
ag b	a->9	e->58	i->1	l->8	o->1	ö->4	
ag c	i->2	
ag d	e->18	o->3	r->3	ä->5	å->1	ö->1	
ag e	f->2	l->1	m->6	n->12	r->13	t->3	
ag f	a->1	i->5	o->5	r->51	u->2	å->11	ö->109	
ag g	a->3	e->9	i->1	j->2	l->10	o->1	r->10	ä->10	å->1	ö->2	
ag h	a->115	e->9	i->1	o->55	u->1	ä->16	å->14	ö->7	
ag i	 ->50	,->1	n->88	
ag j	a->1	u->2	ä->1	
ag k	a->65	l->4	o->43	r->1	u->2	ä->10	ö->1	
ag l	a->4	e->3	i->3	y->7	ä->6	å->1	ö->1	
ag m	a->1	e->30	i->21	o->4	y->4	ä->1	å->23	
ag n	a->5	i->2	o->5	u->6	y->2	ä->13	ö->1	
ag o	c->52	f->1	m->28	r->2	s->1	
ag p	e->5	l->1	o->5	r->2	å->19	
ag r	e->20	i->3	ä->6	å->2	ö->13	
ag s	a->12	e->16	j->14	k->159	o->85	p->2	t->21	v->2	y->6	ä->37	å->4	
ag t	a->52	i->86	o->2	r->115	v->4	y->46	ä->17	
ag u	n->11	p->38	t->19	
ag v	a->12	e->31	i->270	ä->27	å->2	
ag Ö	s->1	
ag ä	g->1	l->1	n->5	r->113	v->2	
ag å	 ->2	t->5	
ag ö	n->6	v->7	
ag, 	a->4	b->2	d->5	e->10	f->11	g->2	h->4	i->5	l->3	m->10	n->3	o->10	p->1	s->16	t->5	u->5	v->7	ä->6	
ag. 	D->1	H->1	P->1	
ag.(	A->1	
ag.)	F->2	H->1	
ag..	 ->1	
ag.A	n->1	r->1	v->1	
ag.B	e->2	
ag.D	e->19	i->1	ä->3	
ag.E	f->2	r->1	
ag.F	r->3	ö->5	
ag.G	e->1	
ag.H	e->6	u->1	y->1	
ag.I	 ->6	n->1	
ag.J	a->13	u->1	
ag.K	a->1	o->3	
ag.L	i->1	å->1	
ag.M	e->1	å->2	
ag.O	c->1	m->1	
ag.P	a->1	
ag.R	a->1	e->1	
ag.S	k->2	y->1	
ag.T	i->2	
ag.U	n->1	
ag.V	a->2	i->6	å->1	
ag: 	d->1	j->1	
ag:D	e->1	
ag; 	s->1	
ag?D	e->1	
ag?F	i->1	r->1	ö->1	
aga 	2->1	H->1	a->3	d->7	j->1	n->1	o->1	r->2	s->1	
aga!	F->1	
aga,	 ->2	
aga.	D->1	F->1	V->1	
agad	e->5	
agan	 ->2	d->224	s->3	
agar	 ->39	,->5	.->5	a->2	e->71	l->3	m->14	n->25	s->2	v->1	ä->1	
agas	 ->3	,->1	.->1	k->1	t->2	
agat	 ->1	e->2	s->2	
agav	 ->3	
agba	r->15	
agd 	a->1	i->1	o->1	p->1	
agd,	 ->1	
agda	 ->6	.->1	
age 	p->1	s->1	
aged	i->4	
agel	,->1	s->5	
agem	a->9	
agen	 ->126	!->1	,->15	.->22	:->2	;->1	d->1	s->55	t->1	
ager	 ->2	.->1	a->69	k->1	
ages	-->1	
aget	 ->136	)->4	,->19	.->34	:->1	;->1	?->1	s->18	t->1	
agfö	r->5	
agg 	d->1	f->1	i->1	m->1	o->1	s->1	
agg,	 ->7	
agg.	D->1	F->1	K->1	M->1	N->1	
agg;	 ->1	
agga	 ->2	d->2	n->1	
agge	n->2	
aggn	i->1	
aggo	r->1	
aggr	e->1	
agh 	m->1	
aghe	t->12	
agin	ä->1	
agis	k->6	
agit	 ->95	,->2	.->4	a->1	s->27	
agiv	a->2	i->1	
agli	g->35	
agma	r->1	t->1	
agn 	f->3	
agna	 ->24	,->1	.->2	d->4	r->2	t->3	
agne	 ->7	-->1	n->2	r->1	s->1	
agni	n->69	s->1	t->1	
agog	e->1	i->4	
agol	f->4	
agom	 ->1	å->3	
agor	 ->2	?->1	d->52	n->2	
agos	k->1	
agra	f->3	n->1	r->2	
agre	n->1	
agro	t->1	
agru	p->1	
ags 	a->9	d->1	f->8	i->2	m->1	o->3	p->2	r->2	s->3	u->2	v->2	
ags,	 ->2	
ags.	F->1	
agsa	m->3	n->1	r->1	v->1	
agsb	e->1	o->1	
agsd	e->1	
agse	k->5	
agsf	a->1	ä->1	ö->3	
agsg	i->8	r->2	
agsi	n->1	
agsj	u->2	
agsk	o->1	r->1	
agsl	i->1	ä->2	
agsm	ä->2	
agsn	a->1	e->1	
agsr	e->5	å->2	
agss	i->1	t->3	
agst	a->1	e->2	i->131	
agsä	n->3	
agt 	-->1	4->1	a->15	b->2	d->2	e->1	f->30	i->4	j->1	m->3	n->10	o->1	s->2	ä->1	
agt,	 ->9	
agt.	 ->1	J->1	
agte	x->2	
agts	 ->36	,->2	
ague	,->1	
agån	g->10	
ahan	d->1	
ahus	 ->1	
ahål	l->43	
ai L	a->7	
aide	r->37	
aids	 ->2	-->1	p->2	
ail 	m->1	
aill	e->1	
ailu	r->1	
ain"	,->1	
ain,	 ->1	
aine	 ->2	,->1	
ains	a->2	t->30	
aint	-->1	
aire	.->1	
aiva	 ->1	
aivi	t->1	
aiwa	n->1	
aj 1	9->3	
aj 2	0->1	
aj f	ö->1	
aj, 	o->1	
aj.J	a->1	
aj.T	o->1	
ajor	i->42	
ajou	r->1	
ak a	t->4	
ak b	e->2	
ak f	ö->1	
ak g	ä->3	
ak h	a->3	o->1	ä->1	
ak i	 ->1	n->1	
ak j	a->1	
ak k	o->1	u->1	
ak l	o->1	
ak m	e->3	o->1	å->1	
ak n	ä->1	
ak s	a->1	e->1	j->1	o->9	
ak t	i->3	
ak u	t->1	
ak v	a->2	i->4	
ak ä	r->2	
ak ö	v->1	
ak, 	a->1	b->1	h->1	m->1	s->1	v->1	
ak.A	t->1	
ak.D	e->3	
ak.E	t->1	
ak.N	i->1	
ak.T	r->1	y->1	
ak: 	g->1	
ak?N	e->1	
aka 	-->1	E->1	a->2	b->3	d->6	e->3	f->3	g->3	i->4	j->1	k->1	m->5	o->8	p->2	r->2	t->10	v->1	ö->1	
aka.	D->1	I->2	L->1	M->1	
aka?	I->1	
akad	e->4	r->3	
akag	å->4	
akam	m->1	
akar	 ->8	e->1	
akas	 ->4	s->1	
akat	 ->5	.->2	s->2	
akav	i->4	
akdö	r->1	
ake,	 ->1	
akel	 ->3	
aken	 ->7	,->2	.->1	:->1	?->1	s->3	
aker	 ->25	,->3	.->5	:->1	n->11	
aket	 ->6	.->1	e->3	
akfö	r->1	
akgr	u->31	
akie	n->1	
akis	 ->3	!->1	b->1	k->1	t->5	
akku	n->2	
akla	s->1	
akli	g->11	
aklu	k->1	
akna	,->1	d->5	r->12	s->20	t->2	
akni	n->14	
akol	o->1	
akom	 ->21	,->1	l->1	r->2	
akon	v->1	
akop	o->5	
akpr	o->1	
akre	r->1	
akro	e->5	f->1	
akry	.->1	g->1	
aks 	b->1	d->1	p->1	s->1	
aksa	m->9	
akso	d->1	
akst	a->1	
akt 	-->1	a->3	b->1	d->4	e->1	f->7	h->2	i->3	l->1	m->9	o->10	p->5	s->1	u->2	v->3	ä->1	
akt,	 ->3	
akt.	B->2	D->2	J->2	M->2	V->1	
akt:	 ->1	
akta	 ->30	.->1	d->1	i->2	n->10	r->24	s->16	t->8	
aktb	a->2	e->2	
aktd	e->1	i->1	
akte	n->12	r->20	t->1	
aktf	a->1	ö->1	
akth	a->1	e->1	å->1	
akti	e->3	g->34	k->12	o->17	s->74	v->37	
aktk	o->1	
aktl	i->14	ö->3	
aktm	e->2	i->1	
akto	r->24	
aktt	a->8	
aktu	a->1	e->31	m->68	
aktä	r->9	
aktö	r->13	
akul	ä->1	
akut	a->1	
akuu	m->2	
akäm	n->1	
akåt	 ->2	s->1	
al -	 ->2	
al C	o->1	
al D	e->1	
al I	n->2	
al K	a->1	
al U	l->1	
al a	r->1	t->1	v->25	
al b	e->5	i->5	r->1	
al c	o->1	
al d	e->4	u->2	
al e	f->2	l->1	n->1	
al f	o->1	r->9	å->1	ö->9	
al g	ö->1	
al h	a->2	ä->1	
al i	 ->8	n->12	
al k	a->2	o->2	v->2	
al l	ä->3	
al m	a->1	e->16	i->1	o->1	ä->1	å->3	ö->1	
al n	i->3	o->1	y->1	
al o	c->22	m->11	r->1	
al p	e->1	l->3	o->2	r->5	å->2	
al r	a->1	e->3	i->1	o->3	ä->2	
al s	a->9	e->1	i->3	j->1	k->3	o->26	t->5	v->2	y->1	ä->2	
al t	i->7	r->3	y->1	
al u	n->1	p->1	t->11	
al v	a->2	e->2	
al ä	n->1	r->6	
al å	k->1	s->1	t->1	
al ö	v->3	
al!H	ä->1	
al" 	m->1	o->1	
al, 	T->1	a->2	d->2	e->1	g->1	h->2	l->1	m->1	n->1	o->6	r->1	s->2	t->1	v->2	
al- 	o->7	
al-F	i->3	
al-S	h->1	
al-s	o->2	
al. 	J->1	
al.D	e->5	
al.E	n->1	
al.F	r->1	ö->4	
al.H	e->2	u->1	
al.I	 ->1	n->1	
al.J	a->2	
al.K	a->1	o->1	
al.M	e->1	
al.P	e->1	
al.S	a->1	j->1	t->1	å->1	
al.V	i->3	
al: 	O->1	p->1	
al; 	a->1	
alFi	n->1	
ala 	E->1	K->1	a->8	b->9	d->10	e->18	f->13	g->7	h->3	i->10	j->1	k->9	l->6	m->36	n->1	o->84	p->22	r->7	s->50	t->4	u->19	v->7	ä->2	å->3	ö->1	
ala"	;->1	
ala,	 ->5	
ala.	D->4	I->1	J->1	K->1	S->1	
ala?	D->3	
alac	i->15	
alad	 ->1	e->34	
alaf	r->1	
alag	 ->3	,->1	e->1	
alai	 ->7	
alam	,->1	
alan	 ->2	.->2	d->52	g->1	k->1	s->35	
alar	 ->69	,->2	.->4	?->1	e->30	n->13	s->1	t->2	
alas	 ->10	,->1	i->6	
alat	 ->20	,->3	.->2	e->1	l->1	s->6	
alay	a->1	
alba	n->18	r->1	
albe	l->1	s->2	
albl	o->1	
ald 	f->4	i->2	k->1	p->2	r->1	ä->1	
ald,	 ->6	
ald.	J->1	
alda	 ->13	,->1	?->1	g->1	
alde	 ->2	l->3	m->16	n->5	s->3	z->3	
aldi	g->2	r->17	s->1	
aldj	u->1	
aldo	m->1	
aldr	i->31	
alei	d->2	
alej	d->1	
alek	o->4	
alem	 ->2	
alen	 ->21	,->3	.->3	?->1	s->1	t->1	
aleo	t->1	
aler	 ->11	,->1	.->3	m->1	n->5	
ales	 ->8	.->2	;->1	a->1	e->1	m->2	t->22	ä->2	
alet	 ->53	,->11	.->5	s->3	
aleu	r->1	
alfa	b->1	
alfo	n->15	r->3	
alfr	a->3	i->2	å->5	
alfå	n->4	
alfö	r->11	
alib	e->1	i->1	
alic	i->2	
alie	n->36	r->4	s->1	
alif	i->15	
alig	 ->2	a->2	t->1	
alin	a->1	i->2	r->1	
alis	e->64	k->5	m->11	t->66	
alit	a->8	e->50	i->14	
alj 	o->1	ö->1	
alj,	 ->2	
alj.	V->1	
alja	n->1	
alje	r->26	
aljf	l->1	
aljk	o->2	
alka	n->7	
alke	m->1	
alko	h->1	r->1	
alkr	e->4	
all 	7->1	E->2	K->1	a->37	b->78	c->3	d->34	e->9	f->67	g->52	h->46	i->50	j->14	k->82	l->23	m->18	n->7	o->21	p->12	r->12	s->66	t->38	u->32	v->64	ä->11	å->10	ö->11	
all"	,->1	
all,	 ->12	
all.	 ->2	B->1	D->4	E->1	H->1	J->3	M->1	S->1	V->2	
alla	 ->357	!->1	,->5	.->4	d->10	n->6	r->7	s->6	t->5	
alld	e->23	
alle	g->1	h->3	l->10	n->9	r->45	s->5	t->56	u->2	
allf	ä->1	
alli	a->7	b->1	e->1	h->1	n->1	t->4	
allk	l->2	
allm	o->1	ä->121	ö->1	
allo	k->1	
allp	o->1	
allr	a->9	i->1	
alls	 ->14	,->1	.->2	f->1	h->1	i->1	m->1	s->3	t->5	ä->1	
allt	 ->173	,->7	.->6	:->1	f->39	i->83	j->3	m->1	s->63	
allv	a->74	
ally	 ->1	!->1	.->1	b->1	s->1	
alma	n->427	
alme	d->1	
alna	 ->1	
alni	n->15	
alog	 ->17	,->1	.->7	e->8	
alpa	r->1	t->1	
alpo	l->44	
alpr	o->2	
alre	s->4	
alri	k->4	
alrä	k->1	
als 	a->2	b->1	f->4	g->1	h->1	i->2	k->1	m->5	o->4	p->2	s->2	å->2	
als.	D->1	
alse	k->2	
alsf	a->1	
alsk	a->5	n->1	o->1	t->1	u->1	
alsl	ö->1	
also	c->1	
alsp	a->1	u->6	
alsr	u->1	
alss	t->1	
alst	a->3	ö->2	
alsu	m->1	
alsy	s->1	
alt 	2->1	7->1	9->1	E->1	a->8	b->1	d->1	f->2	h->5	i->9	m->1	n->1	o->4	p->4	r->3	s->9	t->2	u->3	v->2	ä->2	
alt,	 ->5	
alt.	D->2	J->1	O->1	V->2	
alta	 ->6	,->1	k->1	r->2	s->1	
alte	r->13	s->3	
alti	d->1	
altn	i->47	
alts	 ->4	.->1	
aluf	ö->1	
alun	d->3	
alut	a->23	b->2	
alv 	d->1	m->1	t->2	
alva	 ->4	
alve	r->1	
alvh	j->1	
alvi	n->1	
alvm	i->1	
alvo	f->1	l->1	
alvt	 ->2	i->3	
alvv	ä->2	
alvå	r->5	
alvö	,->1	.->1	n->1	
alyd	a->1	e->2	
alys	 ->26	,->4	.->5	?->2	a->2	e->21	
alös	a->1	
am "	K->1	
am -	 ->5	
am 1	9->1	
am 8	0->1	
am D	e->1	
am a	c->1	l->1	r->1	s->2	v->5	
am b	e->5	l->1	u->1	
am c	o->1	
am d	a->1	e->21	i->2	
am e	f->1	m->17	n->15	r->1	t->23	u->2	
am f	l->1	o->1	r->1	ö->45	
am g	e->1	r->1	ö->2	
am h	a->4	e->1	ä->4	å->1	
am i	 ->13	n->5	
am k	a->1	o->2	v->1	
am l	a->2	i->1	ä->1	ö->2	
am m	a->2	e->10	i->1	o->1	y->1	å->4	
am n	i->1	o->1	u->1	ä->2	å->2	
am o	c->9	m->6	
am p	o->1	r->1	å->10	
am r	a->1	e->8	i->1	ä->1	
am s	a->4	i->3	k->4	l->1	o->12	p->1	t->7	y->2	ä->3	å->2	
am t	a->1	i->47	r->3	
am u	n->1	t->3	
am v	a->4	e->2	i->3	å->2	
am ä	n->2	r->2	v->1	
am å	k->1	s->1	t->1	
am ö	k->1	v->3	
am!D	e->1	
am, 	K->1	a->2	b->2	d->3	e->1	f->2	i->1	j->1	m->2	n->1	o->7	p->1	r->1	s->7	u->2	v->2	
am..	(->1	
am.D	e->5	
am.F	r->3	ö->1	
am.G	e->1	ö->1	
am.H	e->1	u->1	
am.I	 ->1	
am.J	a->2	
am.K	o->1	u->1	
am.M	e->2	
am.N	a->1	ä->1	
am.O	m->1	
am.R	e->1	
am.S	l->1	t->1	y->1	
am.T	i->1	
am.V	i->2	
am?J	a->1	
am?V	i->1	
ama 	-->1	h->1	o->1	p->1	s->1	u->1	
ama.	J->1	V->1	
amaf	f->1	
aman	s->1	
amar	 ->2	,->3	.->1	b->83	n->2	
amas	 ->2	k->1	
amat	i->6	
amav	t->3	
amba	l->1	n->47	s->1	
ambi	t->26	
ambu	l->1	r->2	
ame-	f->1	
amel	s->1	
amen	 ->60	,->4	s->2	t->609	
amer	 ->41	a->2	i->15	
amet	e->1	r->1	
amex	i->2	
amfa	r->1	
amfi	n->1	
amfu	n->5	
amfö	r->179	
amgi	c->1	
amgå	 ->1	n->38	r->12	t->1	
amhe	t->97	
amhä	l->49	r->1	v->4	
amhå	l->17	
amhö	l->2	
amid	i->1	
amik	 ->1	
amil	j->15	
amin	a->2	e->10	g->8	i->1	
amis	k->4	
amka	r->1	s->1	t->2	
amko	m->10	
amla	 ->38	d->2	g->12	r->3	s->1	t->5	
amle	v->1	
amli	g->2	n->25	
amlä	g->8	
amm 	a->1	
amma	 ->255	,->4	.->2	d->1	l->4	n->250	r->68	s->2	t->4	
amme	 ->2	n->36	r->22	t->73	
amn 	K->1	b->1	i->1	k->1	m->3	o->1	p->1	s->2	
amn,	 ->2	
amn.	D->1	M->1	V->1	
amna	 ->3	d->1	r->22	v->2	
amnb	e->1	
amne	n->2	t->2	
amni	n->3	
amnk	o->2	
amnu	p->4	
amo,	 ->1	
amod	 ->2	
amor	d->38	
amot	 ->25	!->7	,->16	e->26	
amp 	J->1	f->2	i->3	m->5	
ampa	g->1	n->6	
ampe	n->16	r->3	
ampl	a->8	
ampo	r->1	
ampr	o->12	
ampå	l->1	
amra	t->1	
amre	 ->1	s->1	
amru	n->1	
amrä	t->1	
amrå	d->9	
ams 	B->1	
amsk	j->1	r->1	y->4	
amst	e->32	ä->14	å->5	ö->1	
amsy	n->3	
amt 	G->1	H->1	a->12	b->4	d->2	e->7	f->12	h->1	i->3	j->1	k->5	l->3	m->5	n->1	o->9	p->2	r->6	s->7	t->4	u->8	v->1	y->1	ä->3	å->1	ö->1	
amt,	 ->2	
amt.	P->1	U->1	Å->1	
amta	g->5	l->16	
amti	d->174	
amtl	i->25	
amtr	ä->2	
amtv	i->2	
amty	c->6	
amus	 ->1	
amut	f->1	
amve	r->4	t->2	
amvi	l->3	
amål	 ->1	,->2	.->2	e->6	s->2	
amåt	 ->12	,->3	.->7	
amöt	e->84	
amöv	e->2	
an "	e->1	
an -	 ->6	
an 1	0->2	5->1	7->1	9->22	
an 4	 ->1	
an 8	 ->2	
an A	l->1	m->1	
an B	r->2	
an C	E->1	e->1	
an D	a->3	e->1	
an E	G->1	K->1	M->1	U->1	r->1	u->13	
an F	l->1	o->1	
an G	a->1	o->1	
an H	a->2	u->23	
an I	m->2	s->11	
an J	u->1	
an K	o->2	
an L	a->1	
an N	i->1	
an P	a->1	l->1	o->2	r->1	
an R	o->1	
an S	P->1	c->1	e->1	h->1	y->2	
an V	e->1	
an W	i->3	
an a	 ->1	b->1	c->10	g->2	k->1	l->12	m->1	n->41	p->1	r->8	t->102	v->33	
an b	a->13	e->50	i->10	l->12	o->6	r->2	y->2	ä->2	ö->20	
an c	e->2	h->1	
an d	a->3	e->140	i->6	o->3	r->9	y->1	ä->13	å->9	ö->3	
an e	f->7	k->3	l->4	m->7	n->43	r->10	t->10	x->4	
an f	a->13	e->1	i->15	l->5	o->12	r->31	u->4	y->3	ä->2	å->20	ö->102	
an g	a->10	e->28	i->1	j->3	l->1	o->10	r->4	ä->5	å->12	ö->36	
an h	a->115	e->7	i->7	j->5	o->4	u->5	ä->21	å->1	ö->3	
an i	 ->83	b->1	d->3	f->2	g->1	n->153	s->2	t->1	
an j	a->42	u->7	ä->2	
an k	a->45	l->3	n->1	o->70	r->8	u->6	v->7	y->1	ä->1	ö->4	
an l	a->6	e->12	i->5	o->4	y->7	ä->22	å->2	ö->5	
an m	a->34	e->48	i->4	o->6	y->7	ä->2	å->42	ö->3	
an n	a->10	i->9	o->3	u->14	y->3	ä->11	å->14	ö->1	
an o	c->107	f->2	l->3	m->125	p->2	r->7	s->1	v->2	
an p	a->6	e->2	l->3	o->6	r->8	u->1	å->53	
an r	a->3	e->36	i->9	o->1	u->1	ä->5	å->5	ö->7	
an s	a->32	e->17	i->13	j->1	k->77	l->6	n->9	o->20	p->6	t->33	v->3	y->3	ä->23	å->6	
an t	a->48	e->3	i->50	j->2	o->1	r->5	v->35	y->5	ä->5	
an u	n->21	p->31	r->3	t->38	
an v	a->42	e->19	i->102	o->1	r->1	ä->11	å->1	
an y	t->2	
an Ö	s->1	
an ä	g->7	n->7	r->74	v->15	
an å	 ->2	r->3	s->5	t->13	
an ö	k->1	n->1	p->2	v->19	
an! 	A->5	B->2	D->33	E->5	F->12	G->2	H->1	I->10	J->74	K->5	L->6	M->5	N->5	O->2	P->4	R->4	S->9	T->8	U->4	V->17	Ä->7	Å->3	Ö->1	
an!A	m->1	
an!D	e->2	
an!E	f->1	n->1	
an!J	a->6	
an!M	i->1	
an!S	a->1	
an!T	a->1	i->1	
an!U	n->1	
an!V	i->2	
an" 	a->1	g->1	
an",	 ->1	
an".	R->1	
an, 	K->2	U->1	a->12	b->2	d->10	e->9	f->26	g->3	h->42	i->6	j->4	k->34	m->20	n->7	o->12	p->5	r->1	s->17	t->4	u->7	v->9	ä->14	
an- 	o->1	
an-C	l->1	
an-K	e->1	
an. 	D->1	
an.(	L->1	P->2	
an.)	 ->1	
an.A	l->1	v->1	
an.D	e->16	ä->2	å->1	
an.E	f->1	n->1	
an.F	r->1	ö->4	
an.H	e->3	u->2	
an.I	 ->2	l->1	n->1	
an.J	a->14	
an.K	o->3	
an.L	å->1	
an.M	e->3	
an.N	i->1	ä->1	
an.O	c->1	
an.S	e->1	k->1	l->2	o->1	å->3	
an.T	a->1	y->1	
an.U	n->2	t->1	
an.V	a->3	i->4	å->2	
an: 	A->1	K->1	V->2	n->2	v->1	
an; 	J->1	d->1	s->1	
an? 	2->1	
an?F	r->1	
an?H	e->1	u->1	
an?J	a->1	
an?O	m->1	
an?S	e->1	
an?V	e->1	
an?Ä	r->1	
anNä	s->1	
ana 	-->2	E->1	M->1	T->1	a->4	b->4	d->10	e->3	f->10	g->2	h->5	i->2	k->1	l->1	m->2	o->3	p->5	r->5	s->9	t->1	v->2	å->2	
ana,	 ->2	
anad	a->2	e->4	
anal	,->1	.->2	e->4	f->1	i->3	y->58	
anam	m->4	
anan	d->1	e->1	
anar	 ->31	,->1	
anas	 ->4	
anat	 ->4	i->1	
anbe	r->2	
anbi	l->8	n->1	
anbl	a->2	i->1	
anbo	e->1	
anbr	o->1	y->1	
anbu	d->4	l->1	n->1	
anc,	 ->1	
anca	,->1	s->1	
ance	,->1	.->1	r->3	
anci	s->1	
and 	-->4	8->1	E->1	S->1	T->1	a->31	b->7	d->20	e->6	f->5	g->4	h->11	i->17	k->6	l->3	m->55	n->6	o->36	p->5	r->2	s->36	t->9	u->6	v->9	ä->14	ö->1	
and)	,->1	
and,	 ->35	
and.	A->1	D->6	E->1	G->1	I->6	J->6	K->1	L->1	M->2	N->2	O->2	S->1	U->1	V->1	Å->1	
and?	F->1	
anda	 ->16	,->5	.->5	d->9	h->43	l->9	m->1	n->4	r->27	s->1	t->24	
ande	 ->1434	!->9	(->1	,->101	.->115	:->15	;->3	?->4	b->2	f->11	h->1	k->9	l->45	m->5	n->251	r->15	s->115	t->386	v->2	
andf	u->1	
andi	c->1	d->14	e->1	g->2	k->4	n->1	s->1	
andl	a->172	i->187	ä->1	
andm	ä->1	
andn	i->10	
ando	m->14	
andr	a->336	e->1	i->7	
ands	 ->11	,->1	a->4	b->44	k->14	m->9	p->3	v->1	ä->1	
andu	p->2	t->1	
andv	i->2	
andz	i->4	
ane 	o->2	
ane,	 ->1	
anel	e->1	
anen	 ->16	,->2	.->7	s->2	t->8	
aner	 ->22	"->1	,->2	.->4	a->37	i->20	n->22	
anes	i->1	
anet	 ->3	,->2	.->2	
anfa	l->2	t->12	
anfl	y->1	
anfö	r->50	
ang 	a->1	b->1	e->1	f->4	g->2	h->3	i->1	j->1	k->1	m->2	n->1	o->4	s->5	u->1	ä->4	
ang,	 ->8	
ang.	.->1	D->4	E->1	H->1	J->2	O->2	Ä->1	
anga	v->1	
ange	 ->15	,->1	l->22	m->4	n->21	r->8	s->9	t->12	
angi	v->5	
angr	e->6	i->7	ä->1	
angå	e->26	r->2	
anha	n->47	
anhe	d->2	
anhä	n->5	
anhå	l->54	
anhö	j->4	
ani 	s->1	
ani,	 ->4	
anie	n->9	
anif	e->1	r->1	
anik	 ->1	
anin	e->1	g->33	v->1	
anio	;->1	
anis	a->43	e->18	m->11	t->2	
anit	e->1	ä->1	
aniu	m->2	
aniv	å->1	
anj 	f->2	m->1	
anj.	D->1	
anje	n->1	r->1	
anjo	r->1	
anjä	m->1	
ank 	e->1	v->1	
ank"	 ->1	
ank-	 ->1	
anka	 ->2	.->1	l->9	r->17	
anke	 ->48	,->2	b->1	f->1	g->1	n->24	p->1	r->8	s->1	
ankf	a->7	o->1	ö->1	
anki	r->1	
ankl	a->4	
ankn	y->1	
anko	.->1	m->3	p->1	
ankr	a->9	e->2	i->39	
anks	c->1	e->1	
ankt	 ->1	i->8	
anla	g->1	
anle	d->50	
anli	g->15	t->1	
anlä	g->13	n->2	
anlö	p->4	
anma	n->1	r->26	
anmä	l->19	r->10	
ann 	d->1	e->1	o->1	t->1	ä->1	
ann,	 ->1	
ann-	g->1	
anna	 ->8	b->1	k->2	l->1	n->44	r->20	t->72	
anne	n->25	r->4	s->1	
annh	e->1	
anni	e->14	n->10	v->1	
annl	a->1	y->1	ä->1	
anno	l->9	r->4	
anns	 ->14	a->1	k->1	
annä	m->2	
ano 	P->2	o->1	u->1	
anoi	s->1	
anon	 ->2	,->1	.->1	?->1	e->1	y->4	
anor	.->4	d->9	
anos	 ->1	!->1	
anpa	s->14	
anpå	 ->1	
anrö	j->6	
ans 	-->1	H->1	a->18	b->16	d->3	e->5	f->21	g->3	h->2	i->8	k->7	l->4	m->31	n->1	o->9	p->6	r->1	s->15	t->1	u->9	v->5	ä->1	å->1	
ans,	 ->18	
ans.	D->2	E->1	L->1	M->1	
ans;	 ->1	
ans?	.->1	
ansa	t->10	
ansc	h->7	
ansd	e->1	
anse	 ->1	.->1	e->2	n->23	r->215	s->5	t->2	u->1	
ansi	e->78	k->1	n->1	o->1	t->7	ä->1	
ansj	o->17	
ansk	 ->7	a->139	e->65	l->1	n->23	o->9	r->1	t->6	u->1	
ansl	a->23	e->1	i->1	o->1	u->29	å->5	
ansm	i->1	ä->6	
ansp	e->1	o->108	r->7	
ansr	ä->22	
anst	a->8	o->2	r->46	ä->38	å->1	
ansv	a->306	ä->11	
ansä	t->5	
anså	g->12	t->1	
ansö	k->10	v->1	
ant 	-->3	E->2	a->12	b->3	c->1	d->4	f->17	g->1	h->2	i->5	k->4	m->1	n->3	o->5	p->4	s->24	t->3	u->2	ä->2	ö->1	
ant!	"->1	
ant,	 ->7	
ant.	D->2	H->1	S->1	V->1	
ant:	 ->1	
anta	 ->36	b->3	g->71	l->58	r->9	s->24	t->1	
ante	 ->3	,->2	n->9	r->114	
anti	 ->9	,->1	-->3	.->1	b->1	d->1	e->18	f->10	k->4	m->1	n->14	q->1	s->12	t->5	
antk	u->1	
antl	i->3	
antn	i->1	
anto	g->23	r->1	
antr	a->3	ä->35	
antv	e->2	
anty	d->2	
antö	r->3	
anua	r->16	
anut	s->1	
anva	p->4	
anvi	s->1	
anvä	n->184	
anyo	n->3	
anz 	F->3	
anze	s->1	
anço	i->1	
anös	t->19	
anöv	r->1	
ao t	i->1	
aord	i->1	
aos 	n->1	o->1	
ap -	 ->1	
ap a	t->2	v->20	
ap b	ö->2	
ap d	e->1	ä->2	
ap e	l->1	
ap f	r->1	ö->2	
ap g	r->1	
ap h	a->1	
ap i	 ->5	n->2	
ap k	o->1	
ap m	e->1	å->1	
ap n	ä->1	
ap o	c->12	m->3	
ap s	k->2	o->9	
ap t	i->1	
ap u	n->1	p->1	
ap v	a->1	
ap ä	r->1	
ap" 	f->1	
ap"!	I->1	
ap",	 ->1	
ap, 	d->2	e->3	f->2	h->1	i->1	o->3	u->1	v->2	ä->1	
ap. 	S->1	
ap.D	a->1	e->6	
ap.E	u->1	
ap.I	 ->2	
ap.J	a->2	
ap.S	l->1	
ap.T	i->1	
ap.V	i->2	
ap: 	K->1	
apa 	O->1	a->2	b->3	d->4	e->39	f->8	g->1	h->3	i->3	j->1	k->5	l->1	n->8	o->2	r->1	s->9	t->6	v->1	y->1	ä->1	
apac	i->5	
apad	e->5	
apan	 ->2	,->1	d->24	s->1	
apar	 ->25	.->2	e->2	l->166	
apas	 ->13	
apat	 ->7	.->1	s->2	
apay	a->2	
apea	u->1	
apen	 ->54	,->10	.->11	?->1	h->1	i->1	s->72	t->1	u->1	
aper	 ->4	,->1	.->1	i->1	n->16	
apes	t->1	
apet	 ->61	)->1	,->13	.->6	?->1	s->15	
apit	a->27	e->6	u->2	
apka	y->11	
apla	n->1	
apli	g->37	
apne	n->2	
apol	i->2	
app 	d->1	h->1	u->1	
app,	 ->1	
app.	V->1	
appa	 ->4	d->3	r->3	s->9	
appe	l->1	n->1	r->8	
apph	e->3	
appj	a->1	
appl	a->2	å->6	
appn	i->1	
appo	r->112	
apps	s->1	
appt	 ->5	
appv	e->2	
appy	 ->1	
apri	l->3	
apro	b->1	c->2	d->1	j->1	p->1	
aps 	f->1	
aps-	 ->1	
apsa	v->2	
apsb	e->3	
apsd	i->1	
apsf	r->1	
apsi	n->14	
apsk	o->3	
apsl	a->3	
apsm	a->2	e->1	ä->16	å->1	
apsn	i->11	
apso	r->1	
apsp	e->2	o->2	r->3	
apsr	a->1	e->9	ä->8	
apss	t->3	y->1	
apså	t->2	
apte	n->2	
ar "	ö->1	
ar (	C->2	F->1	
ar -	 ->13	
ar 1	,->1	0->1	3->1	5->2	7->1	9->3	
ar 2	6->1	
ar 3	-->1	
ar 4	0->1	
ar 9	7->1	
ar A	l->2	
ar B	N->1	r->2	
ar C	e->1	
ar E	u->14	v->1	
ar F	l->1	ö->1	
ar G	o->1	
ar I	n->1	
ar K	u->1	
ar L	a->1	o->2	y->1	
ar P	a->1	o->1	r->1	
ar R	E->1	h->1	o->1	å->1	
ar S	e->1	o->1	w->1	
ar T	h->1	
ar W	a->1	
ar a	b->1	c->2	g->1	k->3	l->44	n->49	r->7	s->1	t->128	v->69	
ar b	a->11	e->63	i->11	l->21	o->1	r->9	u->1	y->4	ä->4	å->2	ö->7	
ar c	i->1	o->1	
ar d	a->1	e->302	i->11	o->7	r->9	ä->33	å->5	ö->2	
ar e	f->15	g->1	k->2	l->10	m->9	n->119	r->19	t->57	u->2	x->10	
ar f	a->16	e->2	i->6	l->10	o->6	r->54	u->8	ä->1	å->28	ö->212	
ar g	a->3	e->28	i->6	j->46	l->2	o->8	r->4	ä->3	å->14	ö->2	
ar h	a->38	e->24	i->10	j->1	o->8	u->4	ä->20	å->6	ö->14	
ar i	 ->143	.->1	a->1	d->4	f->1	g->4	h->1	n->155	s->1	t->6	v->1	
ar j	a->78	u->24	
ar k	a->13	l->6	o->84	r->7	u->15	v->3	ä->1	ö->2	
ar l	a->37	e->10	i->10	o->4	u->1	y->18	ä->18	å->3	ö->6	
ar m	a->44	e->101	i->51	o->15	y->14	ä->4	å->9	ö->8	
ar n	a->8	e->3	i->12	o->5	u->18	y->9	ä->24	å->34	ö->5	
ar o	a->2	b->1	c->154	e->1	f->6	k->1	l->5	m->138	r->12	s->24	
ar p	a->14	e->8	l->1	o->4	r->15	u->4	å->109	
ar r	a->4	e->39	i->3	y->1	ä->22	å->14	ö->10	
ar s	a->42	e->20	i->63	j->5	k->46	l->7	m->1	n->1	o->101	p->9	t->42	u->3	v->4	y->4	ä->15	å->21	
ar t	a->32	e->3	i->122	j->2	o->1	r->9	u->1	v->9	y->8	ä->2	
ar u	n->24	p->43	r->1	t->52	
ar v	a->50	e->23	i->158	u->1	ä->18	å->14	
ar y	t->2	
ar Ö	V->1	
ar ä	g->5	l->1	m->1	n->22	r->28	v->10	
ar å	 ->1	l->1	r->3	s->2	t->7	
ar ö	k->6	n->2	p->1	s->2	v->29	
ar! 	A->1	B->1	D->2	E->1	F->3	H->1	J->4	N->1	P->1	S->2	T->1	V->1	
ar!D	e->1	
ar!J	a->1	
ar!M	e->1	i->1	
ar!T	i->1	
ar" 	m->1	o->1	
ar).	)->1	
ar, 	P->1	T->1	W->1	a->12	b->3	d->13	e->9	f->13	g->2	h->2	i->10	j->5	k->14	l->8	m->18	n->5	o->38	p->4	r->1	s->20	t->3	u->10	v->10	ä->9	å->3	
ar- 	s->1	
ar. 	A->1	E->1	M->1	V->1	
ar.)	S->1	
ar.-	 ->1	
ar..	 ->2	.->1	
ar.A	m->1	t->1	
ar.B	a->1	e->1	l->1	o->1	
ar.D	e->59	ä->4	å->1	
ar.E	f->2	n->2	r->1	u->2	
ar.F	P->1	r->1	ö->14	
ar.G	e->2	ö->1	
ar.H	e->7	u->1	ä->1	
ar.I	 ->10	n->4	
ar.J	a->32	
ar.K	o->3	r->1	
ar.L	i->1	å->2	
ar.M	a->2	e->8	i->1	
ar.N	a->1	i->1	å->1	
ar.O	b->1	c->2	m->6	
ar.P	å->2	
ar.R	e->1	i->1	ä->1	å->1	
ar.S	e->2	k->1	o->1	t->1	å->2	
ar.T	a->2	i->3	
ar.U	n->1	t->1	
ar.V	a->1	i->28	å->1	
ar.Ä	n->2	
ar: 	D->1	F->1	P->1	a->2	d->3	f->1	o->1	u->1	v->2	
ar; 	i->2	m->1	o->1	
ar?I	 ->1	
ar?J	a->1	
ar?K	a->1	o->1	
ar?N	a->1	i->1	
ara 	"->2	1->3	2->1	5->1	7->1	B->1	D->1	E->2	I->1	a->42	b->25	c->2	d->32	e->115	f->63	g->17	h->20	i->22	j->4	k->26	l->18	m->59	n->33	o->30	p->19	r->13	s->56	t->32	u->19	v->31	y->3	Ö->1	ä->18	å->3	ö->7	
ara"	.->1	
ara,	 ->7	
ara.	A->2	D->2	F->1	J->2	M->1	P->1	V->1	
ara:	 ->2	
ara?	D->1	
arab	i->6	l->1	s->2	
arad	 ->2	e->15	o->6	
arag	r->3	
arak	 ->5	.->1	s->3	t->15	
aral	l->5	
aram	e->2	
aran	 ->3	.->1	d->287	n->1	s->6	t->93	
arar	 ->67	,->1	e->26	
aras	 ->11	t->13	
arat	 ->8	e->1	i->1	s->4	
arav	 ->4	
arba	r->2	s->1	
arbe	t->564	
arce	l->2	
arco	u->1	
ard 	C->1	K->1	e->1	f->1	o->1	p->1	s->2	v->1	
ard,	 ->3	
ard-	a->1	
ard.	D->1	
ard;	 ->1	
arda	g->4	
arde	-->1	m->1	n->3	r->19	
ardi	s->9	
are 	-->3	1->2	2->1	3->1	4->1	D->2	E->2	a->39	b->30	d->14	e->22	f->91	g->9	h->26	i->47	j->1	k->34	l->3	m->21	n->11	o->43	p->23	r->10	s->75	t->31	u->12	v->10	ä->31	å->5	ö->2	
are!	S->1	
are"	 ->2	,->1	
are,	 ->77	
are.	 ->3	A->2	B->1	D->19	E->4	F->2	H->1	I->3	J->6	K->2	M->6	N->1	P->1	R->1	S->2	T->2	U->1	V->6	Ä->4	
are:	 ->1	
are?	D->1	K->1	O->1	
areb	e->3	
aref	t->1	
arel	a->1	ä->2	
arem	s->2	
aren	 ->77	)->2	,->17	.->23	;->1	?->1	d->2	h->24	s->5	t->1	
arep	r->1	
arer	 ->15	,->3	.->2	a->4	n->1	
ares	 ->17	,->3	
aret	 ->54	,->2	.->16	
areu	r->1	t->4	
arfo	r->1	
arfä	r->1	
arfö	r->52	
arga	 ->1	n->5	r->2	
argi	n->6	
argo	 ->1	t->1	
argu	m->17	
argö	r->17	
arhe	t->21	
arhu	s->1	
arhä	n->1	
arhå	g->2	l->2	
ari 	1->4	2->5	e->2	f->1	i->3	m->1	n->1	o->3	
ari!	H->1	
ari,	 ->10	
ari.	H->1	V->1	
aria	 ->1	t->2	
aric	i->1	
arie	 ->1	n->1	r->3	t->1	
arig	 ->18	,->3	a->29	e->1	h->5	t->6	
arik	e->24	
arin	 ->1	g->27	h->6	n->1	
ario	 ->1	r->1	t->2	
aris	 ->1	,->1	e->3	f->1	k->18	m->6	t->2	
arit	 ->73	e->53	i->3	
ariu	m->2	
arje	 ->91	
ark 	-->1	b->1	e->3	f->2	h->1	i->3	k->4	l->1	m->1	o->6	p->4	s->5	t->3	v->3	
ark,	 ->4	
ark.	D->2	F->1	J->1	
arka	 ->13	,->1	n->3	r->7	s->7	
arkb	o->1	
arke	 ->1	n->20	r->10	t->1	
arki	.->1	n->2	s->1	v->2	
arkl	a->1	
arkn	a->191	
arko	l->1	m->1	n->3	t->7	v->1	
arks	 ->2	
arkt	 ->21	,->1	.->1	
arl 	H->1	v->3	
arl-	H->1	
arla	g->3	m->600	n->3	
arle	d->1	
arli	g->134	k->1	
arls	r->2	
arlä	g->2	k->1	n->7	
arlø	n->2	
arm 	e->4	
arm-	e->1	
arma	 ->3	c->1	d->4	k->1	n->1	t->6	
armo	d->1	n->18	
armr	a->2	
arms	i->2	t->1	
armt	 ->12	
army	n->14	
armé	 ->1	n->2	
arn 	-->1	i->1	k->1	o->2	s->3	
arn,	 ->3	
arna	 ->354	!->1	"->2	,->43	.->63	?->3	d->1	g->1	r->3	s->66	
arnb	a->1	
arnh	i->1	
arni	e->14	n->7	
arnp	o->2	
arns	 ->1	
aro 	-->1	i->1	n->1	v->1	
aro,	 ->1	
aron	 ->2	,->1	
aror	 ->3	,->1	.->2	
arou	k->1	
arpa	r->1	
arpe	g->1	
arpo	l->1	
arpt	 ->2	
arr 	i->1	
arra	n->6	
arre	s->2	
arri	s->1	ä->4	
arro	g->2	
ars 	1->1	2->1	E->1	a->1	b->3	d->1	e->2	f->6	g->2	h->4	i->4	k->5	l->1	m->3	n->2	o->4	p->2	r->2	s->6	t->2	u->4	v->1	ä->2	å->1	
ars,	 ->4	
ars.	D->1	N->1	V->1	
arsa	m->6	v->1	
arsb	e->2	u->1	
arsc	h->1	
arse	i->1	
arsf	r->47	u->4	ö->4	
arsk	a->9	u->1	ä->3	
arsl	a->1	
arsm	a->1	e->1	i->1	
arso	m->6	r->1	t->1	
arsp	o->5	
arst	a->2	i->1	o->1	å->7	
arsy	d->1	
art 	-->3	E->2	a->58	b->5	d->2	e->4	f->25	g->3	h->6	i->12	k->5	l->2	m->8	n->2	o->15	p->4	r->1	s->31	t->5	u->3	v->2	Ö->1	ä->4	
art!	H->1	
art,	 ->8	
art.	 ->1	A->1	D->1	F->2	H->1	I->1	J->1	K->2	M->1	S->1	V->3	Ä->1	
art:	 ->1	
arta	 ->7	d->3	n->3	r->2	s->2	t->2	
arte	c->4	l->15	m->9	n->8	r->25	x->3	
arth	y->1	
arti	 ->23	,->7	.->4	d->2	e->42	f->2	g->1	i->1	k->108	l->1	n->1	p->2	s->5	
artl	ä->1	
artn	e->28	
arto	n->1	
artp	l->1	
artr	a->2	
arts	i->1	m->2	o->2	s->3	
arty	g->69	
arv 	o->1	
arv,	 ->3	
arv.	"->1	B->1	E->1	
arva	t->9	
arve	n->1	r->1	t->4	
arvi	d->3	
arvl	i->1	
arvs	i->1	s->2	
arvä	r->1	
ary 	o->1	
arzw	a->1	
aräm	b->1	
aråd	a->1	e->1	
aréb	e->1	
arón	 ->2	
as -	 ->2	
as 4	0->1	
as E	u->8	
as S	j->2	
as a	g->1	l->1	n->29	r->6	t->72	u->1	v->105	x->1	
as b	e->11	i->1	l->5	o->5	r->1	ä->3	ö->1	
as c	e->5	
as d	a->6	e->23	i->4	j->1	u->1	ä->7	ö->1	
as e	f->9	g->4	k->6	l->9	n->28	t->9	v->1	x->3	
as f	a->4	i->1	l->2	o->3	r->23	u->6	å->3	ö->74	
as g	a->2	e->18	r->1	u->1	
as h	a->6	i->1	j->2	u->2	y->1	ä->5	å->3	
as i	 ->93	d->1	g->1	n->48	r->1	
as j	a->10	u->4	ä->1	
as k	a->6	l->2	o->25	r->3	u->3	v->3	ä->1	ö->1	
as l	a->5	e->9	i->6	ä->2	
as m	a->3	e->63	i->2	o->4	y->5	ä->1	å->3	ö->5	
as n	a->12	e->1	i->3	o->1	u->4	ä->9	å->9	
as o	b->1	c->65	f->7	h->1	i->2	l->5	m->18	r->6	v->1	
as p	a->3	e->2	l->2	o->6	r->6	å->59	
as r	a->2	e->7	i->1	o->2	u->3	ä->14	ö->2	
as s	a->13	e->3	i->5	j->2	k->14	l->2	n->3	o->27	p->3	t->11	u->4	v->3	y->1	ä->7	å->9	ö->2	
as t	a->3	i->51	j->1	r->4	u->2	v->2	y->3	
as u	n->19	p->22	r->1	t->17	
as v	a->13	e->10	i->15	ä->9	å->2	
as y	r->1	t->3	
as ä	g->2	n->3	r->6	v->2	
as å	l->2	r->2	s->1	t->5	
as ö	d->1	g->1	m->1	n->1	p->1	r->1	v->8	
as!D	e->1	
as!E	u->1	
as!G	e->1	
as!H	e->1	
as".	J->1	
as, 	M->1	a->5	b->2	d->1	e->9	f->8	g->1	h->4	i->6	k->1	l->1	m->7	n->1	o->14	p->2	r->1	s->14	u->7	v->3	ä->1	å->1	
as. 	D->2	M->1	P->1	
as.-	 ->1	
as.A	l->1	t->1	
as.B	e->2	l->2	
as.C	e->1	
as.D	e->25	ä->5	å->1	
as.E	k->1	n->1	t->3	
as.F	l->1	r->3	ö->2	
as.G	e->2	r->1	
as.H	e->6	i->2	
as.I	 ->8	n->2	
as.J	a->8	o->1	ä->1	
as.K	o->4	
as.M	a->1	e->7	i->1	
as.N	i->1	ä->2	
as.O	m->1	
as.P	a->3	e->1	r->2	å->1	
as.R	e->1	
as.S	a->1	l->1	n->1	
as.T	a->1	i->1	
as.U	n->1	
as.V	a->3	i->16	å->1	
as.Y	t->1	
as.Ä	n->1	
as.Å	t->2	
as: 	a->1	e->1	
as; 	e->1	
as?H	a->1	
as?S	k->1	
asab	l->1	
asac	a->1	
asad	e->2	
asar	!->1	,->1	
asas	 ->1	
asat	 ->1	t->1	
asbo	u->5	
asch	e->3	h->1	
asci	s->12	
ase.	O->1	
aseb	a->1	
asen	 ->7	,->1	.->1	
aser	 ->2	,->1	.->1	a->8	n->2	
asha	t->1	
ashi	n->3	
ashu	s->1	
asia	t->2	
asie	n->5	
asif	u->1	
asil	i->1	
asin	 ->1	
asis	 ->3	,->1	m->15	t->12	
ask 	f->1	
aska	d->2	m->1	r->1	
aske	r->2	
aski	e->2	n->6	s->4	
askr	a->1	
asku	s->1	
asm 	f->1	p->1	s->1	
asma	t->1	
asmu	g->1	
asni	n->3	
asoc	h->1	
asor	,->1	
aspe	k->36	
aspi	s->1	
ass 	e->1	f->2	o->1	t->1	v->1	
assa	 ->7	d->4	g->1	k->1	n->2	r->3	s->6	v->1	
asse	-->1	n->2	r->6	
assi	f->9	g->1	o->2	s->7	v->4	
assl	a->1	
assm	e->3	
assn	i->4	
asso	c->1	n->1	r->2	
assp	e->1	
asst	 ->1	
assu	s->1	
ast 	1->1	2->1	5->1	7->1	9->1	a->10	b->2	d->6	e->12	f->11	g->5	h->2	i->13	k->10	l->2	m->11	n->6	o->7	p->5	r->3	s->6	t->16	u->5	v->13	ä->7	å->4	ö->2	
ast!	D->1	
ast,	 ->5	
ast-	 ->1	
ast.	D->1	E->1	K->1	N->1	V->1	
ast?	V->1	
asta	 ->12	d->4	n->2	r->5	s->3	t->5	
aste	 ->146	,->1	.->3	:->1	n->6	r->2	t->4	
asti	a->1	g->2	n->1	o->1	s->12	
astk	u->1	
astl	a->3	ä->2	
astn	a->1	i->7	
asto	d->1	
astr	i->6	o->91	u->15	
asts	l->21	t->51	
astu	 ->1	
astä	n->1	
astå	e->2	
asun	e->1	
asus	 ->3	
asyl	 ->4	,->2	-->1	.->3	b->1	f->2	r->2	s->6	
asäk	e->1	
asät	t->19	
aså 	e->1	h->1	s->1	v->1	
at "	K->1	e->1	
at -	 ->10	,->1	
at 3	9->1	
at 9	0->1	
at A	d->1	
at B	r->1	
at E	r->1	u->5	
at F	l->1	r->1	
at I	t->1	
at K	i->1	
at S	j->1	
at a	d->1	l->5	n->8	r->2	t->41	v->14	
at b	a->1	e->13	i->2	l->1	o->1	r->1	ö->1	
at d	e->32	i->4	o->1	r->2	ä->2	ö->1	
at e	f->2	m->3	n->23	r->4	t->12	x->1	
at f	a->7	i->3	l->2	o->2	r->12	å->6	ö->38	
at g	e->5	r->1	å->1	ö->5	
at h	a->11	e->1	i->2	o->3	u->3	ä->2	å->2	ö->3	
at i	 ->27	c->2	f->1	g->2	n->12	
at j	a->1	u->1	
at k	l->1	o->17	r->1	ö->1	
at l	a->3	e->1	i->2	ä->4	å->1	
at m	a->2	e->12	i->5	o->7	y->4	ä->1	å->5	
at n	e->1	u->1	ä->2	å->6	ö->1	
at o	c->25	l->1	m->19	r->2	s->9	
at p	a->1	r->8	å->21	
at r	e->2	ä->2	å->2	ö->2	
at s	a->2	e->1	i->34	j->2	k->4	o->21	t->9	y->2	ä->11	å->8	ö->1	
at t	a->5	i->18	r->2	ä->1	
at u	n->7	p->6	r->6	t->9	
at v	a->6	i->10	ä->3	å->3	
at y	t->1	
at ä	m->1	n->14	r->1	
at å	r->3	t->2	
at ö	k->1	v->1	
at, 	a->2	b->2	d->1	e->6	f->1	h->2	i->3	k->3	l->1	m->4	n->2	o->12	p->2	s->5	u->3	v->3	ä->3	
at. 	F->1	H->2	O->1	
at..	H->1	
at.B	e->1	i->1	
at.D	e->19	ä->3	
at.E	n->3	
at.F	P->1	ö->2	
at.G	e->1	r->1	
at.H	e->5	u->2	ä->1	
at.I	 ->5	
at.J	a->10	
at.K	o->3	u->1	
at.L	ä->1	
at.M	e->1	
at.N	i->1	
at.O	c->1	m->1	
at.P	r->1	
at.T	a->1	i->1	r->1	
at.V	a->3	i->1	
at.Ä	n->1	
at.Å	 ->1	
at.Ö	v->1	
at: 	"->1	h->1	j->1	
at; 	a->1	
at?.	(->1	
at?J	o->1	
ata 	a->1	f->6	i->1	k->1	m->2	o->8	s->4	å->1	
ata,	 ->1	
atab	a->1	
atal	 ->1	o->2	s->5	y->2	
atan	e->3	
atar	 ->1	
atas	t->89	ä->1	
atch	a->1	e->1	
ate 	c->2	
ateg	i->63	o->8	
atek	o->1	
atel	l->3	
atem	a->2	
aten	 ->27	,->7	.->7	s->5	
ater	 ->78	)->2	,->10	-->1	.->18	;->1	?->1	a->55	g->1	i->28	n->219	s->3	
ates	-->1	
atet	 ->45	,->4	.->5	i->1	
atfö	r->4	
ath 	h->1	n->1	o->1	
ath,	 ->1	
athi	e->2	
ati 	d->1	f->3	i->1	k->1	m->1	o->9	s->1	u->1	
ati"	 ->1	
ati,	 ->4	
ati.	D->2	E->2	F->1	H->1	I->1	K->1	M->1	
atie	n->4	r->4	
atif	i->13	r->1	
atik	,->1	e->4	
atin	 ->11	,->1	.->4	o->4	r->1	s->4	
atio	n->722	
atir	e->1	
atis	 ->4	e->5	k->134	t->9	
ativ	 ->68	,->7	.->9	;->1	a->50	b->1	e->16	f->1	i->2	r->5	t->26	
atjä	n->1	
atla	n->3	
atli	g->100	s->2	
atlä	n->10	
atny	t->1	
ato 	-->1	f->2	h->1	i->1	o->1	s->2	t->1	ö->1	
ato.	J->1	
atoa	k->1	
atob	a->1	e->1	
atog	e->2	
atol	i->4	s->3	
atom	 ->3	)->1	e->3	f->1	
aton	-->1	s->1	
ator	 ->1	,->1	b->1	e->6	i->18	l->1	n->2	s->1	
atos	 ->13	
atpe	n->1	r->9	
atpr	o->1	
atri	o->1	
ats 	-->5	E->1	S->2	a->32	b->1	d->4	e->5	f->22	g->6	h->5	i->29	k->1	l->1	m->11	n->2	o->10	p->10	r->3	s->7	t->24	u->12	v->6	ä->2	å->2	
ats,	 ->28	
ats-	 ->5	
ats.	D->12	E->3	F->1	H->2	J->2	K->2	M->1	R->1	S->1	V->1	Ä->1	
ats?	F->1	K->1	
atsa	 ->7	r->3	s->2	t->1	
atsb	a->2	
atse	n->25	r->79	
atsf	ö->1	
atsk	a->1	
atsm	a->2	i->2	
atsn	i->8	
atso	s->3	
atsp	r->1	
atss	t->22	
att 	"->1	-->8	1->3	2->1	4->1	7->1	8->1	A->3	B->5	C->1	D->3	E->90	F->5	G->1	I->6	J->3	K->2	M->2	N->1	O->3	P->3	R->3	S->3	T->16	V->1	a->210	b->309	c->1	d->1071	e->148	f->474	g->298	h->173	i->204	j->91	k->318	l->148	m->352	n->102	o->90	p->144	r->152	s->474	t->245	u->260	v->573	y->6	z->1	ä->66	å->54	ö->69	
att,	 ->22	
att.	.->1	D->7	F->2	H->2	J->1	K->1	L->2	M->3	N->1	P->2	T->1	U->1	V->2	
att:	 ->2	
att?	V->1	
attB	e->1	
atta	 ->68	.->4	c->2	d->11	n->42	r->49	s->30	t->18	v->7	
atte	 ->3	-->1	b->15	f->3	i->2	l->1	n->129	p->1	r->24	s->8	
atti	g->30	n->1	t->5	
attk	v->1	
attl	e->4	
attn	a->6	e->8	i->68	
attr	a->1	e->1	
atts	 ->2	.->1	
atue	r->2	
atul	a->6	e->31	
atum	 ->9	,->2	.->1	e->2	
atur	 ->5	,->3	-->1	.->3	a->1	e->18	f->2	k->14	l->102	n->1	o->1	v->1	
atus	 ->4	.->1	?->1	e->4	f->1	
atzi	d->2	
atäc	k->1	
atör	e->4	
atöv	e->6	
atür	k->1	
au d	u->1	
au f	ö->4	
au o	c->1	
au s	a->3	
au",	 ->1	
au, 	L->1	a->1	e->1	h->1	o->1	s->2	
au.E	t->1	
auMe	d->1	
aube	t->1	
auct	o->1	
aude	 ->1	
audr	o->1	
auen	,->1	
auer	 ->1	n->1	
aufm	a->1	
auka	s->3	
aukt	o->6	
auma	t->1	
auna	 ->1	
auni	o->3	
aure	r->1	
auro	,->1	
aus 	b->3	
auss	e->1	
ausu	l->6	
auto	m->8	p->1	
autr	e->2	
aux,	 ->1	
av "	p->1	r->2	
av -	 ->6	
av 1	4->1	9->3	
av 2	0->1	
av 4	0->1	
av 5	 ->1	4->1	
av 8	 ->1	
av A	h->2	m->2	r->1	
av B	N->6	S->1	a->2	e->8	o->1	r->2	
av C	a->1	
av D	a->2	e->1	i->2	u->1	ü->1	
av E	G->1	U->17	r->1	u->70	x->2	
av F	N->1	P->2	l->1	ö->8	
av G	a->1	e->2	r->3	
av H	a->1	e->1	i->1	
av I	s->2	
av J	a->1	e->1	o->2	
av K	i->3	o->10	u->1	
av L	a->3	i->1	ö->1	
av M	a->2	c->1	o->1	
av O	L->3	s->1	z->1	
av P	a->2	o->1	é->1	
av R	a->1	i->1	
av S	a->1	c->6	
av T	a->1	e->1	h->4	i->1	o->1	
av U	N->1	
av V	a->2	ä->1	
av W	a->1	i->1	y->1	
av a	c->1	d->2	g->1	l->32	n->26	p->2	r->39	s->1	t->64	v->9	
av b	a->2	e->38	i->14	l->3	o->3	r->10	u->8	y->2	å->2	ö->3	
av c	e->2	i->6	o->1	
av d	a->5	e->544	i->26	j->1	o->12	r->1	
av e	f->4	g->2	k->10	n->109	r->18	t->52	u->7	v->1	x->8	
av f	a->47	i->6	j->2	l->16	o->8	r->28	u->5	y->1	ä->1	å->2	ö->107	
av g	a->3	e->31	i->3	l->1	o->1	r->11	ö->1	
av h	a->11	e->7	i->5	o->1	u->8	ä->2	ö->2	
av i	 ->5	b->1	c->3	d->2	m->4	n->26	
av j	o->5	u->4	ä->2	
av k	a->10	l->4	n->1	o->109	r->5	u->5	v->5	ä->8	
av l	a->19	e->11	i->13	o->5	ä->4	å->1	ö->1	
av m	a->18	e->26	i->38	o->5	y->3	ä->7	å->7	ö->1	
av n	a->14	i->1	o->1	y->11	ä->2	å->6	ö->2	
av o	a->2	b->2	c->7	f->5	k->1	l->14	m->10	n->1	r->11	s->12	t->2	u->1	v->1	
av p	a->22	e->12	i->1	o->8	r->37	å->17	
av r	a->6	e->32	i->7	y->1	ä->12	å->12	ö->1	
av s	a->12	c->1	e->7	i->24	j->3	k->20	l->2	m->2	o->15	p->2	t->72	u->4	v->2	y->20	ä->14	å->10	
av t	a->2	e->8	i->13	j->28	o->2	r->11	u->6	v->1	y->2	ä->1	
av u	n->27	p->6	t->33	
av v	a->22	e->8	i->20	o->4	ä->19	å->24	
av y	t->5	
av Ö	s->2	
av ä	l->1	m->1	n->5	r->1	
av å	l->1	r->7	s->1	t->14	
av ö	b->1	d->1	k->4	p->4	s->2	v->3	
av, 	d->2	e->1	f->1	m->1	o->3	s->1	t->1	ä->1	
av.(	S->1	
av..	 ->1	
av.D	e->4	ä->1	
av.E	f->1	r->1	
av.J	a->1	
av.M	e->1	
av.O	L->1	
av.R	å->1	
av?V	i->1	
ava 	g->1	
aval	e->4	l->1	
avan	c->1	d->1	o->2	t->1	
avar	 ->1	.->1	a->1	e->1	n->2	s->1	
avbr	o->3	u->2	y->3	ö->6	
avde	l->8	
ave 	(->2	m->1	ä->1	
ave,	 ->1	
ave-	 ->1	p->2	
aveN	ä->1	
avec	 ->1	
aven	 ->25	,->2	.->4	:->1	
aver	a->4	e->2	i->6	y->1	
avet	 ->23	,->1	.->6	s->2	t->1	
aveu	r->1	
avfa	l->22	
avfo	l->1	
avfö	r->3	
avga	s->1	v->1	
avge	 ->3	r->5	s->1	t->1	
avgi	c->4	f->4	v->1	
avgj	o->4	
avgr	ä->4	
avgå	.->1	e->1	n->2	r->1	t->1	
avgö	r->61	
avhj	ä->2	
avhä	n->2	
avhå	l->1	
avi 	I->1	
avid	 ->3	
avie	n->1	
avis	a->4	e->4	k->1	
avkl	a->1	
avkr	ä->1	
avku	n->1	
avla	 ->4	"->2	d->1	g->1	n->1	
avle	d->2	
avli	g->1	v->1	
avlo	p->1	
avlä	g->10	
avma	t->1	
avor	i->1	
avpr	i->1	
avra	p->1	
avre	g->2	
avru	n->1	
avrä	t->1	
avs 	a->1	h->2	i->2	m->1	o->1	u->1	v->1	
avs,	 ->4	
avs.	A->1	D->1	R->1	V->1	
avs?	T->1	
avsa	k->4	t->3	
avse	 ->1	d->3	e->47	r->14	s->1	t->14	v->13	
avsf	o->1	ö->1	
avsi	d->1	k->38	
avsk	a->19	e->5	i->1	r->2	y->2	
avsl	a->2	o->2	u->60	ä->2	å->3	ö->6	
avsm	i->2	
avsn	i->4	
avso	m->1	
avsp	e->5	
avst	a->1	o->2	ä->3	å->26	
avsv	a->1	
avsä	g->1	t->4	
avt 	s->1	
avta	l->89	r->1	
avtv	i->1	
avun	d->1	
avva	k->6	
avve	c->8	r->2	
avvi	k->8	s->15	
avvä	g->3	
aw, 	s->1	
aw.M	e->1	
ax a	v->1	
ax e	f->1	
ax i	n->1	
ax-f	r->3	
axa 	e->1	u->1	
axbe	l->1	
axel	r->1	
axer	i->1	
axim	a->6	e->2	i->1	
axis	 ->5	.->2	e->1	
axla	r->1	
ay f	ö->2	
ay h	a->1	
ay, 	J->1	a->1	h->1	s->1	
ay.V	i->1	
ayDe	 ->1	
ayab	e->1	u->2	
ayag	o->4	
ayan	n->2	
aybe	t->1	
ayed	 ->2	
ayer	n->1	
ays 	b->2	d->1	
ays-	d->1	
aza 	o->1	
aza,	 ->1	
aza.	D->1	S->1	
azak	s->1	
azar	e->2	
azis	m->8	t->8	
aça 	M->5	
b Sö	d->2	
b ef	t->1	
b ha	d->1	
b hj	ä->1	
b ka	n->1	
b oc	h->3	
b sk	a->1	
b va	r->1	
b) i	n->1	
b) m	i->1	
b, e	n->1	
b, s	o->1	ä->1	
b, v	i->1	
b-om	r->1	
b.An	s->1	
b.De	t->1	
ba a	n->1	
ba b	e->1	i->1	
ba f	r->1	
ba o	c->1	s->1	
ba p	å->1	
ba r	e->1	
ba t	i->1	
ba u	p->1	
ba v	a->1	
ba å	t->1	
ba-,	 ->1	
baci	l->1	
back	-->1	n->1	
bacè	t->1	
bad 	F->1	e->1	k->1	o->1	
bada	 ->1	
bade	 ->21	.->2	s->4	
bads	 ->1	
baga	t->2	
bain	"->1	
bak 	i->1	
bak,	 ->1	
baka	 ->35	.->4	?->1	d->3	g->4	v->4	
bakd	ö->1	
bakg	r->31	
bako	m->21	
baks	 ->1	o->1	
bakt	e->1	
bakå	t->3	
bal 	n->1	
bala	 ->5	m->1	n->33	
bali	s->5	
ball	m->1	
balt	 ->1	,->1	
ban 	s->1	
ban"	 ->1	
bana	 ->1	l->3	n->1	t->1	
banb	r->1	
band	 ->49	e->4	
bane	r->5	s->1	
bani	e->1	s->1	
bank	 ->1	"->1	e->14	f->1	i->1	s->2	
bann	l->1	
bano	n->5	r->3	
bans	k->4	
bant	a->1	n->1	
bar 	d->2	e->6	f->1	g->1	h->1	k->3	m->3	n->1	o->1	p->2	r->1	s->5	t->1	u->12	v->2	
bar,	 ->1	
bar.	D->2	F->1	H->1	
bara	 ->281	,->2	.->3	:->1	
barb	a->2	
bard	e->1	
bare	 ->8	.->3	
barg	o->1	
barh	e->9	
bari	e->1	s->1	
bark	b->1	
barl	i->12	
barm	a->1	
barn	 ->6	,->3	b->1	p->2	s->1	
barr	i->2	
bart	 ->84	!->1	,->4	.->9	
baré	b->1	
bas 	a->5	f->1	h->1	i->1	o->1	p->1	
bas,	 ->1	
bas.	D->1	
basa	r->2	
base	b->1	n->5	r->8	
basi	s->4	
bask	i->4	r->1	
bass	a->1	
bast	 ->2	e->1	i->2	u->1	
basu	n->1	
bat 	F->1	e->1	f->1	
bats	 ->7	.->2	
batt	 ->53	,->9	.->21	:->1	?->1	B->1	a->1	e->83	i->1	k->1	
baxa	 ->1	
baye	r->1	
bb e	f->1	
bb h	j->1	
bb o	c->3	
bb v	a->1	
bb, 	s->1	v->1	
bba 	a->1	b->2	f->1	o->2	p->1	r->1	t->1	u->1	v->1	å->1	
bbad	e->27	
bbar	 ->4	e->11	
bbas	 ->8	t->3	
bbat	 ->3	s->9	
bbel	 ->1	s->3	t->2	v->1	
bbig	a->1	
bbla	 ->10	s->1	
bbpl	a->1	
bbt 	f->5	g->2	h->1	k->3	l->1	m->2	o->1	p->1	s->14	t->1	u->1	v->2	
bbt,	 ->3	
bbt.	J->1	M->1	O->2	T->1	V->1	
bbva	r->1	
bby,	 ->1	
bbya	r->1	
bbyb	i->1	
bbyg	r->2	
bbyi	s->2	
bbym	a->1	
bbyn	 ->3	
bbyv	e->1	
be P	r->1	
be e	r->5	
be f	r->1	
be h	e->1	o->1	
be k	o->6	
be o	m->2	
be p	a->1	
be s	t->1	
beak	t->30	
bear	b->2	
bebo	e->1	
beby	g->1	
bebå	d->1	
bedd	 ->1	
bedr	e->1	i->15	ä->35	
beds	 ->1	
bedö	m->51	
befa	r->5	t->6	
befi	n->41	
befl	ä->1	
befo	g->32	l->43	r->7	
befr	a->10	i->9	ä->1	
befä	l->1	n->1	s->10	
bega	g->4	
begr	a->1	e->13	i->21	u->2	ä->68	
begä	r->60	
begå	 ->2	r->3	s->3	t->3	
beha	g->2	n->85	
beho	v->67	
behä	f->1	
behå	l->29	
behö	l->1	r->18	v->147	
beiv	r->1	
beka	n->3	
beki	s->2	
bekl	a->42	
beko	m->1	s->1	
bekr	ä->30	
bekv	ä->15	
beky	m->16	
bekä	m->41	n->1	
bel 	H->1	P->1	e->1	i->1	l->1	n->1	o->1	r->1	u->1	
bel!	M->1	
bel,	 ->4	
bel.	D->1	V->3	Ä->1	
bela	g->4	s->10	
belg	i->8	
bell	 ->4	.->2	
belo	p->16	
bels	 ->1	k->2	
belt	 ->19	.->8	;->1	?->1	
belv	ä->1	
bely	s->4	
belä	g->7	
belö	n->2	
bema	n->2	
bemy	n->1	
bemä	r->5	
bemö	d->3	t->7	
ben 	i->1	
bene	f->5	n->1	
beng	a->1	
benh	å->1	
beni	 ->2	.->1	
bens	i->1	
benä	g->1	
benå	d->1	
beor	d->1	
ber 	1->20	V->1	a->4	d->3	e->8	f->4	h->1	i->3	j->9	k->4	l->3	m->4	n->1	o->12	r->2	s->1	v->1	
ber,	 ->13	
ber.	 ->1	D->1	E->1	J->1	N->1	S->1	
bera	d->1	l->31	
berb	a->1	
bere	d->59	t->6	
berg	 ->3	e->1	
beri	k->8	s->1	
bern	a->2	
bero	d->5	e->68	p->1	r->19	t->1	
bert	 ->2	
berv	e->1	
bery	k->1	
berä	k->4	t->31	
berö	m->2	r->42	v->1	
bes 	a->1	ä->1	
bese	g->2	
besi	k->2	t->2	
besk	a->4	e->3	r->23	y->5	
besl	u->220	ä->1	ö->1	
besp	a->5	
best	o->1	r->5	y->1	ä->165	å->53	ö->1	
besv	a->17	i->8	ä->7	
besy	n->1	
besä	t->3	
besö	k->9	r->2	
bet 	F->1	d->1	h->1	m->1	o->3	s->2	t->1	u->2	
bet"	 ->1	,->1	
bet,	 ->3	
bet-	f->1	
bet.	E->1	V->1	
bet?	J->1	
beta	 ->64	,->1	.->3	?->1	d->2	l->90	n->21	r->35	s->2	t->14	
bete	 ->116	,->11	.->29	?->3	c->4	e->3	n->9	r->2	t->51	
beth	 ->1	
betj	ä->1	
beto	n->46	
betr	a->23	y->1	ä->72	
bets	-->2	a->5	b->6	d->4	f->2	g->13	i->2	k->6	l->46	m->17	n->3	o->11	p->14	r->5	t->83	v->5	
bett	 ->3	s->2	
betu	n->1	
betv	i->3	
bety	d->122	
betä	n->268	
beun	d->3	
beva	k->6	r->22	
beve	k->1	
bevi	l->48	s->43	t->1	
bexp	l->1	
bi d	e->1	
bi n	ä->1	
bibe	h->11	
bibl	i->2	
bidr	a->108	o->3	
bief	f->2	
bifa	l->3	r->2	
biga	 ->1	
bigo	t->1	
bigå	 ->1	e->4	s->1	
biha	n->1	
bikm	e->2	
bil 	e->1	f->1	g->2	i->1	k->1	o->1	s->4	v->1	
bil,	 ->2	
bil-	 ->1	
bil.	 ->1	D->1	T->1	
bila	 ->1	g->6	r->82	t->6	
bilb	e->1	r->1	
bild	 ->4	,->1	.->2	a->28	e->7	n->66	
bile	n->7	
bili	n->29	s->11	t->27	
bilj	o->1	
bilk	o->1	y->1	ö->2	
bill	i->6	
bilm	ä->1	
bilp	a->6	r->1	
bils	 ->2	e->1	k->3	p->1	
bilt	 ->2	i->15	
bilv	r->6	
bilä	g->1	
bilå	t->1	
bin,	 ->1	
bina	t->1	
bind	a->14	e->23	
bine	t->3	
bio 	s->1	
biog	r->1	
biol	o->4	
biop	l->1	
bios	f->1	ä->2	
bise	e->1	n->1	
bisk	 ->2	-->1	a->9	
bist	å->23	
bit 	p->1	
bite	r->1	
biti	o->14	ö->12	
bitt	e->2	r->1	
bjek	t->2	
bjud	a->22	e->16	i->1	n->3	
bjöd	 ->1	s->1	
bl.a	.->27	
bla 	a->1	d->2	e->1	f->9	i->2	k->1	o->1	s->4	t->1	
bla"	.->1	
bla,	 ->1	
bla.	D->1	M->1	N->1	Ö->1	
blad	 ->1	
blam	e->1	
blan	c->1	d->99	k->2	
blar	e->2	
blas	 ->1	
blek	a->1	
blem	 ->72	,->13	.->22	:->1	;->2	?->1	a->5	e->65	o->3	
bler	 ->1	a->11	i->3	
bles	 ->1	
blev	 ->15	
bli 	-->1	2->1	a->11	b->5	d->5	e->31	f->12	g->1	h->1	j->1	k->4	l->4	m->21	n->5	o->3	p->3	r->1	s->9	t->3	v->4	ä->1	ö->2	
bli,	 ->1	
bli.	U->1	
blic	 ->1	e->4	i->1	k->24	
blig	a->14	
blik	 ->2	a->6	e->12	
blin	 ->4	.->1	d->1	k->2	t->1	
blio	t->2	
blir	 ->112	,->2	:->1	
bliv	a->1	i->26	
blix	t->1	
bloc	k->6	
blom	m->3	s->3	
blon	m->1	
blot	t->3	
blun	d->4	
bly 	å->1	
bly,	 ->2	
bly.	V->1	
blyg	s->4	
blå 	b->1	
blås	e->2	
bnin	g->1	
bo i	 ->1	
bo k	v->1	
bo v	i->1	
boar	d->1	
bock	"->1	a->1	
boda	 ->2	s->1	
boel	i->1	
boen	d->3	
bogs	e->1	
bojk	o->1	
bok 	a->1	h->1	m->1	o->7	s->3	t->1	ä->2	
bok,	 ->1	
bok.	D->1	H->1	J->1	T->1	V->1	
boke	n->36	
boks	l->1	t->1	
bol 	f->2	
bola	g->12	
boli	s->7	
boll	s->1	
bomb	 ->1	.->1	a->2	e->4	n->1	
bomu	l->1	
bon 	f->1	g->1	k->1	m->1	
bon,	 ->1	
bon.	V->1	
bond	g->2	
bonm	ö->2	
bor 	d->1	i->4	p->1	
bora	t->3	
bord	 ->3	.->1	a->3	e->70	l->1	s->1	
borg	 ->1	a->168	e->3	m->2	
borr	e->1	
bort	 ->20	,->5	.->6	a->1	f->6	o->2	p->1	s->6	
bosa	t->3	
bosn	i->2	
bost	a->1	ä->4	
bosä	t->4	
bot 	p->2	
bota	r->2	
bott	e->5	n->4	
bour	g->5	
bova	r->1	
bove	n->1	
boxn	i->1	
bpla	t->1	
bra 	a->11	b->5	d->5	e->2	f->3	i->3	j->1	m->5	n->2	o->9	s->9	t->1	u->4	v->1	ä->2	å->1	
bra!	M->1	
bra,	 ->8	
bra.	D->1	E->1	J->1	P->1	S->1	V->1	
bran	d->3	s->7	
bred	 ->4	a->6	d->2	e->1	n->4	
brei	s->1	
brep	u->1	
bret	a->1	t->6	
brev	 ->4	.->1	l->1	
brie	f->1	n->3	
brig	h->1	
brik	e->3	
brin	g->13	
bris	t->62	
brit	a->14	t->17	
bro 	m->1	o->1	
broa	r->1	
brod	e->2	
brok	i->2	
brom	e->4	s->6	
bron	-->1	
bror	,->1	
brot	h->1	t->53	u->1	
brua	r->16	
bruk	 ->9	!->1	,->9	a->17	e->20	n->1	s->23	
brun	a->1	
brut	a->1	e->2	i->2	t->1	
bryg	g->3	
bryo	s->1	
bryr	 ->2	
bryt	a->8	e->8	n->2	
brän	d->3	n->5	s->7	
bräs	c->2	
bråd	s->20	
bråk	e->1	
brås	 ->2	
bröd	.->3	
brös	t->1	
bröt	 ->5	s->2	
bser	v->2	
bsid	a->1	i->22	
bsol	u->40	
bsor	b->1	
bsta	n->4	t->2	
bstr	a->1	
bsur	d->1	t->2	
bt f	r->4	ö->1	
bt g	e->2	
bt h	å->1	
bt k	a->2	o->1	
bt l	ä->1	
bt m	å->2	
bt o	c->1	
bt p	å->1	
bt s	k->2	o->9	v->1	ä->2	
bt t	a->1	
bt u	t->1	
bt v	i->1	ä->1	
bt, 	a->1	h->1	k->1	
bt.J	a->1	
bt.M	e->1	
bt.O	m->2	
bt.T	y->1	
bt.V	i->1	
bu i	n->1	
bud 	e->1	f->5	m->9	o->4	r->1	v->1	ä->1	
bud,	 ->4	
bud.	D->2	V->1	
budd	h->1	
bude	t->9	
budg	e->106	
budo	r->1	
buds	f->3	i->3	k->10	m->10	p->1	
bugg	e->1	
bukt	e->2	
bul 	f->1	
bula	n->1	r->1	
bult	e->1	
bund	e->13	i->3	n->4	s->8	
bure	t->1	
burg	 ->4	,->4	.->1	a->1	h->1	
buri	t->1	
burn	a->1	
bus 	ä->1	
buss	a->2	
buti	k->1	o->1	
bvar	n->1	
bven	t->12	
bvär	l->1	
by, 	d->1	
byar	b->1	
bybi	l->1	
byen	s->1	
bygd	 ->2	.->2	e->31	s->10	
bygg	a->57	d->4	e->12	n->19	s->3	t->5	
bygr	u->2	
byis	t->2	
byma	s->1	
byn 	h->1	l->1	å->1	
byrå	 ->2	e->1	k->30	n->2	
byta	 ->2	
byte	 ->10	,->1	t->6	
bytt	s->1	
byve	r->1	
byxf	i->1	
bält	e->10	
bänk	e->1	
bär 	a->51	b->2	d->5	e->15	f->5	i->9	l->1	m->2	n->1	o->4	p->4	s->3	u->1	v->1	ä->1	ö->1	
bär,	 ->1	
bär.	D->1	F->1	
bära	 ->25	n->2	s->3	
bärl	i->4	
bärs	 ->2	
bäst	 ->5	a->37	
bätt	r->153	
bävn	i->10	
båda	 ->23	,->1	d->1	n->1	
både	 ->46	
båta	r->8	
båte	n->1	
bé a	v->1	
bébé	 ->1	
böck	e->3	
böde	l->1	
böje	l->1	
böjt	 ->1	
böld	 ->1	
bör 	"->1	-->1	E->3	a->10	b->8	d->16	e->5	f->18	g->12	h->6	i->14	k->7	l->6	m->24	n->4	o->6	s->10	t->6	u->12	v->29	ä->4	å->4	ö->2	
bör,	 ->1	
bör.	F->1	
böra	n->1	
börd	.->1	a->17	e->6	o->2	
börj	a->115	
börl	i->10	
börs	e->2	
böte	r->1	
c - 	o->1	
c Br	a->1	
c bl	i->1	
c bö	r->1	
c då	 ->1	
c i 	E->1	d->1	
c l'	e->1	
c os	v->1	
c se	r->1	
c", 	f->1	
c) l	i->1	
c, d	v->1	
c-di	r->1	
c-sy	s->1	
c-tr	a->1	
c. o	c->1	
c. Ä	m->1	v->1	
c.De	t->1	
c.En	 ->1	
c?At	t->1	
cCar	t->1	
cNal	l->5	
ca 3	0->1	
ca C	o->1	
ca M	o->3	
ca s	a->1	
ca, 	o->1	
ca. 	1->1	
cal 	c->1	
calv	i->1	
canc	e->2	
cann	a->1	
cant	e->1	
cao 	t->1	
cap 	ä->1	
capi	t->10	
cas 	s->1	
case	.->1	
caya	b->2	g->4	
ccep	t->89	
cces	s->5	
ce b	ö->1	
ce d	e->4	
ce f	ö->1	
ce n	a->1	
ce o	c->1	r->11	
ce t	a->2	
ce, 	D->1	
ce..	.->1	
ce.A	l->1	
ce.D	e->1	
ce.J	a->2	
ce.O	f->1	
ce.S	t->1	
cedo	 ->1	
cedu	r->1	
ceko	r->1	
cekv	a->1	
celo	n->2	
cemb	e->19	
ceme	n->2	
cemi	s->1	
cen 	m->1	
cen,	 ->1	
cena	r->5	
cene	n->1	
cenn	i->7	
cens	a->1	i->1	
cent	 ->77	,->2	.->10	a->8	e->14	i->1	r->109	s->5	
cept	 ->2	.->2	a->44	e->48	i->6	
cer!	D->1	
cer,	 ->1	
cera	 ->12	d->31	n->3	r->7	s->5	t->17	
cerb	ö->1	
ceri	n->13	
cern	e->2	
cert	i->6	
cess	 ->22	"->1	,->2	.->13	?->1	e->66	i->5	r->3	u->1	
ceut	i->1	
ch "	U->1	s->1	t->1	
ch (	A->1	
ch -	 ->3	o->3	
ch 0	 ->1	
ch 1	-->1	0->2	3->1	4->1	6->1	7->2	9->13	
ch 2	 ->1	,->1	.->1	0->3	1->3	2->1	5->1	7->1	9->1	
ch 3	.->1	0->2	3->1	4->1	5->1	:->1	
ch 4	.->1	1->2	5->4	7->1	8->2	
ch 5	 ->1	.->1	3->1	
ch 6	0->1	8->1	
ch 7	 ->4	,->2	
ch 8	 ->1	,->1	2->6	6->2	9->1	
ch 9	 ->2	2->1	4->1	
ch A	l->2	m->1	n->1	
ch B	P->1	a->1	e->1	r->2	u->1	
ch C	.->1	E->1	a->1	y->1	
ch D	a->2	e->2	
ch E	L->2	U->4	d->1	l->2	m->1	r->1	t->1	u->24	
ch F	N->1	P->1	i->2	r->11	
ch G	a->2	e->1	o->1	r->3	
ch H	e->1	i->1	u->1	
ch I	I->2	n->4	r->2	s->5	t->1	
ch J	a->1	ö->1	
ch K	a->1	i->6	o->1	u->1	
ch L	a->3	e->5	
ch M	A->1	a->3	e->1	
ch N	o->1	y->1	
ch O	L->1	n->1	
ch P	P->1	S->2	a->9	o->2	r->1	
ch R	a->3	
ch S	a->10	c->1	i->1	j->1	o->1	p->1	t->2	w->1	y->8	
ch T	a->4	s->1	u->1	y->2	
ch U	z->1	
ch V	i->1	ä->1	
ch W	y->1	
ch X	 ->1	
ch a	b->1	c->1	d->2	g->2	k->4	l->18	m->4	n->58	p->1	r->15	s->4	t->150	v->32	
ch b	a->13	e->52	i->10	l->8	o->5	r->15	u->3	y->2	ä->4	å->1	ö->6	
ch c	a->2	e->6	h->2	
ch d	a->4	e->467	i->11	j->4	o->9	r->4	u->1	y->1	ä->83	å->24	ö->1	
ch e	f->34	g->1	j->1	k->22	l->1	n->90	r->17	t->33	u->9	x->4	
ch f	a->14	e->3	i->12	l->10	o->7	r->83	u->9	y->2	ä->1	å->12	ö->168	
ch g	a->7	e->43	i->4	j->1	l->3	o->2	r->10	ä->1	å->4	ö->17	
ch h	a->44	e->54	i->1	j->4	o->11	u->15	y->2	ä->9	å->16	ö->6	
ch i	 ->74	b->3	c->2	d->5	f->1	k->1	l->1	m->2	n->142	r->1	s->2	
ch j	a->149	o->5	u->7	ä->1	
ch k	a->21	i->1	l->4	n->1	o->129	r->18	u->7	v->10	ä->6	ö->1	
ch l	a->17	e->16	i->11	j->1	o->9	u->1	y->3	ä->14	å->19	ö->2	
ch m	a->21	e->143	i->39	o->24	u->1	y->8	ä->12	å->22	ö->9	
ch n	a->11	e->8	i->9	o->5	u->11	y->13	ä->16	å->5	ö->6	
ch o	a->4	b->2	c->9	d->1	e->2	f->6	j->1	k->4	l->8	m->41	n->1	p->2	r->8	s->5	t->1	u->3	
ch p	a->25	e->9	l->3	o->17	r->32	å->29	
ch r	a->7	e->66	i->9	o->4	u->1	ä->61	å->39	ö->1	
ch s	a->43	e->29	i->10	j->6	k->30	l->24	m->2	n->4	o->134	p->9	t->61	u->5	v->12	y->16	ä->33	å->28	ö->2	
ch t	.->1	a->20	e->6	h->1	i->60	j->4	o->6	r->18	u->17	v->3	y->14	ä->3	
ch u	n->25	p->24	t->57	
ch v	a->52	e->23	i->123	ä->26	å->12	ö->1	
ch y	n->1	r->1	t->5	
ch Ö	V->1	s->6	
ch ä	g->2	n->12	r->10	v->31	
ch å	 ->4	k->1	s->3	t->29	
ch ö	k->3	m->1	n->1	p->13	r->1	s->4	v->20	
ch! 	U->1	
ch)D	e->1	
ch, 	d->1	f->3	h->1	i->1	n->1	r->1	s->4	t->1	u->1	
ch.E	f->1	
ch.J	a->1	
ch/e	l->1	
ch: 	V->1	
ch?F	r->1	
chI 	o->1	
chII	.->1	
chab	l->1	
chan	d->1	s->12	
chap	e->1	
char	a->1	d->2	t->1	
che 	B->1	
chec	k->1	
chef	 ->1	e->16	
chem	a->1	
chen	 ->4	.->1	;->1	g->10	
cher	 ->3	a->1	n->2	
chez	 ->1	
chho	f->1	
chie	l->1	
chis	t->1	
chle	r->4	
chne	r->12	
choc	k->4	
chok	l->1	
chre	y->3	
chro	e->14	
chrö	d->1	
chs 	i->1	
cht 	m->1	o->1	
cht.	D->1	
chte	r->2	
chtf	ö->3	
chti	d->1	
chul	z->3	
chwa	r->1	
chwe	i->1	
chwi	t->1	
chyr	e->1	
chör	l->1	
chüs	s->4	
cial	 ->30	-->1	a->78	b->2	d->16	f->28	i->41	p->5	t->18	u->1	
cide	n->1	
ciel	l->49	
cien	,->2	t->2	
cier	i->1	
ciet	y->1	
cifi	c->2	k->27	
cil 	-->1	
cill	 ->1	
cilo	v->1	
cine	r->1	
cio 	S->1	V->3	f->1	h->1	s->2	
cio,	 ->3	
cio.	J->1	N->1	
cio:	 ->1	
cioe	k->3	
cios	 ->2	
cip 	a->3	e->3	f->1	i->7	o->4	r->1	s->5	ä->4	
cip,	 ->3	
cip.	J->1	S->1	V->2	
cipe	n->102	r->48	s->1	
cipi	e->8	
cipl	i->14	
cips	k->1	
cirk	a->4	e->1	l->2	u->3	
cis 	W->1	a->1	d->4	e->1	f->2	h->1	i->1	l->5	p->1	s->21	v->1	
cis-	p->1	
cisa	 ->1	
cise	r->11	
cism	,->1	e->2	
cist	 ->3	e->3	i->5	
cit.	F->1	
cita	m->8	t->1	
cite	r->7	t->7	
civi	l->19	
ck -	 ->1	
ck K	i->1	
ck a	l->1	n->1	t->12	v->7	
ck b	a->2	e->1	
ck d	e->6	
ck e	f->3	j->1	m->1	n->3	t->1	
ck f	r->7	å->1	ö->21	
ck g	a->1	r->1	å->2	
ck h	a->4	u->1	ö->2	
ck i	 ->6	n->11	
ck j	a->3	u->2	
ck k	a->3	l->1	o->3	ä->1	
ck l	ä->2	
ck m	e->2	i->1	o->2	y->3	å->1	ö->1	
ck n	e->1	u->1	y->1	å->3	
ck o	c->10	s->2	
ck p	a->1	å->2	
ck s	e->1	k->2	n->1	o->3	t->3	v->1	ä->3	å->15	
ck t	i->15	v->1	ä->1	
ck u	p->1	t->1	
ck v	a->8	i->8	ä->1	
ck ä	n->1	r->1	
ck å	t->2	
ck" 	-->1	
ck, 	1->1	R->1	f->6	h->6	i->3	k->4	m->2	n->1	s->3	t->1	
ck-p	o->1	
ck. 	M->1	
ck.A	v->1	
ck.D	e->2	
ck.F	r->1	
ck.H	e->2	
ck.J	a->2	
ck.K	i->1	o->1	
ck.Ä	v->1	
cka 	A->1	G->2	K->2	L->1	P->2	S->1	a->8	d->7	e->7	f->24	h->9	i->5	k->11	l->3	m->15	n->3	o->5	p->5	r->6	s->11	t->7	u->5	v->14	ä->2	å->1	
cka"	,->1	
cka,	 ->5	
cka.	(->1	B->1	
cka?	"->1	
ckad	 ->2	.->1	e->15	i->1	
ckan	 ->23	.->1	d->21	
ckar	 ->24	s->1	
ckas	 ->23	!->1	,->3	.->1	
ckat	 ->4	s->21	
ckba	r->5	
ckbi	l->1	
ckbä	r->1	
ckde	l->8	
cke 	b->1	e->2	f->3	i->2	k->2	l->2	o->1	s->3	t->3	u->1	v->1	ö->1	
cke-	a->2	d->3	f->1	m->1	s->12	
cke.	F->1	H->1	V->1	
ckel	f->3	n->3	p->1	r->1	
cken	 ->18	.->2	s->1	
cker	 ->105	,->2	.->1	:->1	a->3	i->1	t->2	
cket	 ->445	!->1	,->22	.->5	;->1	?->1	m->1	
ckfr	i->1	
ckfö	r->7	
ckhe	e->14	t->1	
ckho	l->3	
ckit	 ->1	
ckla	 ->31	.->1	d->10	n->5	r->3	s->22	t->6	
ckle	r->4	
ckli	g->106	n->175	
ckna	 ->3	d->6	n->1	r->2	s->6	t->11	
ckne	s->1	
ckni	n->47	
ckor	 ->25	,->2	.->2	n->9	s->1	
ckos	a->1	
ckpr	o->3	
ckra	 ->5	s->1	
cks 	a->4	d->2	e->1	i->1	m->2	n->1	o->1	p->1	r->1	s->1	t->1	u->2	v->2	ö->1	
cks.	P->1	U->1	
cks;	 ->1	
cksa	m->9	
cksb	å->1	
cksc	e->1	
cksd	r->3	
cksf	a->2	
cksi	l->3	
cksk	ö->1	
ckso	n->2	
cksr	i->2	
cksv	a->1	
ckså	 ->572	,->10	.->5	
cksö	d->1	
ckt 	e->1	f->1	h->2	k->1	n->2	s->3	u->1	v->1	ä->1	
ckte	 ->17	s->5	
ckts	 ->3	!->1	
ckup	a->2	e->3	
ckvi	d->3	
ckön	s->5	
clin	g->1	
co, 	e->1	
co-a	f->1	
cob 	S->2	
comb	a->1	
comm	o->1	
comp	a->1	
cond	i->1	
cont	r->2	
copy	r->1	
core	b->1	
corp	u->4	
corr	e->1	
cost	-->5	
coup	 ->1	
cour	s->1	
cove	r->1	
cque	s->3	
cqui	s->1	
cric	k->1	
ct. 	D->1	
ctne	s->1	
ctor	i->1	t->1	
cu m	e->1	
cu, 	e->1	
cy, 	s->1	
cyav	t->1	
cycl	i->1	
cyde	l->1	
cyfö	r->1	
cyke	l->3	
cykl	a->4	
cète	 ->1	
d "a	l->1	n->1	
d "e	n->1	
d (a	r->1	t->1	
d (e	f->1	
d (k	o->1	
d (r	å->1	
d - 	E->1	a->1	d->1	e->1	m->2	o->1	u->1	v->1	Ö->1	ä->1	
d 12	 ->2	
d 13	 ->2	
d 14	,->1	
d 16	4->1	
d 19	9->1	
d 2 	i->1	m->1	p->1	
d 20	 ->1	0->1	
d 24	 ->1	
d 27	 ->2	
d 28	 ->1	
d 30	 ->1	
d 36	7->1	
d 5 	0->1	
d 7 	p->1	
d 70	0->1	
d 80	 ->2	
d A.	 ->1	
d Ad	e->1	
d Am	o->1	s->1	
d BN	I->1	
d BS	E->1	
d Ba	l->1	r->2	
d By	r->3	
d Co	r->1	
d Da	l->1	v->1	
d E-	k->1	
d ED	D->1	
d EG	-->3	
d EU	-->3	
d Er	i->4	
d Eu	r->17	
d FP	Ö->1	
d Fr	a->4	
d GA	-->1	
d Ge	n->1	
d Gu	i->1	
d Ha	a->1	i->4	
d In	g->2	t->1	
d Is	l->1	r->1	
d Jö	r->1	
d Ko	u->3	
d Ku	l->2	
d Ky	o->1	
d LT	C->1	
d La	n->4	
d Le	a->1	
d Li	b->1	t->1	
d Ma	a->1	d->1	l->1	
d Me	d->1	
d Mi	d->1	
d OL	A->1	
d Os	l->1	
d Pa	d->1	t->1	
d Ry	s->1	
d Sa	v->1	
d Sv	e->1	
d Sy	d->1	r->4	
d Th	e->1	
d Ti	b->1	
d Tu	r->2	
d US	A->4	
d Va	n->1	
d Ve	r->1	
d Wi	d->1	
d a)	 ->1	
d ac	q->1	
d ad	m->2	
d al	l->41	t->1	
d an	a->1	d->18	g->1	k->1	l->6	n->19	s->13	t->7	v->6	
d ar	b->5	g->2	t->8	
d at	t->188	
d au	t->2	
d av	 ->136	.->1	f->1	s->20	t->1	
d ba	k->2	l->1	r->2	s->1	
d be	d->4	g->1	h->11	k->4	r->2	s->6	t->27	v->4	
d bi	b->2	d->3	l->4	n->1	
d bl	a->1	i->3	o->1	
d bo	m->2	
d br	a->3	i->3	o->1	y->1	ä->1	å->1	
d bu	d->1	
d by	g->2	
d bä	t->1	
d bå	d->2	
d bö	r->7	
d ca	.->1	
d ci	r->1	
d da	g->8	t->1	
d de	 ->87	f->1	l->5	m->16	n->109	r->4	s->29	t->90	
d di	r->7	s->1	
d do	k->2	m->3	
d dr	a->1	o->2	
d du	b->2	
d dy	l->1	s->1	
d dä	r->9	
d då	 ->4	
d ef	f->3	t->8	
d ek	o->2	
d el	e->1	l->12	
d en	 ->102	a->1	b->2	d->1	e->4	h->4	l->2	o->1	t->1	
d er	 ->9	.->2	a->3	b->1	t->1	
d et	t->42	
d eu	r->5	
d ev	e->1	
d ex	i->1	k->1	p->3	
d fa	l->1	m->1	r->3	s->1	t->2	
d fe	d->2	
d fi	c->1	n->6	
d fl	e->9	y->1	
d fo	n->1	r->6	
d fr	a->9	i->14	u->1	å->40	
d fu	l->3	n->8	
d fy	r->1	s->1	
d fä	l->1	
d få	 ->1	r->2	t->1	
d fö	l->2	r->173	t->1	
d ga	m->1	r->1	
d ge	m->6	n->7	r->2	
d gi	g->1	l->1	
d gj	o->2	
d gl	ä->2	
d go	d->6	t->1	
d gr	a->3	u->5	ä->1	ö->1	
d gä	l->60	
d gö	r->2	
d ha	 ->1	d->1	l->1	m->1	n->12	r->24	
d he	l->1	m->2	n->1	
d hi	t->1	
d hj	ä->26	
d ho	c->2	n->1	s->1	
d hu	n->1	r->4	
d hä	l->1	n->20	r->1	v->1	
d hå	l->1	
d hö	g->2	j->1	n->1	r->2	
d i 	E->4	F->1	L->1	M->3	S->1	a->2	b->4	d->16	e->9	f->7	h->4	j->1	k->4	l->2	m->4	o->1	p->3	r->3	s->8	t->3	u->4	v->3	ä->1	å->1	
d ib	l->1	
d id	é->3	
d if	r->1	
d im	p->2	
d in	 ->1	f->10	g->2	h->1	n->2	o->6	r->3	s->11	t->28	v->1	
d is	 ->2	
d iv	e->1	ä->1	
d ja	g->15	
d jo	r->3	
d ju	l->1	r->1	s->1	
d jä	m->3	
d ka	m->1	n->18	p->1	t->2	
d ki	n->1	
d kl	a->2	i->1	
d kn	a->1	
d ko	l->1	m->52	n->20	r->1	s->1	
d kr	a->6	i->4	ä->1	
d ku	l->3	n->1	s->1	
d kv	a->9	i->4	
d kä	n->1	r->2	
d kö	p->1	
d la	d->1	g->3	n->1	
d le	d->3	g->1	
d li	g->1	k->3	n->1	v->4	
d lu	n->1	
d lä	g->2	m->1	n->1	t->1	
d lö	p->1	s->3	
d ma	i->1	j->7	k->1	n->12	r->3	t->2	
d me	d->86	l->8	n->2	r->3	t->1	
d mi	g->5	k->2	l->9	n->24	t->2	
d mo	d->1	n->1	r->2	t->14	
d my	c->9	
d mä	n->1	
d må	l->2	n->4	s->13	
d mö	j->3	t->4	
d na	m->5	t->12	z->1	
d ne	g->3	
d ni	 ->4	,->1	
d no	t->1	
d nu	 ->2	m->1	v->1	
d ny	a->1	f->1	k->1	l->2	p->1	t->1	
d nä	m->2	r->7	s->1	
d nå	g->11	
d nö	d->5	j->2	t->1	
d oc	h->101	k->6	
d oe	r->1	
d of	f->2	
d oj	ä->1	
d ol	i->5	
d om	 ->67	.->1	b->1	f->2	r->5	s->5	
d op	t->1	
d or	d->6	m->1	o->1	
d os	s->13	ä->1	
d ot	i->1	
d pa	l->2	r->15	s->1	
d pe	n->3	r->5	
d pl	a->2	e->1	
d po	l->8	
d pr	e->1	i->7	o->8	ö->1	
d ps	y->1	
d pu	b->1	n->5	
d på	 ->48	f->1	l->1	
d ra	d->1	
d re	a->1	d->2	f->3	g->9	k->1	n->1	p->3	s->11	v->1	
d ri	k->3	
d ro	l->3	
d rä	d->1	t->15	
d rå	d->7	
d rö	s->1	t->1	
d s.	k->1	
d sa	k->4	m->15	
d se	 ->2	d->6	k->2	r->1	
d si	d->8	f->1	g->9	n->11	t->10	
d sj	u->1	ä->3	ö->1	
d sk	a->12	e->1	j->1	r->2	u->8	y->1	
d sl	a->1	u->2	ö->1	
d sm	ä->1	å->3	
d sn	e->2	
d so	c->7	m->138	
d sp	e->2	ä->3	
d st	a->8	i->1	o->22	r->9	y->1	ä->1	å->3	ö->9	
d su	b->3	
d sv	ä->1	å->1	
d sy	f->3	m->1	s->8	
d sä	g->8	k->8	l->1	r->3	
d så	 ->8	,->1	d->7	
d t.	e->1	o->1	
d ta	 ->2	c->1	g->10	l->3	n->43	r->1	
d te	k->1	m->1	r->1	x->1	
d ti	d->18	l->94	
d tj	ä->1	
d to	l->1	n->1	p->2	
d tr	a->5	e->6	o->2	
d tu	n->1	r->1	
d tv	i->1	å->7	
d ty	p->1	
d tä	c->1	n->2	t->1	
d un	d->10	g->1	i->2	
d up	p->15	
d ur	s->2	v->1	
d ut	a->11	b->4	f->1	g->2	n->1	s->8	v->11	
d va	c->1	d->7	l->3	n->1	r->16	
d ve	r->7	t->8	
d vi	 ->34	d->4	k->2	l->15	s->11	t->2	
d vo	n->1	
d vä	l->1	r->1	
d vå	r->22	
d yr	k->3	
d yt	t->5	
d ÖV	P->1	
d Ös	t->1	
d än	 ->5	d->6	n->2	
d är	 ->46	e->2	
d äv	e->2	
d år	 ->1	e->2	t->1	
d åt	 ->4	a->3	e->3	g->3	
d ök	a->1	n->1	
d öm	s->1	
d öp	p->2	
d ös	t->1	
d öv	e->31	r->2	
d! L	i->1	
d! N	i->1	
d) i	 ->1	
d), 	o->1	r->1	s->1	
d, "	a->1	
d, 5	6->1	
d, D	a->1	
d, E	C->1	
d, F	i->1	
d, I	t->2	
d, N	o->1	
d, S	p->2	
d, a	m->1	t->5	
d, b	l->1	o->1	ö->1	
d, d	e->5	v->1	ä->5	å->2	
d, e	f->3	k->1	n->4	t->1	
d, f	a->1	r->1	ö->5	
d, g	ö->1	
d, h	a->4	e->2	u->1	y->2	
d, i	 ->2	n->2	
d, k	a->1	o->1	r->1	
d, l	ä->1	
d, m	a->1	e->17	i->2	
d, n	ä->2	å->1	
d, o	c->25	m->4	
d, p	l->1	r->1	å->1	
d, r	e->1	ä->1	
d, s	a->1	k->2	o->10	p->2	t->2	ä->1	å->4	
d, t	i->1	o->1	r->2	y->1	
d, u	n->2	p->1	t->1	
d, v	a->3	i->6	
d, ä	r->2	v->1	
d- (	P->1	
d-af	f->1	
d-fö	r->1	
d-ko	s->1	
d. V	i->1	
d. Ö	s->1	
d. ö	s->1	
d."J	a->1	
d."M	e->1	
d.(S	a->1	
d., 	f->1	
d.- 	(->1	
d.. 	(->1	
d..(	D->1	
d.Al	l->1	
d.An	d->1	
d.At	t->2	
d.Be	d->1	
d.De	 ->4	n->8	s->1	t->36	
d.Di	r->2	
d.Dä	r->3	
d.Då	 ->1	
d.Ef	f->1	
d.Em	e->1	
d.En	 ->1	
d.Eu	r->3	
d.Fa	k->1	
d.Fr	å->2	
d.Fö	r->5	
d.Ge	n->1	
d.Ha	d->1	n->1	
d.He	r->13	
d.Hu	r->1	
d.I 	T->1	d->1	k->1	s->2	v->1	
d.In	f->1	i->1	n->1	
d.Ir	l->1	
d.Ja	g->23	
d.Ka	n->1	
d.Ko	m->5	n->1	
d.Lå	t->2	
d.Ma	n->1	
d.Me	n->8	
d.Mi	t->1	
d.Mo	t->1	
d.Mä	n->1	
d.Må	n->1	
d.Na	t->1	
d.Ni	 ->2	
d.Nu	 ->2	
d.Nä	r->2	
d.Om	 ->3	r->14	
d.Or	d->1	
d.Pa	r->1	
d.På	 ->1	
d.Re	g->3	
d.Sa	v->1	
d.So	m->2	
d.Su	b->1	
d.Så	 ->1	
d.Ta	c->1	
d.Ti	l->1	
d.Tr	o->1	
d.Un	d->1	
d.Up	p->1	
d.Ut	a->1	g->1	
d.Va	d->1	r->1	
d.Ve	t->1	
d.Vi	 ->11	l->1	s->1	
d.Än	d->1	
d.Äv	e->1	
d.Å 	a->2	
d.År	 ->1	
d: "	D->1	O->1	
d: d	e->1	
d: e	n->1	
d; d	e->3	
d; i	n->2	
d? H	a->1	
d?- 	(->2	
d?. 	(->1	
d?Dä	r->1	
d?Fö	r->1	
d?He	r->1	
d?Ja	g->1	
d?Vi	 ->1	
d?Är	 ->1	
da -	 ->1	
da 1	2->1	
da 2	0->1	
da 6	0->1	
da C	o->5	
da E	U->2	r->1	u->3	
da F	e->1	
da G	o->1	
da a	g->2	k->1	l->6	n->5	r->6	t->26	v->13	
da b	a->2	e->7	i->2	o->2	å->1	
da c	h->2	i->1	
da d	e->50	i->2	j->2	o->5	r->1	
da e	f->2	k->2	l->5	n->19	r->2	t->7	u->3	x->1	
da f	a->3	i->3	o->4	r->7	ö->43	
da g	a->1	e->2	i->1	r->3	ä->1	ö->1	
da h	a->5	i->1	u->2	y->1	ä->2	ö->1	
da i	 ->19	d->1	g->2	n->17	
da j	a->2	o->2	
da k	a->2	o->14	r->3	u->1	v->1	ä->1	
da l	a->4	e->1	i->1	o->2	u->1	ä->4	ö->1	
da m	a->3	e->22	i->6	o->4	y->2	ä->2	å->3	ö->3	
da n	a->1	e->1	i->2	y->2	ä->1	å->3	ö->2	
da o	c->14	d->1	l->1	m->6	r->3	s->6	
da p	a->8	e->5	h->1	l->3	o->5	r->7	u->1	å->5	
da r	a->1	e->17	i->2	y->1	ä->3	å->1	ö->3	
da s	a->2	c->1	e->5	i->20	k->8	m->1	o->15	t->10	u->2	y->1	ä->8	
da t	a->1	e->1	i->41	o->1	r->6	u->1	å->1	
da u	n->4	p->3	r->1	t->8	
da v	a->2	e->2	i->10	ä->2	å->2	
da ä	n->3	r->4	
da å	t->8	
da ö	a->1	r->1	v->2	
da!D	e->1	
da" 	b->1	
da, 	J->1	b->1	d->1	e->2	f->5	h->2	i->2	k->1	m->3	n->1	o->3	p->1	r->2	s->8	t->1	v->4	ä->1	
da. 	E->1	
da.B	e->1	
da.D	e->5	å->1	
da.E	t->1	
da.F	r->2	ö->1	
da.H	a->1	e->4	
da.I	 ->1	b->1	
da.J	a->3	
da.K	ä->1	
da.M	e->2	i->1	
da.N	i->1	ä->1	
da.O	c->2	
da.R	u->1	
da.V	a->1	i->4	
da.Ä	r->1	v->1	
da?D	e->2	
da?F	r->1	
da?I	n->1	
dabo	c->2	
dac 	b->2	o->1	
dac"	,->1	
dac-	s->1	
dad 	a->1	b->1	i->1	p->3	r->1	s->1	
dad.	S->1	
dade	 ->23	,->1	.->1	s->6	
dafo	n->1	
dafr	i->2	
dag 	-->3	I->1	a->11	b->1	d->4	e->5	f->15	g->3	h->21	i->15	j->1	k->6	l->4	m->8	n->2	o->9	p->3	r->4	s->10	t->12	u->4	v->6	Ö->1	ä->16	
dag,	 ->32	
dag.	 ->1	(->1	A->2	D->9	E->1	F->2	G->1	H->3	I->2	J->7	K->1	L->1	O->1	V->1	
dag:	 ->1	D->1	
daga	r->17	s->1	
dage	n->36	
dagl	i->8	
dago	g->1	r->52	
dags	 ->17	,->2	.->1	b->1	l->2	t->2	
dahå	l->43	
dair	e->1	
daki	s->3	
dakt	i->1	ö->2	
dal!	H->1	
dal,	 ->1	
dala	g->4	n->1	
dale	r->5	
daly	d->2	
dalö	s->1	
dam 	-->1	1->1	i->1	o->1	p->1	s->2	t->1	v->1	ä->1	
dam,	 ->3	
dam.	N->1	
dama	f->1	
dame	n->1	r->45	
damf	ö->27	
damm	 ->1	a->3	
damo	t->74	
damr	e->1	
damå	l->13	
damö	t->84	
dan 	-->1	1->15	4->1	A->1	E->1	F->1	P->1	S->1	a->24	b->16	d->30	e->20	f->32	g->10	h->50	i->26	j->4	k->15	l->7	m->14	n->11	o->13	p->11	r->8	s->25	t->21	u->10	v->19	ä->12	å->1	ö->3	
dan,	 ->17	
dan.	A->1	D->8	H->1	I->1	J->5	S->2	
dan?	 ->1	H->1	S->1	
dana	 ->52	n->1	
danb	e->2	
dand	e->105	r->1	
danf	l->1	
dang	e->1	
danh	å->1	
dani	e->1	
danm	a->1	
dano	r->1	
danr	ö->6	
dans	 ->1	k->25	v->7	
dant	 ->53	,->1	a->39	
dape	s->1	
dar 	a->9	b->1	d->6	e->2	g->1	h->1	i->3	j->1	m->5	n->1	o->1	r->3	s->4	
dar,	 ->2	
dar.	D->1	J->1	
darb	e->2	
dard	 ->6	,->2	.->1	;->1	e->5	i->9	
dare	 ->85	,->8	.->9	?->2	b->3	n->5	s->4	u->4	
darf	ö->1	
dari	s->2	t->29	
darn	a->23	
dars	 ->1	k->2	y->1	
das 	a->2	d->1	f->2	g->1	i->7	m->2	n->1	o->1	p->10	r->1	s->1	t->5	u->3	ö->1	
das,	 ->5	
das.	A->1	B->1	D->3	H->2	I->3	M->1	T->1	V->1	Å->1	
das?	H->1	
dast	 ->84	.->1	e->1	
dat 	a->6	b->1	d->1	f->4	h->1	k->1	m->1	n->1	p->4	s->3	u->1	
dat,	 ->4	
dat.	F->1	T->1	
data	 ->1	,->1	b->1	s->1	
date	n->1	r->6	t->4	
dati	o->33	
datl	a->1	i->1	ä->10	
dato	 ->1	r->2	
datp	e->9	
dats	 ->4	,->2	.->2	
datu	m->13	
dbar	 ->1	a->3	t->5	
dbed	d->1	
dbel	ä->1	
dbes	l->16	t->1	
dbet	ä->1	
dbor	g->170	
dbro	t->1	
dbru	k->56	
dbrä	n->1	
dbul	t->1	
dbäv	n->10	
dd a	t->17	v->5	
dd b	a->1	ö->1	
dd e	l->1	
dd f	ö->18	
dd h	ä->1	
dd i	 ->1	n->1	
dd m	e->1	o->3	å->1	
dd o	c->4	
dd s	a->2	o->1	t->1	
dd t	i->3	
dd u	t->2	
dd v	i->2	
dd ä	n->2	
dd ö	v->1	
dd),	 ->1	
dd, 	d->1	e->1	h->1	v->1	
dd.D	e->2	
dd.J	a->2	
dd.M	e->1	
dd.N	a->1	
dd.R	e->1	
dd.V	i->1	
dda 	6->1	a->16	c->1	d->6	e->1	f->2	g->3	i->2	k->3	l->2	m->6	o->1	p->1	r->4	s->5	t->1	u->2	v->1	
dda.	 ->1	M->1	
ddad	 ->1	e->5	
ddag	 ->4	,->2	.->1	e->2	s->4	
ddan	d->1	
ddar	 ->1	e->1	s->1	
ddas	.->2	
ddat	s->1	
dde 	"->1	4->1	A->2	V->1	a->2	d->4	e->1	f->5	i->6	j->1	m->1	p->4	t->7	v->1	
dde,	 ->1	
ddel	 ->1	a->59	e->2	h->1	
dden	 ->2	,->1	
dder	 ->1	
ddes	 ->10	.->1	
ddet	 ->16	,->2	
ddhi	s->1	
ddig	h->1	t->1	
ddin	g->2	
ddit	i->1	
ddni	n->4	
dds 	e->1	
ddsm	e->4	
ddsn	i->6	
ddso	m->1	r->1	
ddsp	r->1	
ddss	t->1	ä->1	
ddst	u->1	
de "	a->2	d->1	f->1	k->2	l->2	s->1	
de (	A->29	m->1	
de -	 ->20	
de 1	1->1	2->1	4->3	5->1	8->1	9->3	
de 2	0->1	5->4	6->1	
de 4	0->1	1->1	
de 8	 ->1	
de 9	 ->1	
de A	h->1	l->2	m->2	
de B	 ->1	u->1	
de C	e->2	
de D	a->1	u->1	
de E	U->1	u->7	
de F	r->1	
de G	a->3	r->2	
de H	a->1	e->1	o->1	
de I	m->1	r->1	
de J	a->1	
de K	a->2	i->1	o->3	
de L	a->1	o->1	
de M	a->4	e->1	
de N	a->2	
de O	L->1	i->1	
de P	a->6	r->14	
de R	a->1	o->2	
de S	a->1	c->2	e->1	v->1	w->1	
de T	r->1	u->1	
de V	a->1	e->1	
de W	e->1	
de a	b->1	d->6	f->1	g->2	i->1	k->5	l->26	m->4	n->60	p->2	r->20	s->2	t->69	v->177	
de b	a->11	e->83	i->18	l->8	o->2	r->16	u->2	y->6	ä->5	å->9	ö->3	
de c	e->3	h->1	
de d	a->10	e->107	i->16	j->1	o->5	r->13	ä->12	å->4	ö->1	
de e	f->11	g->5	j->1	k->22	l->9	m->2	n->52	p->1	r->3	t->16	u->55	v->1	x->21	
de f	a->36	e->9	i->22	j->3	l->29	o->14	r->99	u->6	y->8	ä->1	å->17	ö->179	
de g	a->12	e->23	i->1	j->3	l->1	o->10	r->32	ä->2	å->5	ö->5	
de h	a->67	e->13	i->8	j->1	o->7	u->2	y->2	ä->18	å->5	ö->7	
de i	 ->117	c->8	d->3	f->1	g->1	n->136	s->3	t->5	
de j	a->17	o->4	u->5	ä->1	
de k	a->42	e->1	i->5	l->4	n->2	o->113	r->18	u->33	v->8	ä->3	
de l	a->13	e->12	i->13	o->10	y->2	ä->15	å->4	ö->1	
de m	a->30	e->90	i->33	o->8	u->4	y->18	ä->38	å->46	ö->5	
de n	a->49	e->3	i->6	o->9	u->10	y->28	ä->22	å->7	ö->3	
de o	b->3	c->121	e->1	f->11	l->49	m->105	n->2	p->2	r->23	s->5	t->1	v->3	
de p	a->26	e->28	l->5	o->36	r->66	u->8	å->59	
de r	a->8	e->102	i->21	o->7	u->3	ä->41	å->8	ö->2	
de s	a->24	e->45	i->26	j->4	k->48	l->4	m->21	n->2	o->102	p->4	t->92	u->3	v->12	y->26	ä->27	å->7	
de t	.->1	a->23	e->7	i->87	j->8	o->3	r->22	u->3	v->23	y->4	ä->1	
de u	l->1	n->17	p->23	r->5	t->56	
de v	a->40	e->31	i->65	o->3	r->1	ä->19	å->4	
de y	r->3	t->11	
de Ö	s->1	
de ä	g->1	l->1	m->1	n->18	r->53	v->2	
de å	 ->1	r->19	s->4	t->54	
de ö	a->1	k->1	m->1	n->4	p->3	s->3	v->33	
de! 	J->5	N->1	
de!A	l->1	
de!J	a->1	
de!N	i->1	
de",	 ->1	
de(A	5->1	
de, 	,->1	D->1	E->1	F->1	G->1	L->1	a->9	b->6	d->10	e->6	f->9	h->10	i->14	j->2	k->7	l->1	m->13	n->8	o->25	p->4	s->16	t->7	u->3	v->12	ä->3	ö->1	
de- 	o->1	
de-F	r->2	
de-L	o->1	
de-l	ä->1	
de. 	D->2	M->1	O->1	V->2	
de.-	 ->1	
de..	 ->1	
de.A	t->1	v->3	
de.D	e->39	ä->4	
de.E	f->2	m->1	n->5	u->1	
de.F	P->1	r->2	ö->7	
de.G	e->1	r->1	
de.H	a->2	e->7	o->1	u->5	
de.I	 ->3	d->1	n->2	
de.J	a->35	
de.K	a->2	o->2	
de.L	i->1	y->1	å->2	
de.M	a->4	e->10	i->3	å->1	
de.N	i->1	u->1	ä->2	
de.O	c->3	m->3	
de.P	a->1	l->1	o->1	r->1	
de.R	e->1	
de.S	a->1	c->1	e->1	l->2	o->4	t->1	å->2	
de.T	V->1	a->4	i->1	o->1	r->2	v->1	
de.U	n->2	
de.V	a->3	i->10	
de.Å	t->1	
de: 	"->2	A->3	D->2	F->3	G->3	H->1	I->1	J->2	K->3	M->1	N->2	P->1	S->2	T->1	U->1	V->3	b->1	f->1	h->1	i->1	k->1	t->1	Å->2	
de; 	d->2	h->1	m->1	p->1	
de?D	e->1	
de?F	ö->1	
de?H	e->3	
de?J	a->1	
de?V	i->1	
deHe	r->1	
dePr	o->1	
dead	l->1	
deal	,->1	a->1	e->2	i->1	
deau	x->1	
deba	t->170	
debe	s->1	
debu	d->9	
debä	n->1	
dece	m->19	n->22	
dede	l->2	
deel	l->2	
deer	s->2	
defi	n->36	
defo	n->1	
defr	i->1	
defu	l->7	
defö	r->13	
dege	m->3	n->1	
degr	a->1	
dehö	j->1	
deir	a->2	
deko	d->8	l->1	
dekr	i->1	
dekv	a->5	
del 	(->2	-->1	K->1	a->84	b->3	d->1	f->22	h->3	i->13	k->4	l->1	m->8	n->1	o->15	p->8	s->16	t->5	u->3	v->1	ä->8	ö->1	
del,	 ->23	
del.	B->1	D->5	E->2	J->2	M->3	N->1	S->1	V->5	
del?	J->1	
dela	 ->21	d->11	g->1	k->8	n->44	r->73	s->10	t->17	y->2	
delb	a->19	
dele	g->20	n->36	s->23	
delf	r->1	
delg	i->1	
delh	a->3	o->1	
dell	 ->3	"->2	.->1	e->6	å->4	ö->1	
deln	 ->2	i->41	
delp	u->2	
delr	a->1	
dels	 ->15	-->1	d->1	e->134	f->4	h->2	i->2	k->5	l->6	m->11	n->1	o->5	p->6	s->46	t->46	v->1	
delt	a->56	i->2	o->2	
delu	t->2	
delv	i->11	
delö	s->1	
dem 	2->1	a->6	d->7	e->6	f->8	g->2	h->3	i->10	j->1	k->1	l->1	m->5	n->1	o->10	p->7	r->1	s->61	t->5	u->4	v->2	ä->1	
dem,	 ->11	
dem.	(->1	A->1	B->2	D->6	E->1	F->2	H->1	J->4	K->1	M->3	N->2	O->1	R->1	V->6	
dem:	 ->2	
dem?	D->1	
dema	g->4	r->1	s->1	
deme	n->5	
demi	,->1	n->1	s->1	
demo	g->3	k->136	n->14	
den 	"->3	(->1	,->1	-->11	1->33	2->18	3->7	4->2	5->1	6->1	7->1	9->2	B->2	E->4	G->2	J->1	K->5	L->1	P->3	R->1	T->1	X->1	a->147	b->88	c->3	d->63	e->174	f->191	g->100	h->118	i->180	j->4	k->84	l->24	m->96	n->77	o->131	p->106	r->64	s->278	t->90	u->39	v->55	z->1	ä->52	å->13	ö->31	
den"	 ->1	
den)	 ->1	(->2	,->1	.->1	
den,	 ->121	
den.	 ->3	.->3	A->6	D->39	E->7	F->12	H->11	I->9	J->18	K->7	L->2	M->10	N->3	O->4	P->4	R->1	S->8	T->3	U->2	V->16	Ä->1	
den:	 ->6	F->1	
den;	 ->4	
den?	D->3	N->1	V->2	
denN	ä->1	
dena	 ->53	,->13	.->13	;->1	?->1	s->1	u->1	
denb	u->2	
deni	e->2	
denn	a->522	e->5	
dens	 ->58	,->2	a->4	e->7	i->2	
dent	 ->5	,->1	e->5	i->20	l->25	s->1	
deol	o->5	
depa	r->9	
der 	-->4	1->8	2->2	4->1	E->6	F->2	I->2	L->7	N->2	U->2	a->40	b->23	d->165	e->53	f->97	g->14	h->29	i->69	j->5	k->26	l->9	m->70	n->19	o->65	p->34	r->19	s->147	t->48	u->21	v->37	ä->11	å->11	ö->1	
der"	 ->1	
der)	 ->2	F->2	J->1	K->1	T->1	
der,	 ->69	
der-	p->1	
der.	 ->4	.->1	A->4	B->2	C->1	D->26	E->3	F->5	H->1	I->7	J->12	K->3	M->3	N->2	O->1	R->1	S->2	T->2	U->4	V->5	Ä->3	
der:	 ->1	
der;	 ->1	
der?	.->1	H->1	Ä->1	
dera	 ->30	,->1	.->1	d->7	l->10	n->1	r->27	s->93	t->8	
derb	a->1	l->2	ö->11	
derd	e->4	o->2	
dere	g->3	
derg	r->4	ä->1	
derh	u->2	å->3	
deri	,->1	e->2	n->59	
derk	a->4	u->1	
derl	a->7	e->2	i->10	ä->37	å->3	
derm	a->3	e->1	i->1	å->1	
dern	 ->7	,->1	a->260	e->1	i->24	t->1	
dero	r->4	
derr	e->2	ä->1	
ders	 ->26	a->1	k->6	m->1	p->2	t->39	å->1	ö->48	
dert	a->1	e->17	i->1	
deru	t->3	
derv	i->1	ä->1	
derä	t->3	
derö	s->1	
des 	-->2	1->3	2->1	A->1	S->1	V->1	a->30	b->6	d->12	e->10	f->19	g->2	h->8	i->33	j->1	k->7	l->1	m->8	n->4	o->12	p->5	r->2	s->9	t->13	u->9	v->6	ä->2	
des,	 ->8	
des.	)->1	D->2	I->1	J->1	M->2	R->1	U->1	
desa	m->2	
desb	e->1	
desd	i->2	
desg	e->1	
desk	a->113	i->1	y->1	
desp	e->7	
dess	 ->101	a->344	k->1	t->1	u->36	v->4	
dest	a->1	o->2	r->1	å->1	
desv	i->2	
det 	"->4	(->7	-->8	2->2	A->1	B->2	C->1	E->4	G->1	I->1	K->1	M->3	P->3	S->2	T->1	a->404	b->115	c->5	d->63	e->127	f->423	g->243	h->162	i->211	j->16	k->111	l->39	m->139	n->90	o->132	p->99	r->52	s->384	t->93	u->57	v->175	y->6	ä->339	å->13	ö->29	
det!	.->2	
det)	 ->1	N->1	
det,	 ->119	
det.	 ->6	(->2	-->1	.->2	A->6	B->1	D->26	E->10	F->2	H->12	I->7	J->20	K->1	L->1	M->13	N->3	O->2	P->5	S->5	T->2	U->2	V->21	Ä->1	Å->2	Ö->1	
det:	 ->3	
det;	 ->1	
det?	.->2	D->2	H->1	I->1	J->1	N->1	V->1	
deta	k->1	l->34	
dets	 ->115	,->1	a->5	
dett	a->829	
deur	o->2	
deut	r->1	
deva	l->6	
devi	s->2	
dez,	 ->1	
dez-	k->2	
dfil	m->1	
dfin	a->2	
dfrå	g->10	
dful	l->1	
dfäl	l->4	
dföd	d->1	
dför	 ->10	,->2	a->227	d->2	e->2	s->1	t->2	u->2	
dga 	E->2	d->4	f->5	g->1	k->2	m->3	o->3	p->1	s->2	u->2	ä->2	ö->1	
dga,	 ->1	
dga?	D->1	
dgad	 ->4	e->2	
dgan	 ->9	.->1	
dgar	 ->4	.->1	
dgas	 ->5	,->2	.->6	
dgat	 ->3	
dge 	F->1	a->3	
dger	 ->10	
dges	 ->5	
dget	 ->9	,->4	.->6	a->3	b->1	e->16	f->11	k->17	m->1	p->14	s->4	t->1	u->10	å->10	ö->1	
dgiv	a->23	i->2	n->3	
dgni	n->71	
dgor	 ->1	
dgrä	n->1	
dgrö	n->1	
dgän	g->2	
dgån	g->2	
dgår	d->2	
dgåt	t->1	
dgör	 ->1	l->2	
dhet	 ->8	.->1	e->3	s->13	
dhis	t->1	
dhjä	l->1	
dhål	l->4	
dhöl	l->1	
di -	 ->1	
di a	t->2	v->1	
di b	e->1	
di h	a->2	
di i	n->1	
di l	o->1	ä->1	
di o	c->5	
di r	e->1	
di s	o->2	
di t	a->2	
di, 	v->1	
di.D	e->1	
di.S	o->1	
di.V	i->1	
di: 	f->1	
di; 	m->1	
dia 	-->1	a->1	h->1	s->2	
dial	 ->1	o->31	
diar	i->21	
dias	 ->1	
diat	ä->1	
dica	p->1	
dice	r->1	
dici	n->1	
dida	t->14	
die 	R->1	a->1	o->1	
die,	 ->1	
dieb	e->1	
diek	t->1	
dien	 ->4	s->3	
diep	r->1	
dier	 ->7	,->2	.->3	n->2	
diet	 ->3	.->1	
diff	e->5	
difi	e->5	
dig 	a->1	b->1	d->4	e->3	f->8	g->1	h->1	i->3	j->1	l->2	m->3	n->1	o->6	p->1	r->4	s->2	t->4	
dig,	 ->2	
dig.	D->1	E->1	M->1	P->1	U->1	
diga	 ->59	,->3	.->4	n->4	r->86	t->1	
dige	n->1	s->1	
digh	e->250	
dign	a->1	
digr	a->2	
digs	t->1	
digt	 ->212	,->10	.->5	?->1	v->7	
dika	l->16	p->4	t->9	
dike	n->1	
dikt	a->3	e->2	i->5	
dile	m->3	
dime	n->13	
dina	v->1	
dinb	u->1	
dinf	l->1	
ding	 ->5	,->3	s->1	t->2	
dins	a->1	k->1	t->1	
dinä	r->1	
diol	o->2	
diox	i->7	
dipl	o->11	
dire	k->248	
diri	g->1	
dirl	ä->2	
dis 	B->1	l->1	p->2	s->1	u->1	v->2	
disc	i->14	
dise	r->9	
disk	 ->9	a->32	r->21	t->10	u->141	
disp	e->1	o->3	
dist	a->1	i->1	r->2	
dit 	F->1	a->1	d->2	f->2	h->1	l->1	r->1	s->3	t->1	
dita	l->1	
dite	r->2	
dith	ö->1	
diti	o->22	
dits	 ->1	
dium	 ->3	.->1	
dive	r->4	
divi	d->14	
diz 	e->1	f->2	
diz,	 ->1	
diz-	k->1	
diär	,->1	
dja 	-->1	D->1	H->1	a->2	d->28	e->4	f->4	i->1	k->4	l->1	m->2	o->5	p->1	r->1	s->5	t->2	u->1	v->1	Ö->1	å->3	
dja.	H->1	J->1	
djan	 ->3	d->3	
djar	 ->6	
djas	 ->6	,->2	
dje 	-->1	a->2	b->2	d->2	f->3	g->3	k->1	l->24	m->4	n->1	o->2	p->6	r->2	s->1	v->4	ä->1	å->1	ö->3	
dje,	 ->4	
dje:	 ->1	
djed	e->6	
djek	t->2	
djel	a->6	
djer	 ->1	
djor	n->1	
djun	g->2	
djup	 ->1	a->13	e->5	g->7	n->5	s->1	t->7	
djur	 ->2	,->2	-->2	.->2	a->1	e->2	f->4	l->2	
djär	v->7	
djäv	u->2	
dkar	e->1	
dkom	m->24	
dkor	e->1	
dkur	s->1	
dkus	t->2	
dkvi	s->1	
dkän	d->25	n->46	s->5	t->18	
dla 	d->7	f->1	g->1	i->2	m->1	o->7	s->1	u->1	v->2	
dla.	D->1	V->1	
dlad	 ->1	e->10	
dlag	 ->1	d->1	
dlan	d->1	
dlar	 ->116	e->4	n->2	
dlas	 ->12	,->1	.->1	
dlat	 ->6	s->1	
dlem	 ->5	,->1	m->14	s->323	
dlen	 ->10	,->2	
dlet	 ->1	
dlid	a->2	
dlig	 ->30	,->1	:->1	a->51	e->16	g->4	h->5	t->91	
dlin	e->1	g->190	j->2	
dlis	t->1	
dläg	g->79	
dlös	a->1	
dmak	t->1	
dmed	e->3	l->1	
dmin	i->25	
dmiu	m->3	
dmon	t->3	
dmot	t->1	
dmän	 ->1	
dmål	e->1	s->1	
dmån	 ->1	
dna 	d->1	e->1	f->1	g->1	k->1	l->1	m->1	r->1	s->2	t->1	u->1	v->1	
dnac	k->2	
dnad	 ->6	e->4	
dnan	d->2	
dnap	p->1	
dnar	 ->1	e->3	n->1	
dnas	 ->2	
dnat	 ->2	s->1	
dnin	g->407	
dniv	å->1	
do R	o->1	
do a	n->1	t->3	
do, 	a->1	
do.D	e->1	
do.F	ö->1	
do.H	e->1	
do.O	m->1	
dock	 ->59	,->2	
doef	f->1	
dofi	l->1	
dog 	i->1	
dog.	D->1	S->1	
dogj	o->1	
dogm	 ->1	a->1	
dogö	r->9	
doku	m->45	
dolf	 ->2	
doll	a->9	
dom 	a->4	b->1	d->1	f->1	g->1	i->1	n->1	o->5	p->1	r->1	ä->1	
dom,	 ->5	
dom.	D->1	
dom/	r->1	
doma	r->28	
dome	n->10	
domi	n->8	
doml	i->3	
domr	å->14	
doms	 ->1	-->3	b->1	f->4	g->1	h->1	l->3	r->1	t->83	
don 	(->2	-->1	b->2	e->1	f->1	i->3	k->1	m->1	o->3	p->3	s->13	u->1	ä->1	
don,	 ->10	
don.	D->3	J->3	L->1	M->1	O->1	V->1	
don?	V->1	
donN	ä->1	
done	n->6	t->1	
dons	i->1	p->1	t->3	ä->1	å->1	
dont	 ->1	
dor 	d->1	f->2	h->1	o->2	p->2	s->6	u->1	v->1	
dor,	 ->4	
dor.	D->1	H->1	K->1	M->1	
dord	e->1	
dore	r->2	
dorn	a->11	
dors	a->1	
dosa	m->1	
dose	d->1	
dosk	o->3	
dost	a->1	e->1	
dou 	f->1	
dovi	s->4	
dox,	 ->1	
doxa	l->5	
doäm	n->1	
dpel	a->1	
dpol	i->1	
dpri	n->1	
dpun	k->119	
dra 	-->1	E->3	L->2	R->1	a->24	b->17	d->24	e->14	f->33	g->14	h->12	i->23	k->13	l->17	m->30	n->10	o->28	p->25	r->18	s->52	t->43	u->4	v->13	y->2	ä->7	å->3	ö->1	
dra,	 ->23	
dra.	D->2	J->1	N->2	U->1	V->1	
dra:	 ->4	
dra;	 ->2	
drab	b->50	e->5	
drad	 ->1	e->24	
drag	 ->61	,->2	.->6	:->1	a->114	e->151	i->12	n->49	s->21	
drah	a->1	
drak	a->1	
dram	 ->1	a->7	
dran	 ->7	,->1	.->1	d->5	
drar	 ->60	,->1	e->6	n->3	
dras	 ->23	,->2	.->5	t->3	
drat	 ->9	a->5	s->10	u->3	
dre 	a->2	b->3	d->1	e->3	f->8	g->1	h->1	i->1	k->4	l->3	m->1	o->4	p->4	r->1	s->4	t->2	u->5	v->1	ä->10	
dre,	 ->2	
dre.	D->2	
dre?	V->1	
drek	o->1	
dren	 ->3	
dres	a->2	
dret	 ->1	
drev	s->1	
dria	t->2	
dric	k->3	
drid	 ->1	,->1	.->1	
drif	t->8	
drig	 ->32	
drik	t->3	
drin	g->315	
driv	a->25	e->18	k->3	n->1	s->7	
drog	 ->5	b->1	e->1	k->1	s->2	
drol	l->2	
drom	e->1	
dron	 ->1	
drop	p->1	
drot	t->4	
druc	k->2	
drun	k->3	
drus	t->1	
dryf	t->1	
dryg	t->3	
dräg	e->36	l->1	
drän	g->1	k->2	
dråp	s->1	
dröj	a->2	d->1	e->3	s->2	
dröm	m->1	
ds a	l->1	n->1	t->1	v->6	
ds b	e->4	l->2	å->1	
ds d	e->2	ä->1	
ds e	f->1	m->1	n->1	
ds f	e->1	ö->4	
ds g	e->1	r->1	
ds i	 ->5	n->4	
ds j	u->1	
ds l	a->1	i->1	
ds m	e->5	y->1	
ds n	y->1	
ds o	b->1	c->1	m->1	
ds p	a->1	å->25	
ds r	e->3	å->1	
ds s	a->1	k->4	o->2	
ds t	a->1	i->1	r->1	
ds u	n->1	t->1	
ds v	e->1	i->1	
ds ä	n->1	
ds å	r->1	t->3	
ds ö	k->1	v->1	
ds, 	m->1	o->1	s->1	t->1	
ds- 	o->2	
ds-i	n->2	
ds-n	y->1	
ds-s	i->1	
ds. 	D->1	
ds.B	e->1	
ds.D	e->1	
ds.J	a->1	
ds.U	n->1	
ds/i	n->1	
ds; 	b->1	
dsNä	s->1	
dsak	 ->6	l->10	t->1	
dsam	 ->2	m->1	t->4	
dsan	d->3	m->1	s->1	
dsar	b->5	
dsat	s->1	
dsav	g->3	t->3	
dsbe	d->1	f->6	h->1	s->3	v->1	
dsbu	s->1	
dsby	g->43	
dsce	n->1	
dsde	l->13	
dsdi	r->3	
dsdo	m->1	
dsdu	g->1	
dsdö	m->1	
dsef	f->4	
dsek	o->15	
dsen	 ->1	,->1	
dset	 ->1	s->1	
dsfa	l->1	
dsfr	i->14	å->1	
dsfö	r->8	
dsgr	ä->1	
dsha	n->6	
dsin	f->2	r->2	s->2	t->2	
dsit	u->1	
dsju	k->1	
dsk 	a->1	k->3	t->1	
dsk-	b->1	
dska	 ->19	,->2	d->2	l->1	n->19	p->13	r->1	s->8	
dsko	g->1	m->1	n->4	
dskr	a->1	i->6	ä->1	
dskt	 ->1	
dskä	r->3	
dsla	 ->4	,->1	.->1	g->3	n->3	
dsli	b->1	g->1	s->1	
dslä	n->2	
dslå	n->1	
dslö	s->2	
dsma	n->10	r->1	
dsme	d->11	
dsmi	n->1	
dsmy	n->2	
dsmä	n->3	s->2	
dsmå	l->1	
dsmö	j->1	t->1	
dsni	v->8	
dsom	r->7	s->1	
dsor	d->20	g->2	i->1	
dspa	k->2	r->1	t->2	
dspe	n->6	r->4	
dspl	a->11	
dspo	l->3	
dspr	i->2	o->32	
dspu	n->1	
dsra	m->5	
dsre	g->3	p->4	
dsry	m->2	
dsrä	t->1	
dsrö	r->1	
dssa	m->4	
dssk	i->1	ä->1	
dsst	a->5	ä->24	ö->1	
dssy	s->2	
dssä	l->1	
dsta	d->2	g->2	
dste	n->1	
dsti	l->1	
dstj	ä->2	
dsto	p->1	w->3	
dstr	ä->1	
dstu	l->1	r->1	
dstä	d->2	m->1	n->2	
dsup	p->2	
dsut	t->1	v->2	
dsve	r->1	
dsvi	l->2	n->1	
dsvä	g->1	
dsyf	t->1	
dsys	t->4	
dsän	d->1	
dsål	d->2	
dsåt	g->1	
dsöd	a->1	
dt f	r->1	
dt h	a->1	
dt o	c->3	
dt s	a->1	
dt t	a->1	
dt u	t->1	
dt, 	O->1	f->2	i->1	
dta 	a->1	d->4	e->6	f->10	g->2	j->1	k->1	l->1	m->3	n->2	o->1	p->2	s->1	u->1	ä->3	å->5	
dta.	D->1	
dtab	e->6	
dtag	b->15	i->8	n->1	
dtal	a->1	
dtar	 ->11	
dtas	 ->14	,->2	.->5	
dter	 ->5	,->1	H->1	b->2	s->5	
dtes	,->1	
dtid	.->1	
dtog	 ->2	s->2	
dtyc	k->6	
dtys	k->1	
du b	a->1	e->1	
du c	o->1	
du m	i->1	
du ä	r->2	
dual	i->1	
dubb	e->6	l->11	
duce	n->22	r->13	
duel	l->7	
duer	,->1	
duga	,->1	
dugl	i->6	
duka	r->1	
dukt	 ->5	,->1	e->14	i->32	s->2	
dumh	e->3	
dump	a->1	n->3	
dumt	 ->1	
duna	n->1	
dunk	l->1	
dupp	b->1	g->1	r->2	
durr	e->1	
duss	i->1	
dust	r->114	
duts	l->1	
duty	p->1	
dvag	n->1	
dval	 ->20	a->3	e->1	
dvat	t->1	
dver	k->19	
dvet	a->4	e->21	n->17	
dvik	a->31	e->3	i->1	l->4	
dvin	n->2	
dvis	 ->3	
dvok	a->5	
dvri	d->12	
dvrä	n->1	
dvs.	 ->45	
dvun	n->1	
dvän	d->126	
dvär	d->1	
dväs	t->2	
dwil	l->1	
dyka	 ->2	
dyke	r->5	
dyli	k->3	
dyna	m->5	
dyr 	h->1	
dyra	 ->2	r->2	
dyrk	a->1	
dyrt	 ->1	.->1	
dyst	r->1	
dzio	-->4	
dzji	k->5	
däck	 ->1	
dämp	a->2	
där 	-->1	1->1	2->1	5->1	8->1	E->4	F->1	L->1	a->9	b->7	d->43	e->8	f->6	g->3	h->9	i->5	j->3	k->8	l->1	m->29	n->5	o->3	p->4	r->2	s->16	t->4	u->5	v->27	Ö->1	ä->4	å->1	
där!	D->1	
där,	 ->10	
där.	 ->1	D->2	F->1	I->1	J->3	S->3	V->3	
där?	J->1	
dära	v->2	
däre	f->7	m->13	
därf	ö->184	
därh	ä->1	
däri	 ->1	b->6	f->2	g->15	
därm	e->40	
därp	å->2	
därr	ä->1	
därt	i->1	
därv	a->2	b->1	i->4	l->1	
då 2	4->1	
då A	s->1	
då D	a->1	
då E	G->1	r->1	u->1	
då a	k->1	l->2	n->3	r->2	t->11	
då b	a->2	e->6	l->3	o->1	ö->4	
då d	e->16	å->1	
då e	n->6	
då f	a->1	i->2	o->1	r->4	å->2	ö->4	
då g	e->3	ö->1	
då h	a->6	e->1	
då i	 ->5	d->1	n->10	
då j	a->2	u->1	
då k	a->10	o->4	v->1	
då l	a->1	
då m	a->2	e->3	y->1	å->2	ö->1	
då o	c->7	e->1	l->1	m->2	
då p	e->1	o->1	r->1	å->1	
då r	i->1	ä->3	
då s	e->1	j->1	k->7	n->1	o->3	ä->2	å->1	
då t	a->4	i->4	r->1	v->1	y->1	ä->1	
då u	n->3	p->2	
då v	a->1	e->3	i->9	r->1	
då ä	n->1	r->2	v->1	
då ö	v->1	
då, 	f->1	m->1	n->1	
då..	.->1	
då.D	e->1	
då?I	n->1	
dåli	g->19	
dåtg	ä->6	
dåva	r->1	
dé -	 ->1	
dé a	t->2	
dé j	a->1	
dé k	o->1	
dé o	m->1	
dé s	o->3	
dé ä	r->1	
dé, 	m->1	
dée,	 ->1	
déer	 ->6	,->1	n->1	
dén 	a->6	b->3	m->1	o->3	v->1	
dén,	 ->1	
dö i	 ->1	
död 	i->1	o->2	v->2	
död.	A->1	J->1	M->1	
döda	 ->1	"->1	,->1	d->3	n->1	s->2	t->1	
dödf	ö->1	
döds	d->1	f->1	
döen	d->1	
dölj	a->6	e->3	s->1	
döma	 ->26	,->1	.->1	n->7	s->2	
dömb	a->1	
dömd	,->1	e->2	
döme	.->1	r->9	s->1	
döml	i->2	
dömn	i->28	
döms	 ->3	
dömt	 ->4	s->1	
döpa	 ->1	
döpe	r->2	
döpt	e->1	
dör 	M->1	e->1	f->1	m->1	u->1	
dörr	 ->1	,->1	a->3	e->4	
döst	r->1	
dött	.->2	r->1	
dövt	 ->1	
e "a	l->1	v->1	
e "d	e->1	
e "f	ö->1	
e "k	o->2	
e "l	ä->2	
e "s	v->1	
e (A	5->29	
e (B	e->1	
e (C	5->2	
e (K	u->2	
e (a	r->1	
e (f	i->1	
e (m	a->1	
e - 	,->1	a->5	d->4	e->2	f->2	h->2	i->1	j->3	k->1	m->1	n->3	o->4	p->2	s->5	t->1	u->2	v->1	ä->2	
e -,	 ->1	
e 10	0->1	
e 11	 ->1	5->1	
e 12	 ->1	
e 14	 ->4	
e 15	 ->3	
e 18	 ->1	
e 19	5->1	9->4	
e 20	 ->1	0->1	
e 21	 ->1	
e 25	 ->4	
e 26	 ->1	
e 35	 ->1	
e 4,	 ->1	
e 40	 ->1	
e 41	 ->1	
e 8 	t->1	
e 9 	m->1	
e Ah	e->1	
e Al	t->2	
e Am	s->3	
e B 	t->1	
e BN	P->1	
e Ba	n->1	r->1	
e Be	r->1	s->1	
e Bu	s->1	
e Ce	n->2	
e Cu	r->1	
e Da	n->1	
e De	 ->1	
e Di	r->1	
e Du	i->1	
e EM	U->1	
e EU	 ->1	-->2	:->1	
e Ek	o->1	
e Eu	r->23	
e FN	:->1	
e Fo	U->1	r->1	
e Fr	a->2	
e Fu	n->1	
e Ga	m->1	r->2	
e Gr	a->2	o->1	ö->1	
e Ha	i->1	
e He	d->1	
e Hi	t->1	
e Ho	l->1	
e Im	b->1	
e Ir	l->1	
e Is	r->1	
e It	a->1	
e Ja	c->1	
e Jo	n->1	
e Ka	r->2	
e Ki	n->3	
e Ko	c->2	u->1	
e La	n->1	
e Lo	y->1	
e Ma	r->4	
e Me	l->1	
e Na	p->1	t->1	
e OL	A->1	
e Oi	l->1	
e Ou	v->1	
e Pa	l->7	
e Pl	a->1	
e Pr	o->15	
e Qu	e->1	
e Ra	p->1	
e Re	p->1	
e Ro	m->2	o->1	y->1	
e Sa	n->1	
e Sc	h->2	
e Se	i->1	
e Sv	e->1	
e Sw	o->1	
e Tr	i->1	
e Tu	r->1	
e Va	t->1	
e Ve	n->1	
e We	b->1	
e ab	s->2	
e ac	c->11	
e ad	 ->1	j->1	m->5	
e af	f->1	
e ag	e->4	
e ai	d->1	
e ak	t->10	
e al	b->2	l->78	t->1	
e am	b->2	e->3	
e an	 ->2	a->7	b->1	d->14	f->1	g->7	i->1	l->6	m->4	n->1	o->1	p->3	s->51	t->16	v->9	
e ap	p->2	
e ar	a->3	b->21	g->2	t->3	
e as	p->3	t->1	y->1	
e at	t->241	
e au	t->4	
e av	 ->203	.->1	d->1	f->4	g->6	r->1	s->7	t->6	v->3	
e ba	k->2	l->1	n->3	r->101	s->3	
e be	a->3	d->9	f->15	g->14	h->31	i->1	k->5	l->3	r->13	s->41	t->44	v->9	
e bi	d->6	f->1	l->18	n->1	o->2	s->2	
e bl	a->6	e->1	i->40	u->2	
e bo	k->1	r->5	v->1	
e br	a->2	e->2	i->8	o->6	ä->1	
e bu	d->3	r->1	
e by	g->3	r->7	t->1	
e bä	r->2	s->5	t->2	
e bå	d->7	t->4	
e bé	b->1	
e bö	r->18	
e ce	n->4	
e ch	a->1	e->3	
e ci	v->1	
e co	n->2	
e da	g->18	m->3	n->4	t->1	
e de	 ->37	b->7	c->4	f->1	g->1	l->27	m->16	n->84	p->1	r->1	s->12	t->106	
e di	a->1	e->1	p->1	r->9	s->13	t->1	
e dj	ä->1	
e do	c->10	g->1	m->4	
e dr	a->13	o->1	y->1	ö->2	
e du	s->1	
e dy	k->2	
e dä	r->36	
e då	 ->11	.->1	
e dö	l->1	m->1	r->1	
e ef	f->3	t->12	
e eg	e->4	n->2	
e ej	 ->1	
e ek	o->27	
e el	-->1	e->3	i->1	l->18	m->1	
e em	e->2	o->3	
e en	 ->70	b->9	d->18	e->4	g->4	h->3	i->1	l->4	o->4	s->22	t->2	
e ep	o->2	
e er	 ->11	.->1	a->1	b->2	f->2	i->1	k->4	s->1	
e et	a->1	n->2	t->49	
e eu	r->65	
e ev	e->3	
e ex	 ->1	a->4	e->3	i->2	p->16	t->2	
e fa	c->2	k->9	l->19	m->3	n->7	r->13	s->9	t->7	x->1	
e fe	l->1	m->12	
e fi	c->4	l->1	n->48	s->4	
e fj	o->3	ä->1	
e fl	a->4	e->29	y->2	
e fo	l->5	n->1	r->29	
e fr	a->44	e->5	i->12	u->5	ä->9	å->98	
e fu	l->1	n->12	t->1	
e fy	r->11	
e fä	s->2	
e få	 ->28	r->25	t->5	
e fö	l->5	r->401	
e ga	m->6	n->1	r->10	v->3	
e ge	 ->12	m->11	n->36	o->2	r->6	t->2	
e gi	l->1	v->2	
e gj	o->8	
e gl	ö->11	
e go	d->21	t->1	
e gr	a->10	u->27	ä->8	å->1	ö->9	
e gä	l->11	r->5	
e gå	 ->11	n->11	r->8	t->2	
e gö	m->1	r->41	
e ha	 ->37	d->13	f->4	l->4	m->1	n->31	r->157	
e he	l->55	m->6	n->1	r->4	t->1	
e hi	e->1	n->6	s->2	t->4	
e hj	ä->6	
e ho	n->5	p->2	r->1	s->4	t->3	
e hu	r->10	v->1	
e hy	c->1	s->1	
e hä	n->8	r->21	v->1	
e hå	l->10	r->2	
e hö	g->8	j->1	l->1	r->7	
e i 	A->1	B->2	D->2	E->8	F->2	H->2	I->2	K->4	L->1	S->2	T->1	a->11	b->4	d->40	e->11	f->21	g->7	h->6	k->11	l->2	m->9	n->8	o->3	p->5	r->4	s->31	t->9	u->11	v->6	y->2	z->1	Ö->2	ä->1	å->5	
e ia	k->2	
e ic	k->8	
e id	e->1	é->3	
e if	r->4	
e ig	e->1	n->1	
e il	l->1	
e im	p->1	
e in	b->7	d->8	f->23	g->15	i->3	k->1	l->9	n->23	o->13	r->11	s->29	t->92	v->8	
e is	o->1	r->3	
e it	a->6	
e ja	g->73	
e je	t->1	
e jo	r->5	u->2	
e ju	 ->3	d->1	r->1	s->4	
e jä	m->4	
e ka	m->3	n->115	p->2	r->1	t->11	
e ke	m->1	
e ki	n->5	
e kl	a->9	i->1	
e kn	a->2	ä->1	
e ko	l->19	m->152	n->49	r->3	s->8	
e kr	a->11	e->1	i->10	o->1	y->1	ä->12	
e ku	l->5	n->109	s->2	
e kv	a->8	i->2	ä->1	
e kä	l->1	n->9	r->1	
e kö	r->1	
e la	 ->1	d->1	g->15	n->35	s->2	
e le	d->22	g->2	t->1	v->4	
e li	b->5	d->2	g->7	k->1	n->1	v->4	
e lo	g->3	k->8	
e lu	r->1	
e ly	c->8	s->2	
e lä	c->1	g->8	m->6	n->42	r->2	t->5	
e lå	n->5	s->1	t->7	
e lö	f->1	n->1	p->1	s->7	
e ma	j->6	k->9	n->38	r->75	t->1	x->1	
e me	d->158	k->3	l->14	n->5	r->10	s->22	t->3	
e mi	g->7	l->16	n->34	s->9	t->1	
e mo	b->1	d->2	n->1	t->16	
e mu	l->4	
e my	c->22	l->1	n->7	
e mä	k->2	n->33	r->3	
e må	l->18	n->39	s->32	
e mö	j->12	r->1	t->1	
e na	t->56	
e ne	d->2	g->2	k->1	
e ni	 ->7	o->7	v->4	
e no	g->3	r->12	t->4	
e nu	 ->13	v->8	
e ny	a->23	h->3	l->1	s->4	t->1	
e nä	m->7	r->35	s->3	t->1	
e nå	 ->1	g->40	r->1	
e nö	d->7	j->8	
e oa	v->1	
e ob	e->4	
e oc	h->224	k->58	
e oe	r->1	
e of	a->1	f->13	r->1	t->1	
e ol	a->1	i->45	j->3	o->1	y->7	ä->1	
e om	 ->116	,->3	.->1	b->2	e->2	f->7	k->1	p->1	r->36	s->3	ö->1	
e on	s->2	
e op	e->1	i->1	p->1	r->1	
e or	d->26	g->6	i->1	k->1	o->6	s->3	ä->1	
e os	s->14	
e ot	i->1	
e ov	a->2	e->1	i->1	ä->1	
e pa	l->3	r->38	s->1	
e pe	k->4	l->2	n->5	r->39	s->1	
e pi	l->1	
e pl	a->9	i->1	
e po	l->35	p->1	r->2	s->5	t->1	
e pr	a->3	e->13	i->26	o->48	
e pu	b->2	n->14	
e på	 ->176	,->2	b->2	g->4	m->1	p->5	s->3	
e qu	a->2	
e ra	d->1	m->8	p->10	s->3	t->1	
e re	a->9	d->10	f->17	g->81	k->2	l->2	n->4	p->1	s->31	v->3	
e ri	k->24	s->5	
e ro	l->9	s->1	t->1	
e ru	b->2	l->1	n->1	t->1	
e ry	k->1	
e rä	c->8	d->1	k->4	t->50	
e rå	d->23	
e rö	r->3	s->3	
e sa	d->2	g->5	k->6	m->31	n->6	t->1	
e se	 ->16	d->14	k->4	n->40	r->4	s->4	t->3	x->3	
e si	f->2	g->31	k->1	n->2	s->4	t->11	
e sj	u->2	ä->11	
e sk	a->71	e->10	i->4	j->5	o->2	r->2	u->29	y->7	ä->6	å->2	ö->1	
e sl	a->1	i->1	u->8	ä->1	
e sm	å->22	
e sn	a->12	
e so	c->13	m->213	p->1	r->2	
e sp	a->1	e->5	r->2	ä->1	å->2	
e st	a->35	e->3	i->1	o->29	r->22	y->4	ä->11	å->15	ö->28	
e su	m->2	n->1	v->2	
e sv	a->9	e->1	å->7	
e sy	f->6	m->1	n->6	r->1	s->23	
e sä	g->18	k->15	l->1	m->4	n->2	r->3	t->29	
e så	 ->21	d->1	l->9	r->1	
e sö	k->1	n->1	r->3	
e t.	e->1	o->1	
e ta	 ->34	c->2	g->8	k->1	l->29	n->5	r->5	s->3	x->2	
e te	c->1	k->6	n->1	r->1	x->3	
e ti	d->33	l->216	o->5	s->1	t->4	
e tj	a->1	ä->12	
e to	g->2	l->4	p->1	t->3	
e tr	a->8	e->13	o->9	ä->2	
e tu	m->3	n->1	r->3	s->1	
e tv	e->2	i->4	ä->4	å->22	
e ty	c->3	d->4	n->1	s->3	v->1	
e tä	c->6	n->3	
e ul	t->1	
e un	d->34	i->4	
e up	p->80	
e ur	a->4	b->1	h->2	s->1	v->1	
e ut	 ->9	,->2	?->1	a->17	b->6	e->3	f->5	g->16	k->2	l->3	m->3	n->3	o->1	r->7	s->10	t->19	v->33	ö->5	
e va	c->1	d->15	l->7	n->3	r->131	t->11	
e ve	c->11	l->3	m->1	r->23	t->15	
e vi	 ->99	,->1	a->1	d->15	k->27	l->104	n->2	r->2	s->11	t->1	
e vo	l->2	n->2	r->4	
e vr	a->1	
e vä	c->1	g->3	l->5	n->9	r->15	s->3	x->1	
e vå	n->1	r->7	
e yr	k->3	
e yt	t->11	
e Ös	t->1	
e äg	n->2	t->2	
e äl	d->1	
e äm	n->1	
e än	 ->49	.->1	d->27	n->5	t->4	
e är	 ->160	.->1	e->2	
e äv	e->9	
e å 	r->1	
e åk	l->1	
e ål	ä->1	
e år	 ->14	.->7	e->28	h->1	s->1	t->1	
e ås	i->3	t->2	
e åt	 ->5	a->8	e->16	f->3	g->42	m->1	t->1	
e öa	r->1	
e ök	a->5	n->2	
e öm	m->1	
e ön	s->11	
e öp	p->11	
e ös	t->3	
e öv	e->52	n->1	r->12	
e! J	a->5	
e! N	i->2	
e!Al	l->1	
e!De	t->1	
e!Ja	g->1	
e!Me	n->1	
e!Ni	 ->1	
e!Sk	a->1	
e!Äv	e->1	
e" s	k->1	o->1	
e", 	i->1	o->2	
e(A5	-->1	
e) f	ö->1	
e) i	 ->1	
e) o	c->1	
e, ,	 ->1	
e, A	l->1	
e, B	e->1	
e, D	a->2	i->1	
e, E	r->2	
e, F	r->1	ö->1	
e, G	r->1	
e, H	a->1	
e, L	e->1	i->1	
e, R	a->1	
e, S	p->1	
e, a	l->1	n->1	r->1	t->15	v->2	
e, b	e->2	l->1	o->3	r->1	y->1	ä->1	å->3	ö->1	
e, d	e->19	v->2	ä->2	å->1	
e, e	f->7	m->1	n->3	t->1	x->1	
e, f	i->1	r->4	ö->10	
e, g	a->1	e->1	ö->1	
e, h	a->7	e->10	u->3	ö->1	
e, i	 ->11	n->13	
e, j	a->4	
e, k	a->5	i->1	o->6	r->1	ä->1	
e, l	i->3	
e, m	e->25	i->1	o->1	u->1	y->1	å->1	
e, n	a->2	y->1	ä->10	å->1	ö->1	
e, o	a->1	c->39	m->6	s->2	
e, p	r->5	å->5	
e, r	ö->1	
e, s	a->2	k->5	o->19	ä->3	å->4	
e, t	a->1	i->1	o->1	r->1	y->3	ä->1	å->1	
e, u	n->2	r->1	t->5	
e, v	a->6	e->1	i->18	ä->1	å->4	
e, ä	n->1	r->10	
e, å	t->4	
e, ö	k->1	
e- o	c->6	
e- p	r->1	
e-Al	p->1	
e-Ar	d->1	
e-At	l->1	
e-Fr	a->2	
e-Le	 ->1	
e-Lo	i->1	
e-Ma	n->1	
e-No	r->1	
e-al	b->1	
e-av	t->2	v->1	
e-da	n->1	
e-de	-->2	
e-di	s->2	
e-fa	l->1	
e-fo	s->1	
e-fö	r->1	
e-lo	b->1	
e-lä	n->1	
e-ma	i->1	
e-me	t->1	
e-pr	o->2	
e-sp	r->3	
e-st	a->9	i->1	o->1	
e. D	e->5	ä->1	
e. M	e->1	
e. O	c->1	m->1	
e. V	i->2	
e. Ä	n->1	
e.- 	(->1	F->1	
e.. 	(->1	P->1	V->1	
e..(	E->1	
e...	)->1	
e.Ak	t->1	
e.Al	l->2	
e.An	n->1	
e.At	t->2	
e.Av	 ->1	s->2	
e.Be	s->1	t->1	
e.Bå	d->1	
e.De	 ->1	n->9	r->1	s->6	t->66	
e.Dä	r->8	
e.Då	 ->2	
e.Ef	t->5	
e.Em	e->1	
e.En	 ->5	d->1	l->2	
e.Et	t->1	
e.Eu	r->4	
e.FP	Ö->1	
e.Fr	u->4	å->1	
e.Fö	r->15	
e.Ge	n->2	
e.Gr	u->1	
e.Ha	n->2	
e.He	l->1	r->12	
e.Ho	n->1	
e.Hu	r->1	v->4	
e.I 	E->1	d->3	o->1	s->2	v->2	
e.Id	é->1	
e.Im	m->1	
e.In	f->1	o->1	
e.Ja	g->60	
e.Ka	n->2	
e.Ko	m->7	
e.Li	k->2	
e.Ly	c->1	
e.Lä	g->1	
e.Lå	t->4	
e.Ma	l->1	n->7	
e.Me	d->2	n->16	r->1	
e.Mi	n->7	
e.Må	n->1	
e.Ni	 ->4	
e.Nu	 ->2	
e.Nä	r->3	
e.Oc	h->3	
e.Of	f->1	
e.Om	 ->7	
e.Pa	r->1	
e.Pl	a->1	
e.Po	r->1	
e.Pr	o->2	
e.På	 ->2	
e.Re	f->1	s->1	
e.Ro	t->1	
e.Rå	d->2	
e.Sa	m->1	v->1	
e.Sc	h->1	
e.Se	d->1	
e.Sk	a->1	
e.Sl	u->2	
e.So	m->8	
e.St	ä->1	ö->1	
e.Så	 ->2	l->1	
e.TV	-->1	
e.Ta	 ->1	c->3	
e.Ti	l->3	
e.To	p->1	
e.Tr	a->1	o->2	
e.Tv	ä->1	
e.Un	d->2	
e.Up	p->1	
e.Ur	 ->1	
e.Va	d->3	r->3	
e.Vi	 ->23	d->2	n->1	t->1	
e.Vå	r->3	
e.d.	,->1	
e.Än	d->2	
e.Är	 ->1	
e.Äv	e->2	
e.Å 	a->1	
e.År	 ->1	
e.Åt	e->1	g->1	
e.Ös	t->1	
e: "	A->1	v->1	
e: A	n->1	r->2	
e: D	e->2	
e: F	l->1	r->1	ö->1	
e: G	e->2	r->1	
e: H	a->1	
e: I	 ->1	
e: J	a->1	o->1	
e: K	o->2	ä->1	
e: M	a->1	
e: N	a->1	y->1	ä->1	
e: P	o->1	
e: S	t->2	
e: T	u->1	
e: U	t->1	
e: V	a->2	i->2	
e: b	a->1	e->1	
e: d	e->1	
e: f	ö->1	
e: h	u->1	
e: i	 ->2	
e: k	o->1	
e: t	o->1	
e: u	t->1	
e: v	a->1	
e: Å	t->2	
e; d	e->2	
e; h	ä->1	
e; j	a->1	
e; m	i->1	
e; p	u->1	
e?De	n->1	t->1	
e?En	l->1	
e?Fö	r->2	
e?He	m->1	r->3	
e?Hu	r->1	
e?Hä	r->1	
e?I 	f->1	
e?Ja	g->1	
e?Ka	n->1	
e?Oc	h->1	
e?So	m->1	
e?Vi	 ->1	l->1	
eEn 	v->1	
eFru	 ->1	
eHer	r->1	
eNäs	t->2	
ePro	t->1	
ea b	e->1	
ea o	c->3	
ead-	k->1	
eade	r->5	
eadi	n->1	
eadl	i->1	
eage	r->16	
eake	,->1	
eakt	 ->1	a->30	i->12	o->10	
eal 	p->1	
eal,	 ->2	
eala	 ->1	
eale	n->1	t->1	
eali	s->10	t->7	
eami	n->8	
ean-	C->1	
eanu	t->1	
earb	e->3	
earv	e->1	
eate	r->1	
eati	v->2	
eato	 ->8	.->1	b->1	n->1	s->11	
eatt	l->4	
eatö	r->1	
eau 	d->1	f->1	
eau"	,->1	
eau,	 ->2	
eaux	,->1	
eb, 	s->1	
ebal	l->1	
eban	o->1	
ebar	 ->1	
ebas	e->1	t->1	
ebat	t->170	
ebbe	l->1	
ebbp	l->1	
ebef	o->2	r->1	
ebeh	a->1	
eben	g->1	
ebes	t->3	ö->1	
ebet	a->12	
ebil	d->1	
eboa	r->1	
eboe	l->1	n->1	
ebol	a->4	
ebor	g->1	
ebre	i->1	
ebro	n->1	
ebru	a->16	
ebrå	s->2	
ebrö	d->1	
ebud	 ->6	,->2	e->1	
ebyg	d->1	g->24	
ebäl	t->10	
ebän	k->1	
ebär	 ->90	,->1	.->2	a->15	
ebåd	a->1	
ebör	d->7	s->1	
ec l	'->1	
eced	o->1	
ecem	b->19	
ecen	n->7	t->15	
ecia	l->14	
ecie	l->42	
ecif	i->29	
ecir	k->1	
ecis	 ->36	a->1	e->11	t->1	
eck 	h->1	i->1	ä->1	
ecka	 ->6	.->1	n->17	
ecke	n->15	
eckl	a->73	i->175	
eckn	a->29	i->3	
ecko	r->17	
ecov	e->1	
ectn	e->1	
ecu 	m->1	
ecu,	 ->1	
ecyc	l->1	
ed "	a->2	e->1	
ed (	a->1	
ed -	 ->1	
ed 1	2->1	3->2	4->1	6->1	9->1	
ed 2	 ->2	0->2	4->1	7->2	8->1	
ed 3	0->1	6->1	
ed 5	 ->1	
ed 8	0->1	
ed A	.->1	m->2	
ed B	S->1	a->1	
ed D	a->2	
ed E	-->1	D->1	U->1	r->4	u->12	
ed F	r->4	
ed G	A->1	
ed H	a->4	
ed I	n->1	s->2	
ed J	ö->1	
ed K	o->2	
ed L	e->1	i->2	
ed M	a->3	i->1	
ed O	L->1	s->1	
ed P	a->1	
ed R	y->1	
ed S	a->1	y->4	
ed T	h->1	u->2	
ed U	S->4	
ed V	a->1	e->1	
ed a	d->1	l->34	n->28	r->12	t->106	u->2	v->17	
ed b	a->3	e->7	i->5	r->7	u->1	å->1	
ed d	a->4	e->246	i->8	r->2	u->2	y->2	
ed e	f->2	k->1	l->1	n->89	r->13	t->29	u->2	x->5	
ed f	a->4	e->1	i->1	l->3	o->3	r->30	u->9	å->1	ö->39	
ed g	a->1	e->7	i->1	l->2	o->5	r->4	
ed h	a->3	e->3	j->25	o->1	u->5	ä->18	å->1	ö->2	
ed i	 ->27	f->1	m->1	n->23	s->2	
ed j	o->1	u->1	ä->1	
ed k	a->5	i->1	l->1	n->1	o->31	r->7	u->1	v->9	ä->1	ö->1	
ed l	a->3	e->2	i->8	ä->1	ö->2	
ed m	a->6	e->15	i->30	o->5	y->6	å->7	ö->4	
ed n	a->13	e->3	u->3	y->4	ä->1	å->8	ö->7	
ed o	c->18	f->1	j->1	l->2	m->23	r->6	s->8	
ed p	a->13	e->5	l->1	o->3	r->8	s->1	u->2	å->19	
ed r	a->1	e->19	i->2	ä->10	å->5	ö->1	
ed s	.->1	a->10	e->1	i->26	j->1	k->7	l->2	m->1	n->1	o->7	p->5	t->37	u->2	v->2	y->2	ä->9	å->11	
ed t	.->1	a->43	e->2	i->22	o->1	r->6	u->2	v->5	y->1	ä->1	
ed u	n->6	p->6	r->1	t->17	
ed v	a->13	e->6	i->17	ä->1	å->17	
ed y	r->1	t->4	
ed Ö	V->1	s->1	
ed ä	n->4	r->5	
ed å	r->2	t->4	
ed ö	k->1	m->1	p->1	s->1	v->11	
ed, 	a->1	d->2	e->1	f->1	g->1	m->2	n->1	o->3	p->1	s->1	v->1	
ed.D	e->4	ä->1	
ed.E	f->1	
ed.F	ö->1	
ed.H	e->1	u->1	
ed.I	 ->1	
ed.J	a->1	
ed.K	o->1	
ed.V	i->2	
eda 	E->1	a->3	d->5	e->8	f->6	h->1	i->2	m->4	o->4	p->4	s->2	t->30	u->3	å->1	
eda,	 ->3	
edag	o->1	
edak	t->1	
edam	o->74	ö->84	
edan	 ->283	,->11	.->10	?->2	d->18	s->3	
edar	b->2	e->13	f->1	n->8	s->1	
edas	 ->6	,->1	t->1	
edat	 ->1	
edbe	s->16	
edbo	r->170	
edbr	o->1	
edd 	a->16	f->2	t->3	u->2	ä->1	
edda	 ->18	.->1	
edde	 ->14	,->1	l->59	n->2	s->7	
ede 	g->1	o->1	ä->1	
ede.	R->1	
edel	 ->61	,->12	.->9	?->1	a->4	b->18	h->3	l->4	p->2	s->121	t->1	
eden	 ->1	,->1	s->1	
edep	a->2	
eder	 ->48	,->2	a->12	b->11	g->1	i->2	l->18	s->1	t->1	v->1	
edes	 ->44	
edet	 ->3	
edfi	n->2	
edfö	r->20	
edga	t->1	
edge	 ->4	r->10	s->5	t->1	
edgi	v->2	
edgå	n->2	
edgö	r->2	
edhj	ä->1	
edi 	-->1	
edi.	D->1	
edia	 ->5	l->1	s->1	t->1	
edic	i->1	
edie	n->2	r->7	
edig	e->1	h->1	n->1	
edin	f->1	g->8	
edit	e->2	i->1	
edja	 ->1	n->2	
edje	 ->56	,->4	:->1	d->6	l->6	
edjo	r->1	
edkv	i->1	
edkä	n->5	
edla	 ->2	g->1	r->1	
edle	m->343	n->12	t->1	
edli	d->2	g->10	n->2	
edlä	g->4	
edmo	n->3	
edni	n->83	
edo 	a->4	
edof	i->1	
edog	j->1	ö->9	
edom	 ->2	,->2	a->4	e->4	
edov	i->4	
edra	 ->5	d->1	g->160	n->3	r->3	
edre	v->1	
edri	v->15	
edro	g->1	
edru	s->1	
edrä	g->37	
eds 	a->1	b->1	i->1	m->1	r->1	s->1	u->1	å->1	
eds,	 ->1	
eds.	J->1	
edsa	n->1	v->3	
edsb	e->2	
edse	n->2	
edsf	ö->3	
edsk	a->2	r->1	ä->3	
edsp	a->1	r->22	
edss	a->4	t->24	
edst	j->2	ä->3	
edsu	p->1	
edt 	o->2	
edt,	 ->2	
edte	r->14	
educ	e->4	
edur	r->1	
edve	r->19	t->42	
edvr	i->12	
edvä	r->1	
edöm	a->15	b->1	d->1	e->4	l->2	n->28	s->3	t->1	
ee-f	ö->1	
ee-l	o->1	
ee.D	e->1	
eela	n->2	
eell	 ->1	.->1	a->4	
eend	e->63	
eenh	e->5	
eer 	o->1	s->2	
eer,	 ->4	
eerJ	a->1	
eerb	e->3	
eeri	n->1	
eers	 ->3	ä->2	
ees 	W->1	
eexe	m->1	
ef h	a->1	
efad	e->1	
efal	l->20	
efan	t->1	
efar	a->5	
efat	t->12	
efel	 ->1	
efen	 ->1	
efer	 ->4	,->2	.->1	e->7	n->8	
effe	k->148	
effi	c->1	
efin	g->1	i->36	n->31	t->10	
efit	-->5	
efle	k->7	
eflä	c->1	
efog	a->5	e->27	
efol	k->43	
efon	,->1	d->1	
efor	d->8	m->141	
efra	k->10	
efri	a->4	e->6	h->2	
efrä	m->1	
efrå	g->2	
efte	r->373	
eful	l->18	
efus	e->1	i->1	
efäl	h->1	
efän	g->1	
efär	 ->9	l->1	
efäs	t->10	
eföl	l->1	
eför	b->1	e->6	f->8	h->3	k->1	o->1	s->1	v->1	
eg a	t->1	
eg b	o->1	
eg f	r->6	ö->5	
eg g	j->1	
eg h	a->1	ä->1	
eg i	 ->13	
eg j	ä->1	
eg l	ä->2	
eg m	o->4	
eg n	ä->2	
eg o	c->2	
eg p	å->3	
eg s	o->7	
eg t	e->1	i->3	
eg u	n->1	
eg v	i->1	
eg, 	d->1	o->1	u->1	
eg.D	e->2	
ega 	B->3	E->2	F->6	H->1	J->3	K->1	L->1	M->1	N->2	R->2	S->1	a->1	b->1	d->1	f->2	k->1	s->2	t->1	v->4	
ega!	 ->1	D->1	J->1	Ä->1	
ega,	 ->3	
ega.	J->1	
egad	.->1	e->1	
egag	n->4	
egal	 ->4	a->7	i->2	t->9	
egan	 ->16	
egap	r->1	
egas	 ->2	
egat	 ->3	i->42	
egdr	a->1	
ege.	O->1	
ege?	H->1	
egel	 ->3	b->16	m->2	n->6	r->2	s->2	v->19	
egem	e->3	
egen	 ->34	a->1	d->5	e->1	f->5	s->22	t->43	
eger	 ->36	!->65	,->14	.->5	:->1	a->4	i->288	n->9	s->1	
eget	 ->24	,->2	.->1	
egi 	f->5	h->1	i->1	k->1	m->1	o->2	s->4	t->2	
egi,	 ->4	
egi.	D->1	F->1	J->1	
egic	k->1	
egie	r->17	t->2	
egim	e->3	
egin	 ->5	.->2	s->1	
egio	n->252	
egip	l->1	
egis	k->17	t->20	
egit	i->18	
egiu	m->3	
egla	 ->7	d->2	r->13	s->2	
egle	r->126	
egli	n->1	
egna	 ->45	
egni	,->1	
egoi	s->2	
egor	 ->1	i->9	s->2	
egra	d->3	t->17	v->1	
egre	p->13	r->23	
egri	p->22	t->3	
egru	n->2	
egrä	n->68	
egur	o->1	
egär	 ->11	.->1	a->34	d->3	s->1	t->10	
egå 	e->1	s->1	
egåe	n->15	
egån	g->4	
egår	 ->3	
egås	 ->3	
egåt	t->3	
ehab	i->1	
ehag	l->2	
ehan	d->88	
ehar	 ->2	
ehav	a->2	
ehin	d->1	
ehov	 ->23	,->2	.->3	e->39	
ehre	n->7	
ehäf	t->1	
ehål	l->120	
ehöj	a->1	
ehöl	l->5	
ehör	i->18	
ehöv	a->16	d->2	e->99	s->27	t->3	
eido	s->2	
eijs	 ->1	.->1	
eik.	D->1	
eikh	 ->1	-->1	.->2	
eill	e->1	
ein.	J->1	
einc	i->1	
eind	r->2	u->1	
eine	n->6	
eins	p->1	t->2	
einz	 ->2	
eira	 ->2	,->2	.->1	
eise	r->2	
eisk	 ->102	.->1	a->586	e->2	t->20	
eism	i->2	
eivr	a->1	
eixa	s->5	
eiz,	 ->1	
ej a	n->1	t->1	v->1	
ej b	e->2	o->1	
ej i	 ->1	
ej k	o->1	
ej l	å->1	ö->1	
ej n	ä->1	
ej t	i->1	
ej ä	r->1	
ej, 	b->2	d->1	h->1	j->1	m->2	n->1	s->2	
ej.(	A->1	
ej.E	x->1	
ej.I	 ->1	
ej.R	å->1	
ejda	 ->1	s->1	t->1	
ejdo	s->1	
ejor	d->3	
ejud	i->4	
ejäl	t->3	
ek h	o->1	
ek o	s->1	
ek s	o->1	
eka 	B->1	a->9	d->4	f->5	p->6	r->1	v->1	
eka,	 ->2	
eka.	D->1	M->1	
ekad	 ->1	e->11	
ekan	 ->14	,->1	d->11	i->10	t->3	
ekar	 ->16	,->1	
ekas	 ->5	,->1	t->1	
ekat	 ->11	,->4	.->1	
ekel	 ->2	,->1	s->1	
eken	 ->2	,->1	s->1	
eker	 ->1	n->1	
ekhe	t->4	
ekin	g->1	
ekis	k->6	t->2	
ekla	g->42	m->2	n->15	
ekle	r->1	t->1	
eklö	s->1	
ekni	k->13	s->36	
ekno	l->3	
ekod	 ->5	e->3	
ekok	a->1	
ekol	l->1	o->14	
ekom	 ->2	m->68	p->1	s->1	
ekon	 ->1	c->1	f->2	o->283	s->3	v->1	
ekor	d->2	t->1	
ekos	t->1	y->4	
ekre	t->16	
ekri	s->1	
ekry	t->1	
ekrä	f->30	
eksa	k->1	m->5	
ekt 	a->8	b->6	d->1	e->3	f->28	g->1	h->3	i->3	k->4	l->2	m->7	n->1	o->5	p->3	s->23	t->8	u->3	v->3	ä->1	
ekt"	,->1	
ekt,	 ->8	
ekt.	D->4	F->2	I->1	J->1	M->2	S->1	U->1	
ekt:	 ->1	
ekt;	 ->1	
ekt?	T->1	U->1	
ekta	 ->10	.->1	b->3	d->2	k->3	r->2	
ekte	n->38	r->79	t->14	
ekti	n->1	o->18	v->354	
ekto	r->107	
ektr	i->1	o->9	u->2	
ektu	e->3	
ekty	r->1	
ektö	r->7	
ekul	a->4	
ekun	d->3	
ekva	l->1	t->6	
ekve	n->62	
ekvo	t->1	
ekvä	m->16	
ekym	m->6	r->10	
ekäm	p->41	
ekän	n->1	
el (	k->2	
el -	 ->5	
el 1	 ->2	0->1	1->1	2->2	3->5	4->1	5->3	6->1	
el 2	.->2	2->1	5->4	8->5	9->2	
el 3	.->2	0->1	3->2	7->2	9->1	
el 4	 ->5	.->1	2->1	8->2	
el 5	 ->1	.->1	0->2	2->1	6->1	
el 6	 ->9	.->1	2->1	7->1	
el 7	 ->7	,->1	
el 8	1->10	2->2	7->2	8->2	
el 9	.->1	4->1	5->1	
el B	a->1	
el H	i->1	
el K	o->1	
el N	y->1	
el P	e->1	
el R	i->1	
el a	l->2	n->5	t->14	v->83	
el b	e->4	l->1	ä->1	ö->2	
el d	e->8	r->1	
el e	n->1	t->1	
el f	a->4	o->1	r->5	å->1	ö->28	
el g	a->1	e->3	ö->1	
el h	a->5	i->1	j->1	y->1	ä->2	
el i	 ->20	n->5	
el k	a->4	o->3	v->2	
el l	e->1	i->1	ö->2	
el m	a->1	e->8	å->2	
el n	i->2	u->1	y->1	ä->3	
el o	c->37	m->11	
el p	a->1	e->2	o->1	å->26	
el r	a->1	e->1	i->1	ä->1	ö->1	
el s	a->3	e->1	i->1	k->4	o->17	t->1	ä->3	å->1	
el t	i->7	o->1	r->1	
el u	n->3	p->1	r->1	t->2	
el v	a->2	e->2	i->2	
el ä	n->2	r->15	v->1	
el å	t->1	
el ö	v->1	
el! 	I->1	J->1	
el!M	e->1	
el!T	i->1	
el, 	A->1	a->3	d->3	e->4	f->2	i->2	j->1	k->3	l->2	m->7	n->3	o->10	s->5	u->1	v->4	ä->1	å->1	ö->1	
el- 	o->3	
el-I	)->1	I->1	
el-S	h->5	y->1	
el.B	e->1	
el.D	e->11	ä->1	
el.E	U->1	f->1	u->1	
el.F	r->1	
el.G	e->1	
el.I	 ->1	
el.J	a->4	
el.M	e->4	
el.N	ä->2	
el.S	a->1	c->1	å->1	
el.T	v->1	
el.V	i->10	
el.Ä	n->1	r->1	
el: 	E->1	F->1	U->1	V->1	d->1	
el; 	i->1	
el?E	l->1	
el?J	a->1	
ela 	9->1	B->1	E->19	K->1	M->1	S->1	a->8	b->2	d->20	e->13	f->8	g->3	h->2	i->6	k->11	l->2	m->2	n->1	o->3	p->2	r->4	s->6	t->11	u->9	v->6	å->3	
ela,	 ->1	
ela?	A->1	
elad	,->1	e->11	
elag	 ->1	d->5	
elak	t->24	
elan	d->57	
elar	 ->64	,->3	.->7	:->1	e->10	n->12	
elas	 ->7	,->2	.->1	p->1	t->10	
elat	 ->19	,->1	.->1	e->4	i->22	s->8	
elay	e->2	
elba	r->20	
elbe	r->1	
elbr	o->1	
elbu	n->15	
elby	r->1	
eled	a->2	
elef	a->1	o->1	
eleg	a->17	e->4	
elek	o->3	t->11	
elem	e->9	
elen	 ->25	"->1	,->8	.->3	F->2	ä->1	
eler	 ->1	.->1	n->5	s->3	
eles	 ->23	
elet	 ->1	
elev	a->9	e->1	i->1	
elfe	d->1	
elfr	å->3	
elft	e->1	
elfu	n->1	
elga	d->1	
elge	n->1	
elgi	e->9	s->8	v->1	
elha	v->3	
elhe	t->21	
elhj	ä->8	
elho	e->1	
elig	 ->1	?->1	a->2	e->1	g->26	h->2	i->4	t->5	
elik	e->1	
elil	l->1	
elim	i->6	
elin	j->1	
elis	k->15	
elkr	i->1	
elku	r->1	
elkv	o->1	
ell 	b->5	d->5	e->3	f->11	g->2	i->2	k->6	l->2	m->4	n->10	o->10	p->6	r->12	s->9	t->4	u->2	v->3	å->2	ö->3	
ell"	,->1	.->1	
ell,	 ->4	
ell-	 ->3	
ell.	A->1	D->3	F->1	J->1	M->1	S->1	V->1	Ä->1	
ella	 ->332	,->3	.->1	m->1	n->227	
ellb	e->1	i->1	
elle	k->3	n->3	r->443	
ellf	ö->3	
elli	 ->1	g->5	s->2	t->1	v->1	
ellm	y->1	
ellr	e->6	ä->4	
ells	k->1	
ellt	 ->108	,->6	.->1	;->1	
ellå	n->4	
ellö	s->2	
elma	j->1	s->1	
elme	d->1	
elms	h->1	
elmä	s->2	
eln 	"->1	f->3	i->1	k->1	m->1	o->2	t->5	ä->2	
eln,	 ->2	
eln.	D->1	
elni	n->42	
elns	 ->2	
elod	l->1	
elog	e->2	
elon	a->2	
elop	p->16	
elor	s->3	
elpl	a->1	
elpr	o->1	
elpu	n->2	
elra	p->1	
elre	g->4	
elri	k->1	
elro	l->1	
elru	m->1	
elry	c->1	
elrä	k->1	t->2	
els 	a->7	d->1	e->1	f->2	i->1	k->1	o->1	p->2	s->2	t->2	v->2	å->2	
els-	 ->1	
elsa	t->1	
elsd	r->1	
else	 ->125	,->12	-->1	.->20	a->1	b->1	f->11	h->1	k->2	l->3	m->1	n->53	o->1	r->172	u->1	v->2	x->1	
elsf	l->2	r->2	
elsh	a->1	i->1	
elsi	k->1	n->22	
elsk	-->1	a->7	i->1	o->2	r->4	t->1	v->1	y->1	
elsl	a->5	o->1	
elsm	y->9	ä->3	
elsn	y->1	
elso	m->2	n->5	r->3	
elsp	l->2	o->2	r->2	
elss	e->1	j->1	t->1	ä->43	
elst	 ->35	,->7	.->4	a->4	i->1	o->41	
elsu	t->3	
elsv	a->1	
elsy	n->1	s->2	
elsä	t->102	
elt 	-->1	E->1	a->12	b->1	d->3	e->27	f->12	g->3	h->2	i->10	k->24	l->2	m->4	n->7	o->28	p->3	r->11	s->15	t->5	u->4	v->3	ä->1	å->2	ö->3	
elt,	 ->1	
elt.	 ->1	D->3	E->1	H->2	I->1	J->1	U->1	V->2	
elt;	 ->1	
elt?	J->1	
elta	 ->15	,->2	g->30	r->9	
elti	d->2	s->1	
elto	g->2	
eltr	a->1	
eltä	c->4	
elut	b->2	
elux	,->1	
elva	 ->3	
elve	r->21	
elvi	s->40	
elvä	g->3	n->1	
elys	a->1	e->1	n->1	t->1	
elze	n->1	
eläg	e->20	g->5	n->6	
eläm	n->3	
elän	d->1	
elät	t->1	
elön	a->2	
elös	 ->1	a->1	t->2	
em -	 ->2	
em 2	0->1	
em a	l->2	n->1	t->5	v->6	
em b	e->3	
em d	a->1	e->6	i->1	ä->4	å->2	
em e	f->4	n->5	t->2	
em f	a->1	r->3	u->1	ö->29	
em g	r->2	å->1	ö->1	
em h	a->4	e->1	ä->1	
em i	 ->22	n->7	
em j	a->1	
em k	a->2	o->5	r->1	
em l	ä->2	
em m	e->23	o->1	y->1	å->2	ö->1	
em n	i->1	ä->3	å->1	
em o	c->23	m->3	
em p	u->2	å->11	
em r	e->1	
em s	e->1	k->5	o->101	t->1	å->1	
em t	i->6	
em u	r->1	t->4	
em v	a->2	e->2	i->4	
em ä	r->8	
em å	r->14	t->1	
em ö	v->2	
em, 	a->1	b->1	d->1	e->3	f->2	g->1	h->2	i->1	k->1	m->5	o->4	p->2	s->3	u->1	v->5	ä->1	å->1	
em. 	D->1	H->1	M->1	
em.(	A->1	
em..	 ->1	
em.A	l->1	v->1	
em.B	e->1	u->1	
em.D	e->12	ä->3	
em.E	n->1	u->1	
em.F	r->1	ö->2	
em.G	e->1	
em.H	e->5	
em.I	n->1	
em.J	a->7	
em.K	o->1	
em.M	a->1	e->3	å->1	
em.N	e->1	i->1	å->1	
em.O	m->1	
em.P	r->1	
em.R	e->1	
em.S	l->1	o->1	
em.T	y->1	
em.U	r->1	
em.V	e->1	i->8	
em: 	A->1	d->3	p->1	
em; 	d->2	
em?D	e->1	
em?M	e->1	
ema 	f->1	g->1	h->1	
ema,	 ->1	
emag	o->4	
emal	a->1	
eman	 ->3	.->1	g->17	n->3	
emar	k->1	
emas	k->1	
emat	 ->1	i->16	
emba	r->1	
embe	r->45	
embl	e->1	
embr	y->1	
embu	r->6	
emby	g->1	
emed	a->1	e->1	
emel	l->67	
emen	 ->25	,->4	.->1	i->5	s->390	t->32	
emes	t->4	
emet	 ->90	)->1	,->9	.->15	?->1	s->1	
emfö	r->1	
emhö	g->14	
emi,	 ->1	
emig	r->2	
emik	 ->1	a->5	
emin	a->1	i->4	s->1	
emis	-->1	k->2	m->5	s->1	t->6	
emit	i->3	
emiä	r->10	
emla	n->3	
emli	g->6	
emlä	n->1	s->1	x->1	
emlö	s->5	
emma	 ->9	,->1	:->1	p->1	r->14	
emme	t->1	
emog	r->3	
emok	r->137	
emom	r->3	
emon	s->6	t->8	
emot	 ->96	.->4	i->1	
empe	l->110	r->4	
empl	a->2	e->6	
empo	r->2	
empu	n->1	
ems 	a->2	t->1	
ems-	 ->1	
emsa	n->2	
emsk	 ->1	a->6	
emsl	a->9	ä->27	
emsr	e->1	
emss	t->284	
emt 	h->2	r->1	s->1	
emte	 ->14	d->2	
emti	e->1	o->2	
emto	n->5	
emvi	s->1	
emyn	d->1	
emän	 ->17	,->1	.->1	d->3	n->12	s->3	
emär	k->5	
emäs	s->1	
emål	 ->16	
emån	a->1	
emår	i->1	s->2	
emöd	a->3	
emöj	l->4	
emön	s->1	
emöt	a->4	e->1	s->2	
en "	E->1	L->1	T->2	d->2	e->2	h->1	n->1	r->2	s->1	å->1	
en (	1->3	B->2	E->1	F->1	I->1	K->1	e->1	i->1	m->1	o->1	s->1	
en ,	 ->1	
en -	 ->53	
en 1	 ->11	,->1	0->1	1->2	2->1	3->4	4->7	5->1	6->1	7->3	8->5	9->13	
en 2	 ->2	,->1	0->16	1->1	3->1	4->1	6->2	9->1	
en 3	 ->4	,->1	0->1	1->3	8->1	9->1	
en 4	 ->2	,->2	
en 5	 ->1	
en 6	 ->1	
en 7	 ->2	9->1	
en 9	 ->2	0->1	
en A	B->2	D->1	m->1	n->1	r->1	
en B	a->2	e->4	r->1	
en C	E->1	a->1	h->1	
en D	e->4	u->1	
en E	U->4	n->3	r->1	u->11	
en F	E->1	N->1	ö->1	
en G	a->1	r->3	
en H	a->1	
en I	 ->1	M->1	X->1	s->2	
en J	a->2	o->1	u->1	
en K	a->5	i->4	o->3	
en L	a->1	e->1	o->1	
en M	i->1	
en N	a->2	
en P	R->1	a->1	r->4	
en R	a->2	e->2	o->1	
en S	S->1	c->1	o->1	y->1	ã->1	
en T	h->1	o->1	y->3	
en U	n->2	
en V	i->1	
en W	o->1	
en X	X->1	
en a	b->2	c->4	d->8	g->2	k->10	l->48	m->4	n->179	r->19	s->7	t->270	u->3	v->482	x->1	
en b	a->23	e->153	i->20	l->25	o->19	r->41	u->9	y->8	ä->23	å->3	ö->28	
en c	e->9	h->7	o->6	
en d	a->22	e->283	i->24	j->6	o->10	r->7	u->3	y->1	ä->34	å->8	ö->9	
en e	f->42	g->16	j->1	k->49	l->32	n->132	p->1	r->8	t->21	u->142	v->4	x->19	
en f	a->24	e->8	i->27	j->7	l->7	o->25	r->178	u->20	y->2	ä->4	å->26	ö->576	
en g	a->26	e->139	i->6	j->11	l->11	n->2	o->24	r->46	u->1	y->1	ä->22	å->55	ö->14	
en h	a->250	e->31	i->5	j->5	o->23	u->11	y->2	ä->85	å->19	ö->27	
en i	 ->418	c->4	d->6	f->1	h->2	l->3	m->1	n->322	r->3	s->10	t->4	
en j	a->89	u->16	ä->6	
en k	a->108	e->2	i->1	l->17	n->1	o->234	r->35	u->24	v->7	ä->19	
en l	a->14	e->9	i->30	o->8	u->1	y->4	ä->22	å->24	ö->17	
en m	a->38	e->218	i->56	o->52	u->4	y->72	ä->18	å->107	ö->22	
en n	a->19	e->12	i->7	o->11	u->30	y->74	ä->42	å->18	ö->16	
en o	a->6	b->25	c->442	e->4	f->30	h->1	k->5	l->7	m->272	n->4	p->3	r->42	s->2	t->4	u->3	v->2	ä->1	ö->3	
en p	a->20	e->23	l->17	o->71	r->42	u->28	y->1	å->162	
en r	a->32	e->132	i->28	o->4	u->2	y->1	ä->48	å->9	é->1	ö->11	
en s	a->63	c->2	e->41	i->37	j->31	k->207	l->20	m->5	n->14	o->279	p->19	r->1	t->210	u->7	v->7	y->17	ä->25	å->73	ö->2	
en t	a->27	e->15	i->210	j->5	o->18	r->33	u->8	v->16	y->41	ä->4	
en u	n->64	p->50	r->9	t->90	
en v	a->60	e->43	i->240	o->3	ä->41	å->3	
en w	a->1	
en y	t->5	
en z	i->2	
en Ö	s->1	
en ä	g->2	l->1	n->43	r->212	v->16	
en å	 ->6	b->1	k->2	l->3	r->2	s->11	t->34	
en ö	d->1	k->30	m->1	n->4	p->6	r->1	s->18	v->55	
en! 	E->1	J->1	M->1	N->1	
en!N	ä->2	
en!R	ö->1	
en" 	a->1	e->1	i->1	o->1	s->1	
en",	 ->3	
en".	D->3	O->1	
en) 	(->1	f->1	h->1	z->1	
en)(	P->2	
en),	 ->1	
en).	D->1	H->1	
en)J	a->1	
en)N	ä->1	
en, 	"->1	1->4	8->1	A->2	B->4	C->1	E->2	I->2	J->1	K->2	L->1	N->1	P->3	R->1	S->2	T->2	V->2	W->1	a->18	b->17	d->49	e->33	f->65	g->4	h->25	i->35	j->7	k->18	l->8	m->48	n->20	o->95	p->10	r->4	s->105	t->26	u->23	v->41	y->1	Î->1	ä->27	å->1	ö->1	
en-S	S->1	
en. 	D->5	F->1	H->2	I->1	J->3	L->1	M->2	N->1	O->2	V->2	
en."	 ->1	
en.(	E->1	I->1	
en.)	.->1	A->1	B->4	F->3	G->1	H->1	
en..	 ->9	(->3	H->1	
en.1	5->1	
en.A	l->9	n->2	r->2	t->3	v->6	
en.B	e->2	i->1	r->1	
en.C	u->1	
en.D	e->200	ä->20	å->1	
en.E	U->2	f->3	m->1	n->13	r->2	t->9	u->5	
en.F	E->1	a->2	i->1	o->1	r->6	y->1	ö->33	
en.G	e->1	o->1	å->1	
en.H	a->7	e->44	i->2	o->2	u->2	ä->6	
en.I	 ->28	n->4	
en.J	a->100	o->1	u->1	
en.K	a->5	o->19	r->1	u->1	v->1	
en.L	e->1	i->1	å->7	
en.M	a->7	e->33	i->4	o->4	y->1	ä->2	å->1	
en.N	a->2	i->6	u->4	y->1	ä->7	
en.O	c->10	m->12	r->5	z->1	
en.P	a->4	e->1	l->1	r->3	å->9	
en.R	e->2	i->1	o->1	ä->1	å->4	
en.S	a->5	e->2	i->2	k->1	l->8	n->1	o->8	t->3	u->1	y->2	ä->3	å->4	
en.T	a->4	h->2	i->5	o->2	r->2	v->1	y->3	
en.U	n->6	p->1	t->3	
en.V	a->8	e->1	i->76	å->2	
en.Ä	n->2	r->2	v->4	
en.Å	 ->2	
en.Ö	g->1	v->1	
en: 	"->1	D->1	E->1	H->1	J->2	K->2	R->1	T->1	d->3	f->3	i->1	j->1	m->2	v->4	
en:F	ö->1	
en; 	a->1	d->7	e->1	f->2	i->1	m->1	o->1	p->1	s->1	ä->1	
en?.	 ->1	
en?D	e->7	
en?E	f->1	
en?F	o->1	r->1	ö->2	
en?H	e->2	
en?I	 ->1	
en?J	a->2	
en?K	a->1	o->1	
en?N	ä->1	
en?V	a->1	e->1	i->6	
en?Ä	r->3	
enFr	å->3	
enHe	r->2	
enI 	d->1	
enJa	g->2	
enNä	s->5	
ena 	-->1	B->1	a->5	d->3	e->9	f->13	g->5	h->1	i->16	k->5	l->2	m->7	o->12	p->3	r->3	s->20	t->1	u->3	v->2	y->1	ä->4	ö->2	
ena,	 ->16	
ena.	 ->1	D->2	E->1	F->1	J->4	O->1	V->2	Ä->1	
ena;	 ->1	
ena?	P->1	
enad	 ->5	,->1	?->1	e->26	
enan	d->7	s->1	t->1	
enar	 ->34	,->2	.->2	:->1	e->35	i->5	n->5	s->4	å->1	
enas	 ->10	t->79	
enat	.->1	e->1	s->1	
enau	e->1	
enav	t->3	
enba	r->66	
enbe	r->3	t->5	
enbu	r->2	
ence	r->1	
end 	f->1	i->1	j->1	o->2	u->1	
end!	 ->2	
end,	 ->2	
end-	 ->1	
enda	 ->52	.->1	i->1	s->71	t->33	
endb	e->1	
ende	 ->230	"->1	,->11	.->21	:->22	;->1	f->2	k->1	l->1	m->1	n->36	r->27	s->2	t->38	v->6	
endi	e->1	
endo	m->5	
endr	a->1	
ends	 ->2	
endt	 ->6	,->1	
endé	e->1	
endö	v->1	
enef	i->5	
enel	u->1	
enem	a->1	
enen	 ->2	.->1	
ener	 ->7	-->10	N->1	a->27	e->19	g->109	ö->4	
enet	 ->2	i->1	
enez	u->1	
enfr	å->1	
enfä	r->1	
enfö	r->7	
enga	 ->1	g->18	r->55	
enge	l->10	n->10	
engu	e->2	
engä	l->1	
engö	r->3	
enha	m->1	n->1	
enhe	t->193	
enhä	l->32	
enhå	r->1	
eni 	f->1	s->1	
eni.	A->1	
enie	d->2	
enig	 ->1	a->4	h->9	
enin	d->1	g->88	
enis	t->2	
enjö	r->2	
enke	l->36	
enkl	a->18	i->1	
enko	l->1	n->1	
enkä	n->1	
enli	g->134	
enlö	s->1	
enna	 ->567	,->2	.->8	?->1	
ennd	r->1	
enne	 ->11	.->1	s->22	
enni	e->11	n->10	u->3	
enom	 ->230	,->1	.->2	a->2	b->7	d->6	e->3	f->161	g->16	l->2	r->1	s->18	t->1	
enor	m->32	
enov	e->3	
enpr	o->1	
enre	g->1	n->1	s->1	
enry	 ->1	
enrö	t->1	
ens 	2->1	B->3	E->3	I->1	V->1	X->1	a->41	b->44	c->1	d->33	e->35	f->81	g->17	h->17	i->48	j->4	k->38	l->25	m->56	n->16	o->73	p->31	r->79	s->101	t->30	u->48	v->36	y->7	ä->12	å->10	ö->13	
ens!	V->1	
ens,	 ->22	
ens-	 ->2	
ens.	D->6	F->1	I->1	J->2	M->1	O->1	S->1	
ens/	d->1	
ens:	 ->1	
ens?	E->1	J->1	
ensa	 ->2	m->207	r->1	t->4	v->1	
ensb	e->12	
ensd	e->2	o->1	u->2	
ense	 ->6	,->1	n->170	r->60	
ensf	r->5	ö->3	
ensh	i->2	ä->2	
ensi	b->1	d->4	f->3	n->4	o->26	s->2	t->1	v->12	
ensk	 ->2	a->313	e->2	i->28	o->18	r->38	t->2	u->5	
ensm	e->1	i->1	y->8	å->1	
ensn	a->2	i->7	
enso	m->2	r->1	
ensp	o->76	r->5	
ensr	a->1	e->10	ä->9	
enss	i->1	k->3	t->21	v->1	y->1	
enst	a->6	r->2	
ensu	t->2	
ensv	a->1	e->1	i->9	ä->1	
ensä	r->2	
ent 	(->1	-->3	1->2	A->1	C->1	a->59	b->5	e->6	f->37	g->5	h->11	i->24	k->12	l->1	m->10	o->28	p->4	r->2	s->41	t->15	u->6	v->4	ä->5	å->1	ö->3	
ent,	 ->28	
ent.	 ->1	D->8	E->2	F->4	H->2	I->4	J->5	L->1	M->3	N->1	O->1	P->1	S->1	V->1	
enta	 ->37	,->1	b->1	l->14	n->18	r->51	t->21	v->1	
ente	k->1	m->27	n->36	r->102	t->478	
entf	r->6	
enti	a->3	e->11	f->11	l->3	m->1	n->23	o->41	t->8	
entk	a->1	
entl	i->207	
ento	r->1	
entp	o->2	
entr	a->97	e->22	u->9	
ents	 ->6	a->1	b->1	f->1	i->1	k->7	l->28	u->2	
entt	i->1	
entu	e->21	r->1	s->3	
entv	a->1	ä->1	
enty	d->4	r->9	
entä	r->2	
enum	 ->4	.->1	
enus	d->1	
enut	v->1	
enve	t->1	
envi	s->5	
envä	g->8	
enz 	b->1	e->1	f->2	o->7	t->1	
enz)	(->1	.->1	
enz,	 ->3	
enzF	r->1	
enzb	e->1	
enÄr	a->1	
enäg	n->1	
enäm	t->1	
enät	 ->1	
enåd	a->1	
enèv	e->3	
enör	 ->1	s->2	
eogr	a->8	
eolo	g->5	
eomr	å->3	
eona	z->1	
eoni	 ->1	
eonl	a->1	
eord	r->1	
eore	t->2	
eost	r->2	
eote	 ->1	
ep a	t->1	
ep m	a->1	
epa 	a->1	d->6	m->4	n->2	p->1	v->1	
epa,	 ->1	
epad	e->8	
epar	 ->15	a->3	e->4	t->9	
epas	 ->5	.->2	
epat	 ->2	:->1	s->2	
epes	k->1	
ephe	r->3	
epni	n->1	
epok	 ->1	,->1	e->2	
epol	i->2	
epos	i->1	
epot	i->5	
epp 	a->1	i->5	o->2	p->3	s->1	
epp,	 ->1	
eppa	 ->1	
eppe	n->1	t->10	
epps	b->2	r->2	s->2	v->2	
epre	n->3	s->21	
epri	s->2	
epro	d->1	g->1	
epsi	s->1	
epsk	ä->1	
ept 	i->1	k->1	
ept.	D->1	H->1	
epta	b->37	n->7	
epte	 ->1	m->15	r->45	t->3	
epti	k->3	o->6	s->5	
epub	l->19	
er (	C->2	a->1	i->1	
er -	 ->48	
er 1	 ->1	0->1	9->29	
er 2	 ->1	0->5	7->1	
er 3	2->1	5->1	
er 4	 ->1	0->2	
er 5	 ->1	0->1	
er 6	0->1	
er 7	 ->1	3->1	
er 8	0->3	
er 9	0->2	7->1	
er A	l->2	m->2	r->1	z->1	
er B	N->1	S->1	a->2	r->1	
er C	o->2	
er D	a->1	u->1	
er E	G->2	M->2	U->3	h->1	k->1	l->1	r->2	u->23	x->1	
er F	N->2	a->1	i->1	ö->3	
er G	A->1	a->2	o->1	r->1	u->2	
er H	e->1	i->1	
er I	 ->1	-->1	I->4	s->3	t->1	
er J	a->1	o->2	ö->2	
er K	i->2	v->1	
er L	a->7	i->1	y->1	
er M	a->2	e->1	
er N	a->1	e->1	i->2	
er O	F->1	r->1	s->1	
er P	V->1	a->1	
er R	a->1	u->1	
er S	c->3	e->2	h->1	k->1	y->2	
er T	a->2	o->1	u->3	
er U	N->1	S->2	r->1	
er V	i->1	
er [	S->1	
er a	b->1	c->1	k->3	l->49	m->1	n->50	r->14	s->1	t->785	u->1	v->90	
er b	a->13	e->51	i->19	l->11	o->8	r->9	u->3	y->3	ä->3	å->1	ö->10	
er c	a->10	i->2	
er d	a->6	e->495	i->6	j->3	o->18	r->3	u->3	y->2	ä->23	å->12	ö->2	
er e	c->2	d->1	f->20	g->4	j->8	k->7	l->37	m->14	n->120	r->14	t->59	u->26	x->8	
er f	a->15	e->3	i->10	l->10	o->19	r->130	u->4	y->2	å->15	ö->307	
er g	a->3	e->35	i->3	j->1	l->2	o->8	r->18	y->3	ä->3	å->8	ö->12	
er h	a->79	e->36	i->4	j->1	o->10	u->29	y->1	ä->16	å->2	ö->5	
er i	 ->224	c->1	f->3	g->6	h->1	l->2	m->1	n->231	r->1	
er j	a->104	o->3	u->10	ä->4	
er k	a->32	e->1	l->3	n->2	o->110	r->18	u->7	v->5	ä->8	ö->1	
er l	a->8	e->10	i->15	o->2	u->2	y->2	ä->14	å->14	ö->3	
er m	a->46	e->140	i->80	o->21	u->1	y->15	ä->9	å->33	ö->9	
er n	a->8	e->5	i->26	o->2	u->10	y->4	ä->28	å->24	
er o	a->2	b->2	c->407	f->5	k->1	l->5	m->120	r->15	s->52	u->1	ö->1	
er p	a->10	e->7	l->4	o->7	r->26	u->3	å->162	
er r	a->10	e->38	i->10	o->1	u->3	ä->11	å->12	ö->7	
er s	a->38	e->17	i->90	j->11	k->53	l->6	m->2	n->3	o->394	p->10	t->53	u->1	v->4	y->11	ä->13	å->37	ö->3	
er t	.->1	a->16	i->163	j->2	o->13	r->25	u->2	v->12	y->3	ä->1	
er u	n->36	p->35	r->4	t->70	
er v	a->59	e->16	i->159	o->2	ä->14	å->22	
er y	t->1	
er Ö	s->4	
er ä	l->1	m->2	n->66	r->58	v->13	
er å	r->19	t->17	
er ö	k->3	n->1	p->5	r->1	v->24	
er! 	D->16	E->6	F->4	G->2	I->7	J->16	K->1	L->2	M->1	N->1	P->1	S->1	T->3	U->1	V->6	Ä->2	Å->1	
er!"	D->1	O->1	
er!D	e->5	
er!E	f->1	
er!J	a->3	
er!M	y->1	
er!V	i->2	
er" 	h->1	m->1	s->2	
er")	,->1	
er",	 ->1	
er".	D->1	
er) 	B->1	V->1	o->2	
er)F	r->2	
er)J	a->1	
er)K	o->1	
er)T	a->1	
er, 	"->1	M->1	T->1	a->24	b->13	d->30	e->22	f->26	g->7	h->23	i->24	j->4	k->12	l->6	m->48	n->12	o->63	p->7	r->5	s->72	t->19	u->19	v->23	ä->10	å->3	ö->1	
er-b	i->1	
er-k	o->1	
er-n	a->1	
er-p	r->11	
er-r	e->1	
er. 	(->1	D->4	E->2	F->1	H->1	J->1	M->2	S->2	T->1	V->1	Ä->1	
er.(	A->1	I->1	
er.)	 ->1	
er.-	 ->3	
er..	 ->1	(->2	H->1	V->1	
er.9	0->1	
er.A	l->3	n->1	t->3	v->4	
er.B	a->1	e->6	l->1	
er.C	S->1	
er.D	a->1	e->114	o->1	ä->7	å->1	
er.E	U->2	f->1	n->10	t->4	u->5	x->1	
er.F	r->9	å->1	ö->16	
er.G	e->3	
er.H	a->1	e->11	ä->6	
er.I	 ->17	n->5	t->1	
er.J	a->59	
er.K	a->2	i->1	o->19	v->1	
er.L	i->1	å->4	
er.M	a->1	e->17	i->3	ä->1	
er.N	a->2	u->1	ä->9	
er.O	c->4	m->9	r->2	
er.P	a->2	l->1	r->3	u->1	å->1	
er.R	e->2	å->1	
er.S	a->2	l->2	o->4	t->4	å->2	
er.T	a->3	e->1	i->11	r->1	
er.U	n->6	
er.V	a->12	i->35	å->1	
er.Ä	n->2	r->3	v->4	
er.Å	 ->2	
er: 	"->1	A->1	D->1	I->1	K->1	V->2	a->1	d->4	e->2	f->1	i->1	k->1	v->2	
er; 	a->1	d->3	e->1	o->1	v->1	
er?-	 ->1	
er?.	 ->1	
er?B	o->1	
er?D	e->1	
er?E	u->1	
er?H	e->3	
er?J	a->1	
er?K	o->1	
er?M	e->1	
er?P	å->1	
er?T	a->1	
er?V	e->1	i->1	
er?Ä	v->1	
erHe	r->1	
erJa	g->1	
erMe	d->1	
erNä	s->2	
era 	-->3	2->1	E->7	F->1	I->2	L->1	a->62	b->11	c->1	d->89	e->60	f->41	g->16	h->17	i->22	j->1	k->24	l->10	m->33	n->6	o->50	p->35	r->15	s->44	t->18	u->12	v->22	Ö->2	ä->7	å->5	ö->11	
era!	 ->1	
era"	.->1	
era,	 ->12	
era.	 ->1	B->1	D->5	E->2	F->1	H->2	I->2	J->6	L->2	M->3	P->1	V->1	
erad	 ->65	,->2	.->6	e->162	
erah	u->1	
eral	 ->5	a->25	d->18	e->3	i->12	l->9	s->2	t->4	
eran	-->1	b->8	d->55	s->12	t->3	v->18	
erar	 ->249	!->1	,->9	.->10	e->4	k->4	t->1	
eras	 ->215	,->13	.->22	
erat	 ->90	,->11	.->10	;->1	i->15	o->2	s->26	u->13	ö->2	
eray	,->1	
erb,	 ->1	
erba	l->1	r->3	y->1	
erbe	l->3	m->1	r->7	t->7	
erbi	l->1	s->6	
erbj	u->19	ö->1	
erbl	i->1	å->2	
erbr	i->1	y->3	
erbö	l->1	r->11	
erce	n->1	
erda	m->41	
erde	l->4	
erdo	 ->1	m->2	
erdr	i->14	
erds	t->3	
erdö	r->1	
ere 	a->1	k->1	
ere.	M->1	
ered	a->10	d->35	e->12	s->2	
ereg	l->3	
erel	l->16	
eren	d->12	g->2	s->246	t->5	
erer	a->19	ö->1	
eres	u->1	
eret	 ->1	,->1	t->6	
erex	t->6	
erfa	l->3	r->27	
erfe	k->7	
erfi	n->3	r->2	s->1	
erfl	y->2	ö->1	
erfo	r->27	
erfr	å->8	
erfu	n->2	
erfö	l->5	r->22	
erg 	f->1	g->1	k->1	o->1	
erga	v->2	
erge	 ->3	n->5	r->22	s->3	
ergi	 ->13	,->2	-->1	.->5	a->7	b->3	c->1	e->4	f->7	i->1	k->39	m->2	n->4	o->2	p->7	s->13	v->8	ä->1	å->1	
ergn	e->1	
ergr	i->14	u->1	ä->4	
ergä	l->1	
ergå	 ->1	n->11	r->3	t->1	
erha	n->6	
erhe	a->1	t->281	u->2	
erhu	s->2	
erhä	m->2	n->1	
erhå	l->12	
erhö	g->2	l->3	r->12	
eri 	-->1	a->1	f->2	i->1	k->1	m->2	n->1	o->5	ä->2	ö->1	
eri,	 ->7	
eri-	 ->1	
eri.	J->1	L->1	M->1	
eria	l->23	
erib	e->4	
erie	l->4	n->1	r->39	s->1	t->9	
erif	e->6	i->1	
erig	e->26	
erik	a->26	o->2	
eril	 ->1	a->1	
erim	s->8	å->1	
erin	 ->1	.->1	f->4	g->711	r->15	s->9	t->1	ä->3	
erio	d->86	
erip	o->1	
eris	e->4	k->1	
erit	e->1	
eriu	t->1	
eriö	s->8	
erk 	-->1	a->1	b->1	f->3	g->1	i->8	k->1	m->2	o->1	p->1	s->4	u->1	ä->2	
erk,	 ->3	
erk.	B->1	D->1	S->1	V->1	
erk?	R->1	
erka	 ->40	,->1	d->2	n->21	r->121	s->11	t->11	
erke	n->6	t->40	
erkl	a->6	i->205	
erkn	i->15	
erko	m->7	
erkr	a->1	ä->1	
erks	a->52	t->19	
erkt	y->8	
erku	r->1	
erkä	n->42	
erla	g->8	
erle	v->10	
erli	g->114	n->7	
erly	s->2	
erlä	g->7	m->18	n->18	t->18	
erlå	t->11	
erma	j->1	n->10	t->1	
erme	n->1	r->3	
ermi	d->9	n->1	s->1	
ermo	,->1	d->1	r->1	
ermå	l->1	
ermö	t->2	
ern 	(->1	-->1	E->2	b->1	d->1	e->1	f->6	g->1	h->3	i->3	k->3	l->2	m->1	n->1	o->9	p->1	r->1	s->6	t->2	u->1	v->2	ä->1	
ern,	 ->9	
ern.	)->1	.->1	D->4	H->1	J->2	O->1	V->1	Ö->1	
ern/	N->2	
erna	 ->948	!->2	"->1	,->168	.->192	/->1	:->3	;->4	?->8	H->1	r->2	s->146	t->94	
ernd	 ->3	
erne	a->1	r->3	t->10	
ernf	r->1	
erni	s->24	t->1	v->1	é->1	
erns	 ->13	
ernt	 ->4	.->1	u->1	
ernö	r->1	
erod	d->5	
eroe	n->69	
erog	a->1	
eroi	s->1	
erom	r->1	
eron	i->1	
erop	a->1	
eror	 ->18	,->1	d->5	
erot	t->1	
erpa	r->2	
erpo	l->1	p->1	s->2	
erpr	e->1	i->1	
err 	A->1	B->10	C->3	E->2	F->1	G->2	H->2	J->1	K->6	L->1	M->1	N->1	P->8	R->1	S->5	W->1	f->5	g->1	k->82	l->15	m->2	o->5	p->3	r->12	t->320	v->3	
erra	n->2	r->45	s->1	
erre	g->5	p->2	s->1	z->1	
erri	k->130	t->17	
erro	n->1	r->11	
errä	t->1	
errå	d->14	
erró	n->3	
errö	s->1	
ers 	a->10	b->10	e->3	f->5	i->3	j->1	k->1	l->4	n->1	o->2	p->6	r->4	s->5	t->1	u->5	v->2	å->1	ö->1	
ers,	 ->1	
ers-	b->1	
ersa	i->1	l->1	m->3	t->5	
erse	 ->2	l->3	n->2	r->1	
ersh	i->1	
ersi	e->9	f->2	k->18	o->13	
ersk	a->24	o->1	r->20	å->6	
ersl	u->1	
ersm	å->1	
erso	m->190	n->108	
ersp	e->22	
erst	 ->18	a->22	i->5	r->42	ä->40	å->14	ö->6	
ersu	n->3	
ersv	ä->7	
ersy	n->1	
ersä	t->35	
erså	t->1	
ersö	k->48	
ert 	C->1	G->1	a->1	b->8	d->1	e->1	f->5	g->2	h->1	i->6	k->4	l->1	m->1	o->6	p->4	s->10	t->1	u->5	v->2	y->1	ä->3	ö->1	
ert!	J->1	
ert,	 ->4	
ert.	J->1	
erta	 ->3	g->10	l->7	n->3	r->2	s->1	
erte	c->17	r->20	
ertg	r->3	
erth	e->1	u->1	
erti	d->67	f->6	k->3	l->1	n->1	s->3	
ertk	o->17	
erto	g->1	n->1	
ertr	a->3	e->1	ä->7	
ertu	t->1	
erty	g->38	
ertä	n->2	
erup	p->34	
erus	a->2	
erut	b->2	v->1	
erva	k->25	t->11	
erve	c->1	n->7	r->5	
ervi	c->7	n->74	s->1	
ervj	u->3	
ervr	i->1	
ervt	r->1	
ervu	n->3	
ervä	g->35	l->3	n->3	r->7	
ery,	 ->1	
eryk	t->1	
eräg	a->1	
eräk	n->4	
erän	 ->2	a->3	i->12	
erät	t->35	
erår	i->12	
eråt	 ->1	
eröm	t->1	v->1	
erör	 ->9	d->21	s->8	t->4	
erös	 ->2	a->1	t->2	
eröv	a->1	r->2	
es -	 ->2	
es 1	9->3	
es 2	 ->1	
es 3	,->1	
es A	d->1	
es D	e->3	
es G	i->1	
es S	p->1	
es V	i->1	
es W	i->1	
es a	l->1	n->7	r->2	t->9	u->1	v->27	
es b	a->1	e->5	l->1	o->1	r->1	y->1	ä->1	
es d	e->14	i->1	ä->3	å->1	ö->1	
es e	g->1	k->1	l->6	m->2	n->5	t->5	
es f	a->1	i->2	l->1	o->3	r->11	ö->24	
es g	e->2	ö->1	
es h	a->5	e->1	i->1	ä->1	å->1	ö->2	
es i	 ->37	g->1	h->1	n->15	
es j	u->2	
es k	l->4	o->7	r->1	u->2	v->1	
es l	e->4	o->1	
es m	a->3	e->5	o->2	y->1	ö->4	
es n	a->1	o->1	y->6	å->2	ö->2	
es o	b->1	c->14	f->1	m->4	r->1	
es p	h->1	o->2	r->2	å->5	
es r	e->5	i->2	o->1	y->1	ä->5	ö->2	
es s	a->1	e->1	i->1	j->1	k->1	l->2	o->9	p->2	t->4	v->1	ä->1	
es t	i->14	j->1	v->2	y->3	
es u	n->3	p->6	r->1	t->5	
es v	a->3	i->5	o->1	ä->3	
es y	t->1	
es ä	n->2	r->2	
es å	t->1	
es ö	g->1	k->1	v->5	
es".	K->1	
es, 	W->1	a->1	e->2	g->1	j->3	o->6	s->1	t->1	v->1	
es- 	o->6	
es-C	a->1	
es.)	Å->1	
es.A	n->1	
es.D	e->1	ä->1	
es.F	l->1	
es.H	u->1	
es.I	 ->1	
es.J	a->1	
es.K	o->1	
es.M	e->1	ä->1	
es.O	m->1	
es.R	e->1	å->1	
es.U	n->1	
es.V	a->1	i->1	
es; 	o->1	
esa 	b->1	d->1	e->1	f->1	i->3	m->1	o->3	p->1	t->1	ö->1	
esa,	 ->2	
esa.	J->1	
esam	m->7	
esan	 ->1	
esar	b->1	e->1	
esat	s->7	
esau	r->1	
esbe	d->1	s->1	
esdi	g->2	
ese 	i->1	
eseg	r->2	
esek	t->3	
esen	 ->1	t->48	
eser	 ->3	,->1	n->1	v->6	
eset	i->1	
esfo	r->1	
esfr	å->4	
esfö	r->1	
esge	m->1	
esgi	l->1	
esgå	 ->2	s->1	
esha	n->4	
esid	e->9	i->5	u->1	
esik	t->2	
esis	k->12	
esit	t->2	
eska	d->1	p->113	r->1	t->5	
eske	d->3	
eski	f->3	
eskr	e->3	i->48	
eskv	a->1	
esky	d->3	l->3	
eskå	l->1	
esla	g->26	
esli	v->2	
eslo	g->11	
eslu	t->241	
eslä	k->1	
eslå	 ->15	r->38	s->16	
eslö	t->3	
esma	n->2	
esmi	n->9	t->1	
esmä	n->1	r->1	s->1	
esnå	l->4	
esol	u->100	
eson	a->1	e->3	
esor	 ->1	
esp.	 ->2	
espa	r->5	
espe	g->1	k->80	r->7	
espo	,->1	l->3	n->2	s->1	
espr	å->9	
esqu	e->1	
esra	p->2	
esrö	r->1	
ess 	a->9	b->7	d->5	e->6	f->11	g->4	h->2	i->11	k->7	l->3	m->9	n->4	o->6	p->5	r->8	s->21	t->3	u->3	v->3	ä->2	å->3	ö->2	
ess"	.->1	
ess,	 ->2	
ess.	A->1	D->4	H->1	M->2	N->1	V->4	
ess?	J->1	
essa	 ->366	!->1	,->4	.->7	d->1	n->22	r->1	
essb	e->5	
esse	 ->21	,->5	.->3	?->1	n->116	r->25	t->5	
essh	ä->1	
essi	m->2	o->9	v->8	
essk	a->1	o->2	
essm	e->1	
essn	i->1	
esso	r->6	
essr	e->1	ä->2	
esst	r->1	
essu	e->1	t->61	
essv	ä->4	
est 	M->1	a->7	b->3	d->4	e->1	f->4	g->2	h->1	k->2	l->4	m->2	n->1	o->2	p->1	r->2	s->3	t->3	u->2	v->1	ä->1	
est,	 ->1	
est?	N->1	
esta	 ->27	,->2	d->2	n->3	r->1	s->1	t->5	u->1	
este	i->1	l->3	n->8	r->32	
esti	e->1	n->22	
estn	i->1	
esto	 ->2	d->1	r->3	
estr	a->3	i->6	u->1	å->1	
ests	.->1	
estu	n->7	
esty	r->1	
estä	l->16	m->159	n->6	
estå	 ->4	e->11	n->28	r->18	
estö	r->1	
esul	t->116	
esur	s->50	
esut	b->7	
esva	l->1	r->17	
esvi	k->8	s->2	
esvä	r->7	
esyn	n->1	
esys	t->1	
esät	t->6	
esök	 ->6	a->1	e->1	t->1	
esör	j->2	
et "	E->1	K->3	O->1	e->3	k->1	r->2	
et (	B->2	C->1	E->2	F->1	I->2	S->1	a->1	d->1	f->2	h->1	i->2	k->1	t->1	Ö->1	
et ,	 ->1	
et -	 ->33	
et 1	9->14	
et 2	1->1	2->1	
et A	B->1	k->1	l->3	
et B	N->1	e->1	r->1	
et C	a->1	
et D	a->1	e->1	
et E	U->1	l->1	q->8	r->1	u->4	
et F	ö->1	
et G	r->2	
et I	 ->1	t->1	
et K	o->1	u->3	
et L	e->2	
et M	i->1	o->3	
et P	o->4	
et R	I->1	a->1	
et S	E->1	a->1	j->1	t->1	v->1	
et T	V->1	u->1	
et V	a->1	e->1	o->1	
et a	b->4	c->4	k->7	l->32	m->2	n->104	r->24	t->258	v->337	
et b	a->15	e->112	i->5	l->27	o->6	r->16	u->3	y->3	ä->11	å->1	ö->25	
et c	e->3	h->1	i->5	
et d	a->15	e->48	i->7	j->1	o->7	r->6	y->2	ä->14	å->14	ö->2	
et e	f->12	g->12	k->8	l->21	m->3	n->82	r->7	t->13	u->31	v->2	x->13	
et f	.->1	a->94	e->12	i->191	j->4	l->4	o->16	r->83	u->9	ä->1	å->26	ö->506	
et g	a->8	e->37	i->5	j->4	l->14	o->21	r->13	y->1	ä->209	å->17	ö->24	
et h	a->207	e->18	i->8	j->2	o->13	u->2	y->1	ä->68	å->2	ö->15	
et i	 ->227	b->3	d->1	g->2	l->2	m->1	n->254	r->3	t->3	
et j	a->16	o->1	u->15	ä->3	
et k	a->62	e->1	l->12	n->1	o->134	r->45	u->11	v->6	y->1	ä->9	ö->1	
et l	a->16	e->5	i->27	o->2	u->1	y->3	ä->33	å->7	ö->6	
et m	a->13	e->215	i->12	o->25	u->3	y->17	ä->1	å->85	ö->31	
et n	a->10	e->2	i->8	o->11	u->35	y->23	ä->23	å->11	ö->13	
et o	a->5	b->3	c->361	e->1	f->9	g->1	k->1	l->3	m->108	n->4	p->2	r->13	s->2	t->3	ö->1	
et p	a->8	e->8	l->7	o->85	r->16	å->79	
et r	a->4	e->34	i->14	y->1	ä->23	å->22	ö->19	
et s	a->40	e->30	i->10	j->8	k->168	l->12	m->2	n->8	o->223	p->16	t->124	u->3	v->13	y->18	ä->60	å->36	ö->2	
et t	a->9	e->1	i->120	j->2	o->3	r->33	u->3	v->8	y->21	ä->6	å->1	
et u	n->21	p->41	r->4	t->46	
et v	a->94	e->27	i->198	o->13	ä->38	å->4	
et y	t->7	
et Ö	s->1	
et ä	c->1	g->3	m->1	n->27	r->787	v->13	
et å	l->4	r->6	t->20	
et ö	d->2	g->1	k->3	n->2	p->3	s->14	v->13	
et!(	P->1	
et!.	 ->1	(->1	
et!H	e->1	
et!K	u->1	
et!P	r->1	
et" 	(->1	g->1	m->1	o->1	ä->1	
et",	 ->2	
et".	E->1	J->1	
et) 	(->1	C->1	h->2	p->1	s->1	
et),	 ->3	
et).	D->1	H->2	L->1	
et)N	ä->1	
et, 	C->1	D->1	E->1	G->1	H->1	I->3	J->1	W->1	a->21	b->6	d->36	e->20	f->34	g->7	h->25	i->22	j->5	k->17	l->4	m->41	n->12	o->66	p->9	r->5	s->93	t->7	u->21	v->36	ä->12	å->1	ö->2	
et- 	o->1	
et-f	r->1	
et. 	(->1	D->8	E->1	J->1	K->1	M->1	S->1	V->2	a->1	
et.(	A->1	F->1	P->1	
et.)	A->1	B->2	R->1	
et.-	 ->1	
et..	 ->2	.->1	
et.1	9->1	
et.A	l->1	n->2	t->1	v->8	
et.B	e->2	l->1	r->1	
et.D	e->116	ä->9	å->1	
et.E	G->1	f->4	k->1	n->8	t->5	u->9	
et.F	l->2	r->12	ö->14	
et.H	a->4	e->23	i->1	u->2	ä->4	
et.I	 ->23	b->1	n->3	
et.J	a->79	u->1	
et.K	o->5	u->1	ä->1	
et.L	a->1	i->2	å->3	
et.M	a->8	e->28	i->6	
et.N	a->1	i->4	u->6	ä->5	ö->1	
et.O	c->7	m->5	r->2	
et.P	a->3	o->1	r->2	u->1	å->5	
et.R	a->1	e->2	ä->1	
et.S	k->2	l->1	o->4	t->3	å->8	
et.T	a->4	h->1	i->2	r->2	u->1	y->2	
et.U	n->1	r->1	t->1	
et.V	a->4	i->49	ä->1	å->2	
et.Ä	n->1	v->1	
et.Å	 ->1	r->1	t->1	
et.Ö	s->1	
et: 	"->1	F->1	J->1	U->1	d->2	e->1	f->1	k->1	o->1	t->1	v->1	ö->1	
et; 	D->1	a->1	d->1	f->2	u->1	
et? 	R->1	
et?.	 ->1	(->1	
et?A	t->1	
et?D	e->3	
et?H	e->1	u->2	
et?I	 ->1	
et?J	a->2	
et?K	o->1	ä->1	
et?N	i->2	ä->1	
et?O	c->1	
et?R	I->1	
et?S	k->1	
et?V	a->1	i->2	
et?Ä	r->1	
etJa	g->1	
eta 	-->1	a->11	b->2	d->3	e->10	f->25	h->2	i->9	k->3	m->17	n->1	o->8	p->11	r->4	s->2	t->4	u->1	v->7	å->6	ö->1	
eta,	 ->4	
eta.	 ->1	D->1	T->1	
eta?	V->1	
etab	l->13	
etad	e->2	
etag	 ->55	,->14	.->15	a->23	e->66	n->9	s->25	
etak	t->1	
etal	a->73	j->35	l->11	n->15	t->2	
etan	d->16	e->5	k->9	s->6	
etap	p->5	
etar	 ->22	,->1	.->1	e->9	i->3	k->1	n->5	
etas	 ->1	.->1	
etat	 ->12	s->2	
etbe	h->1	
etc.	 ->3	D->1	E->1	
etc?	A->1	
etde	r->1	
ete 	(->2	-->3	a->2	b->3	d->2	f->9	h->6	i->9	k->6	l->3	m->22	o->14	p->6	r->1	s->22	t->1	u->1	v->2	ä->1	å->1	
ete,	 ->11	
ete.	 ->1	.->1	A->1	D->5	F->1	H->1	I->1	J->3	K->1	L->3	M->2	N->1	P->1	R->2	S->1	U->1	V->2	Å->1	
ete?	H->1	I->1	S->1	
etec	k->12	
etee	n->3	
eten	 ->296	)->1	,->31	.->53	:->1	a->3	h->1	s->111	t->4	
eter	 ->236	,->31	.->39	?->1	a->11	i->4	l->1	n->121	s->4	
etes	s->12	
etet	 ->49	"->1	,->3	.->8	e->1	s->1	
etfr	å->2	
etfö	r->9	
eth 	S->1	
etik	 ->2	
etin	g->2	
etis	e->2	k->7	
etit	i->1	
etjä	n->1	
etko	n->16	
etkr	a->1	
etli	g->36	
etma	t->1	
etmä	s->1	
etna	 ->17	
etni	s->14	
etod	 ->13	e->16	
eton	a->45	i->1	
etor	i->3	
etpl	a->3	
etpo	l->1	s->10	
etra	k->23	n->1	r->1	
etro	a->12	l->1	
etru	s->1	
etry	c->3	g->1	
eträ	d->73	f->79	t->1	
ets 	"->1	-->1	B->1	L->1	a->15	b->28	c->1	d->21	e->4	f->40	g->31	h->8	i->3	k->7	l->12	m->16	n->4	o->41	p->13	r->20	s->37	t->12	u->9	v->4	y->3	ä->2	å->2	ö->2	
ets,	 ->2	
ets-	 ->5	
ets.	E->1	
etsa	k->1	m->6	n->5	r->5	s->3	v->2	
etsb	a->1	e->5	u->1	ö->5	
etsc	e->1	h->3	
etsd	o->4	
etse	n->6	
etsf	i->1	l->15	o->1	r->9	å->1	ö->4	
etsg	a->3	i->8	r->8	
etsh	a->2	
etsi	n->2	t->1	
etsk	a->2	l->2	o->3	r->8	
etsl	a->3	i->2	o->2	ä->1	ö->43	
etsm	a->13	e->2	y->8	ä->2	
etsn	i->2	o->6	ä->1	
etso	m->5	r->11	
etsp	a->4	e->2	l->9	o->6	r->76	
etsr	a->3	e->3	i->1	u->2	ä->3	å->18	
etss	a->1	i->2	k->2	p->1	t->3	y->3	
etst	a->40	i->48	ä->2	ö->2	
etsu	t->5	
etsv	a->1	e->1	i->5	
etsy	n->1	
etså	t->2	
ett 	"->1	5->1	A->1	E->15	a->128	b->87	c->4	d->47	e->80	f->125	g->40	h->35	i->54	j->8	k->48	l->40	m->113	n->34	o->75	p->89	r->41	s->206	t->55	u->49	v->47	w->1	y->5	ä->20	å->23	ö->16	
ett,	 ->7	
ett.	 ->1	.->1	D->2	F->1	H->1	J->1	M->2	Ä->1	
ett:	 ->2	
etta	 ->925	!->1	,->39	.->74	:->1	?->1	
ette	 ->1	-->1	r->18	t->1	
etti	c->1	d->1	g->3	o->2	
etto	n->4	
etts	 ->11	,->1	.->3	
ettv	i->1	
etun	g->1	
etut	s->10	
etvi	s->27	v->3	
ety 	ä->1	
ety-	p->1	
etyd	a->17	d->1	e->91	i->7	l->13	
etän	k->293	
etär	a->6	
etår	e->10	
etêt	e->2	
etöv	e->1	
euge	n->2	
eum 	v->1	
eund	r->3	
euro	 ->16	!->1	,->6	.->8	f->1	n->6	o->1	p->375	s->2	
euss	a->1	
eutb	i->1	
euti	q->1	
eutr	a->2	o->1	
euts	c->1	l->2	
eutv	e->4	
ev a	n->1	v->2	
ev d	i->1	j->1	ä->2	
ev f	a->1	r->1	ö->1	
ev i	n->3	
ev k	v->1	
ev n	y->1	
ev o	b->2	c->1	m->1	
ev s	o->1	
ev t	i->2	v->1	
ev u	n->2	
ev.F	r->1	
eva 	d->1	e->2	f->1	h->1	i->4	l->1	m->2	n->1	p->1	s->1	u->1	v->1	
eva,	 ->1	
eva?	N->1	
evak	a->3	n->3	
eval	d->6	
evan	d->3	t->9	
evar	a->22	
evat	t->2	
evde	 ->2	
eveb	r->1	
evek	a->1	
evel	 ->1	s->1	
even	e->1	t->20	
ever	 ->12	.->1	a->3	e->4	
evid	e->18	
evig	 ->1	t->2	
evil	j->48	
evis	 ->26	,->1	.->2	a->6	b->7	e->5	i->22	n->1	
evit	t->1	
evli	g->3	
evlå	d->1	
evna	d->12	
evol	u->1	
evs 	a->1	o->1	s->3	u->1	
evt 	d->1	e->2	i->1	
eväc	k->3	
evär	d->8	t->6	
evån	a->2	
ew Y	o->1	
ewie	s->1	
ewoo	d->2	
ex a	l->1	n->4	v->1	
ex e	u->1	
ex f	l->1	
ex m	i->1	å->10	
ex p	l->1	o->1	
ex t	i->1	u->1	
ex ö	v->1	
ex, 	s->1	
ex. 	E->1	F->1	N->1	U->1	a->2	d->2	e->1	i->1	k->2	m->2	n->2	o->1	p->1	u->1	v->1	
ex.J	a->1	
exa,	 ->1	
exak	t->18	
exam	e->6	i->10	
exan	d->2	
exas	 ->2	
exce	p->5	
exem	p->117	
exib	e->11	i->10	l->6	
exik	o->1	
exil	r->1	t->1	
exis	m->1	t->19	
exkl	u->3	
exmå	n->1	
expa	n->6	
expe	d->1	r->44	
expl	i->1	o->2	
expo	n->2	r->4	
ext 	a->1	f->1	i->1	k->1	l->1	o->3	s->5	
ext,	 ->5	
ext.	M->1	
exte	n->17	r->17	
exto	n->1	
extr	a->6	e->30	
exue	l->3	
exvä	r->1	
ey C	a->3	
eyer	 ->2	.->1	
eyhu	n->1	
ez G	o->1	
ez a	n->1	
ez o	c->1	
ez t	o->1	
ez, 	i->1	u->1	
ez-k	a->2	
ezue	l->1	
eäga	r->2	
eåte	r->1	
f - 	a->1	
f Hi	t->2	
f av	 ->1	
f el	l->1	
f ex	t->1	
f fö	r->5	
f ha	d->1	r->2	
f i 	f->1	
f in	n->1	t->1	
f ku	n->1	
f li	k->1	
f no	l->1	
f oc	h->3	k->1	
f om	 ->1	
f so	m->4	
f th	e->1	
f ut	a->1	
f äg	t->1	
f, h	a->1	
f, m	e->1	
f, o	c->1	
f, p	å->1	
f, s	o->1	
f- o	c->2	
f-Ma	t->2	
f.De	t->1	
f.Dä	r->1	
f.En	d->1	
f.Ja	g->1	
f.d.	 ->2	
fa a	l->2	r->1	
fa b	u->1	
fa d	e->2	
fa e	k->2	n->3	
fa f	o->1	r->1	ö->1	
fa i	n->1	
fa k	o->3	
fa m	i->1	
fa o	c->1	
fa r	e->1	
fa s	i->2	
fa u	n->1	t->1	
fa, 	o->1	å->1	
fa.M	e->1	
fabe	t->1	
fabr	i->1	
fack	f->4	
fadd	e->1	
fade	 ->7	r->1	s->2	
fael	 ->2	.->1	
fail	u->1	
fakt	a->9	i->49	o->14	u->64	
fala	 ->1	
fald	 ->3	,->5	e->5	i->2	
fall	 ->91	,->11	.->16	a->1	e->100	i->4	s->8	
fals	k->4	
fami	l->15	
fand	e->42	
fann	 ->2	s->14	
fant	 ->1	a->11	l->2	
far 	E->1	L->1	S->1	a->2	b->2	d->9	e->2	h->2	i->3	k->2	l->1	m->1	o->1	p->1	s->4	u->1	ä->1	ö->1	
far,	 ->4	
far.	 ->1	D->4	I->1	J->2	V->1	
far:	 ->1	
far?	K->1	
fara	 ->9	,->2	.->1	n->167	r->3	
fare	 ->1	n->25	
farh	å->2	
fari	t->2	
farl	i->59	
farm	a->1	
farn	a->1	
faro	r->4	
fars	o->1	
fart	 ->1	,->1	.->1	e->2	s->7	y->69	
farv	a->9	
fas 	h->1	o->1	t->1	v->1	
fas,	 ->2	
fas.	D->1	
fasc	i->11	
fase	n->4	
fasn	i->3	
faso	r->1	
fast	 ->24	.->2	a->5	i->1	k->1	l->5	n->1	s->72	ä->1	
fat 	e->1	g->1	i->1	p->1	s->1	
fat.	D->3	V->1	
fats	 ->2	
fatt	a->172	i->30	n->55	
faun	a->1	
favo	r->1	
faxa	 ->1	
fbes	t->1	
fdra	b->1	
febr	u->16	
fede	r->12	
fekt	 ->7	.->2	a->1	e->37	i->115	
fel 	a->4	o->3	s->3	u->1	
fel!	 ->1	
fel,	 ->4	
fel.	D->2	G->1	J->1	
fela	k->12	n->1	
felb	a->1	e->1	
fele	n->1	
felk	v->1	
felr	ä->1	
fels	y->1	
fem 	a->3	d->1	g->1	k->2	m->1	p->2	v->2	å->15	
fem,	 ->1	
fem:	 ->1	
femp	u->1	
femt	e->16	i->3	o->5	
femå	r->3	
fen 	D->1	S->1	d->1	g->1	i->1	l->1	m->4	o->2	u->2	v->1	ä->2	
fen,	 ->5	
fen-	S->1	
fen.	D->1	F->1	I->1	Ä->1	
feno	m->3	
fens	 ->1	i->3	
fent	l->80	
fer 	a->1	e->1	f->7	h->2	i->6	m->2	o->3	p->2	s->4	u->1	ä->1	
fer"	 ->1	
fer,	 ->10	
fer.	D->2	N->1	O->1	V->2	
fera	 ->3	.->1	
fere	n->179	r->3	
feri	e->1	n->1	
fern	a->12	
fert	.->1	a->1	
fess	i->2	o->6	
fest	a->1	
fety	-->1	
ff n	o->1	
ff o	c->2	
ff, 	p->1	
ff- 	o->2	
ffa 	a->3	b->1	d->2	e->5	f->3	i->1	k->3	m->1	o->1	r->1	s->2	u->2	
ffa,	 ->2	
ffa.	M->1	
ffad	e->9	
ffan	d->42	
ffar	 ->35	,->4	.->9	:->1	?->1	e->1	
ffas	 ->4	.->1	
ffat	 ->5	.->4	s->1	
ffbe	s->1	
ffek	t->153	
ffen	 ->1	-->1	s->4	t->80	
ffer	 ->9	,->3	e->5	t->1	
ffic	e->1	i->6	
ffla	g->1	
ffli	g->2	
ffpr	o->2	
ffra	 ->4	,->3	d->1	r->1	
ffre	n->14	
ffro	r->15	
ffrä	t->28	
ffär	e->11	s->1	
fhjä	l->1	
fi o	c->1	
fi p	å->1	
fi s	o->1	
fi, 	m->1	
fi.D	e->1	
fi.V	i->1	
fice	 ->1	r->38	
fici	e->8	
fick	 ->26	o->1	
fide	n->2	
fien	d->1	t->33	
fier	a->22	b->2	i->3	
fik 	o->1	s->2	ä->1	å->1	
fik-	 ->1	
fik.	B->1	D->1	
fika	 ->17	t->5	
fike	n->3	
fikl	e->1	
fikt	 ->7	
fil 	u->1	
fil.	D->1	L->1	
film	e->2	
filo	s->5	
fils	k->1	
filt	r->1	
fin 	i->1	s->1	
fin-	r->3	
fin.	V->1	
fina	 ->2	n->81	
fing	-->1	e->1	
fini	e->13	n->1	t->24	
finl	ä->5	
finn	a->60	e->39	s->317	
fins	k->6	
fint	l->10	
fiqu	e->1	
fira	 ->1	r->2	
fisk	 ->3	a->13	b->4	e->39	t->2	
fit-	a->5	
fjol	 ->2	,->1	.->1	
fjor	t->9	
fjär	d->11	
fkri	g->1	
flag	g->28	r->1	s->1	
flam	s->4	
flek	t->7	
fler	 ->24	,->1	a->56	s->1	t->5	å->12	
fles	t->25	
flex	i->27	
flic	k->1	
flig	a->1	h->1	
flik	t->16	
flir	t->1	
flit	 ->1	e->1	
flod	 ->2	e->2	
flor	a->1	
flot	t->4	
flut	e->1	n->13	
flyg	,->1	a->2	b->1	e->2	k->1	n->1	p->4	t->2	
flyk	t->16	
flyr	 ->1	
flyt	a->12	e->1	t->17	
fläc	k->1	
fläk	t->1	
flöd	e->3	i->1	
fman	n->1	
fobi	n->1	
fode	r->10	
fog 	f->1	
foga	 ->6	d->3	n->11	r->7	t->3	
foge	n->27	
foku	s->5	
folk	 ->11	,->1	.->8	a->1	e->20	g->2	h->9	l->1	n->43	o->6	p->10	r->3	s->5	v->2	
fon,	 ->1	
fond	 ->7	e->112	m->3	s->3	u->1	
fone	-->1	
for 	o->1	s->1	
fora	 ->1	
forc	e->1	
ford	-->1	e->5	o->65	r->18	
form	 ->49	,->8	.->7	:->1	a->93	e->129	f->2	i->1	n->26	p->15	s->1	u->18	å->1	
fors	 ->24	,->7	.->10	b->1	k->39	
fort	 ->3	b->1	f->89	g->5	l->1	s->95	
foru	m->5	
forê	t->1	
foss	i->3	
fost	e->1	
fotb	o->1	
fotf	ä->1	
fots	p->2	
fpro	c->2	
fra 	e->1	f->1	s->1	ä->1	
fra,	 ->3	
frad	e->1	
frak	t->11	
fram	 ->205	,->8	.->7	f->143	g->53	h->24	k->11	l->20	m->1	s->48	t->115	å->21	ö->2	
fran	c->2	s->36	
frar	 ->1	
fras	e->1	t->15	
fred	 ->15	,->1	.->4	e->2	l->8	s->63	
free	-->2	.->1	
frek	v->1	
fren	 ->11	,->1	s->2	
fres	t->5	
fri 	f->2	i->2	k->2	r->8	ö->1	
fri,	 ->1	
fri-	 ->8	
fria	 ->25	,->2	s->3	t->1	
frie	l->6	
frig	j->1	ö->5	
frih	a->2	e->113	
frik	a->6	t->1	
fris	l->2	t->14	
frit	t->5	
friv	i->12	
frod	a->4	
fron	t->4	
fror	 ->6	.->2	?->1	n->6	
fru 	A->2	F->1	P->1	R->3	S->3	T->1	W->1	k->42	t->13	
fru,	 ->1	
fruk	t->16	
frus	t->2	
frut	a->1	
frys	a->2	n->1	
fryt	t->2	
fräc	k->1	
främ	j->61	l->34	m->2	s->47	
frät	t->28	
fråg	a->525	e->11	n->8	o->272	
från	 ->596	,->3	.->2	g->1	k->3	t->3	v->9	
fsit	u->1	
fstr	a->1	ö->3	
fstö	d->2	
ft 2	0->1	
ft a	l->1	t->4	v->4	
ft b	e->2	
ft d	e->4	ä->1	
ft e	n->1	r->1	t->2	x->1	
ft f	a->1	l->1	r->4	ö->8	
ft g	e->1	
ft h	a->1	
ft i	 ->5	n->1	
ft k	a->1	o->1	
ft l	a->1	
ft m	e->3	y->1	å->1	ö->1	
ft n	ä->2	å->2	
ft o	c->4	m->2	
ft p	r->2	å->3	
ft r	e->1	
ft s	a->1	e->1	i->1	k->3	o->6	t->3	v->1	å->2	
ft t	a->1	i->4	
ft u	n->1	t->1	
ft v	i->2	ä->1	å->1	
ft ä	r->4	
ft!H	e->1	
ft, 	S->1	f->1	i->1	m->3	o->2	s->2	u->1	v->2	
ft. 	D->1	
ft.A	t->1	
ft.D	e->2	ä->1	
ft.E	f->1	
ft.H	e->1	
ft.J	a->1	
ft.M	e->1	
ft.O	m->1	
ft.V	i->4	
ft: 	d->1	
ft? 	M->1	
ft?N	e->1	
fta 	a->8	b->5	d->3	e->1	f->8	g->2	h->7	i->3	k->1	l->2	m->1	n->2	o->5	p->2	s->8	t->2	u->3	v->2	ä->5	
fta,	 ->1	
fta.	O->1	
ftad	e->6	
ftan	 ->2	d->5	
ftar	 ->37	e->3	l->2	n->2	
ftas	 ->7	.->1	t->1	
ftat	 ->6	s->2	
ftbu	r->1	
fte 	a->9	d->1	g->1	i->1	m->1	o->1	s->2	u->1	v->1	ä->2	
fte,	 ->1	
fte.	D->1	V->1	
ftel	s->1	
ften	 ->32	,->2	.->7	a->1	
fter	 ->203	,->9	.->9	:->1	;->1	b->1	f->11	g->8	h->5	l->6	m->9	n->21	s->205	t->6	å->1	
ftet	 ->25	.->1	
ftfu	l->12	
ftig	 ->12	,->1	a->20	t->16	
ftli	g->8	
ftni	n->113	
ftom	r->1	
fton	e->1	
ftor	,->1	n->2	
fts-	 ->1	
ftsa	n->4	
ftsf	ö->2	
ftsl	ä->2	
ftsm	å->1	
ftso	l->1	
ftsp	l->1	o->1	r->2	
ftsr	e->1	
ftss	e->1	ä->1	
ftst	a->1	
ftsv	e->1	
ftsä	k->1	
ftta	g->1	
fttr	ä->4	
ftve	r->8	
full	 ->15	.->3	a->24	b->3	f->3	g->2	h->1	k->5	o->5	s->41	t->43	v->2	ä->2	
fult	 ->1	
fund	a->1	e->17	
fung	e->54	
funk	t->32	
funn	a->2	e->1	i->9	
fuse	"->1	
fusi	o->8	
fusk	.->1	
futt	i->1	
fyll	a->35	d->1	e->19	s->3	t->4	
fyra	 ->23	,->1	:->1	
fyrt	i->3	
fysi	s->9	
fäde	r->1	
fäkt	a->1	
fälh	a->1	
fäll	d->2	e->92	i->18	t->2	
fält	 ->1	e->5	
fäng	d->1	e->1	
fär 	1->3	7->1	l->1	s->2	t->2	
fära	n->1	
färd	 ->2	,->2	;->1	a->12	i->13	s->6	
färe	n->4	r->8	
färg	,->2	a->1	
färl	i->2	
färr	e->2	
färs	k->1	m->1	
fäst	 ->3	a->8	e->12	n->1	s->1	
få 1	0->1	
få E	u->1	
få G	o->1	
få a	l->1	n->1	r->1	v->2	
få b	e->3	o->2	ä->2	ö->1	
få d	e->14	i->1	o->1	
få e	f->2	n->27	r->1	t->11	
få f	a->1	i->1	l->1	o->1	r->4	u->1	ö->4	
få g	a->1	e->1	
få h	i->1	j->1	
få i	 ->3	g->1	n->3	
få k	o->4	v->2	
få l	a->1	i->1	o->2	ä->3	
få m	a->2	e->2	y->1	å->3	ö->1	
få n	å->3	
få o	b->1	m->1	r->2	s->2	
få p	a->1	e->2	o->2	r->2	u->1	å->1	
få r	e->3	y->1	ä->1	
få s	a->2	e->6	i->2	l->1	t->9	ä->2	å->3	
få t	a->6	i->16	
få u	p->1	t->2	
få v	a->1	e->6	i->3	å->1	
få ä	r->1	
få å	t->1	
få ö	k->1	
få, 	o->2	r->1	
få.E	u->1	
få.G	r->1	
få.V	i->1	
fåge	l->3	
fågl	a->6	
fång	 ->1	a->4	e->1	s->8	
får 	M->1	O->1	a->7	b->3	d->14	e->19	f->6	g->5	h->3	i->39	j->2	k->5	l->2	m->10	n->4	o->5	p->2	r->1	s->15	t->11	u->2	v->21	y->1	ä->2	å->1	
får,	 ->2	
får?	N->1	
fårk	ö->1	
fås 	f->1	
fåta	l->1	
fått	 ->56	.->1	
fére	n->1	
född	.->1	e->1	
föde	l->2	r->2	
födn	i->1	
födo	ä->1	
föds	 ->1	
föga	 ->2	
följ	a->80	d->43	e->17	n->10	s->4	t->4	
föll	 ->6	.->1	
föns	t->1	
för 	"->4	-->4	1->15	2->7	3->1	5->2	7->2	A->4	B->6	C->2	D->3	E->70	F->5	G->2	H->1	I->4	K->7	L->2	O->1	P->3	S->3	T->8	V->1	W->2	a->935	b->83	c->7	d->538	e->240	f->123	g->42	h->84	i->60	j->30	k->161	l->59	m->167	n->76	o->99	p->73	r->109	s->206	t->90	u->101	v->125	y->3	Ö->2	ä->31	å->34	ö->46	
för"	.->1	
för,	 ->27	
för.	 ->1	(->1	.->1	D->4	H->1	J->1	M->3	V->5	
för:	 ->3	
för;	 ->1	
för?	D->1	F->2	I->1	Ä->1	
föra	 ->151	,->1	.->3	k->1	l->1	n->311	r->2	s->42	
förb	a->14	e->33	i->32	j->14	l->15	r->5	u->33	ä->78	
förd	 ->1	,->1	a->5	e->66	j->11	o->2	r->163	u->3	ä->4	ö->20	
före	 ->26	b->25	d->160	f->21	g->19	h->1	k->22	l->29	m->13	n->38	s->164	t->271	
förf	a->83	i->1	j->1	l->18	o->18	r->5	ä->3	å->1	ö->5	
förg	l->2	r->3	ä->1	
förh	a->95	i->30	o->9	å->56	ö->1	
föri	n->15	r->1	
förk	a->9	l->76	n->3	o->2	r->1	u->2	
förl	a->3	e->2	i->79	o->20	u->9	ä->6	å->4	
förm	e->5	i->3	o->11	y->1	å->48	ö->1	
förn	a->1	e->10	u->14	y->49	
föro	l->2	r->77	
förp	a->5	l->21	
förr	 ->3	,->1	a->42	e->4	g->3	i->1	ä->5	å->1	
förs	 ->22	,->2	.->6	a->12	e->31	i->66	k->10	l->484	o->5	t->397	u->9	v->83	ä->59	å->1	ö->64	
fört	 ->28	,->2	.->1	e->3	i->6	j->20	r->65	s->29	v->1	y->3	ä->1	
föru	n->1	t->77	
förv	a->55	e->22	i->19	r->1	ä->53	å->6	
förä	n->73	
förå	l->3	
förö	d->5	v->3	
fött	e->3	
g (1	9->1	
g (E	G->1	
g (a	r->2	
g (r	e->1	
g (å	t->1	
g - 	S->1	a->1	d->5	g->1	i->1	j->1	m->2	o->7	s->2	t->1	ä->1	
g -,	 ->2	
g 1 	m->1	o->1	
g 1,	 ->1	2->1	
g 10	 ->4	.->1	
g 11	,->1	
g 12	 ->1	
g 13	 ->1	
g 15	 ->1	
g 17	 ->1	,->1	
g 18	 ->2	
g 19	 ->2	9->3	
g 2,	 ->2	
g 20	 ->1	0->1	
g 22	 ->1	,->2	
g 23	 ->1	
g 26	 ->1	
g 3 	o->1	
g 34	 ->1	
g 37	/->1	
g 38	 ->2	:->1	
g 4 	o->1	
g 4.	I->2	
g 43	 ->1	
g 44	 ->1	
g 45	.->3	
g 5,	 ->2	
g 6 	o->2	
g 60	0->1	
g 68	5->1	
g 80	 ->2	
g De	t->1	
g Ec	e->1	
g Eu	r->2	
g Fä	s->1	
g Ga	z->1	
g Ha	i->14	
g IN	T->1	
g IV	 ->2	
g Ir	l->1	
g OL	A->1	
g Ta	d->1	
g VI	 ->1	
g [K	O->1	
g ab	s->1	
g ac	c->3	
g aj	o->1	
g ak	t->1	
g al	d->2	l->10	
g an	 ->2	d->1	g->1	l->2	m->1	n->5	s->91	t->7	v->3	
g ar	a->1	b->5	t->1	
g as	s->2	
g at	t->203	
g av	 ->355	e->1	g->1	l->1	r->2	s->7	t->1	v->3	
g ba	d->2	k->4	r->14	s->2	
g be	 ->3	a->2	f->6	g->6	h->4	k->15	r->25	s->8	t->11	u->1	v->2	
g bi	d->1	l->2	
g bl	a->2	e->5	i->6	
g bo	r->5	
g br	a->2	o->2	
g by	r->3	
g bä	r->2	
g bö	r->10	
g ci	t->2	
g da	g->1	
g de	 ->8	b->8	l->18	m->3	n->14	s->3	t->19	
g di	a->2	r->1	s->3	
g dj	u->1	
g do	c->5	
g dr	a->2	o->1	
g dy	l->1	
g dä	r->17	
g då	 ->1	
g dö	d->1	r->2	
g e.	d->1	
g ef	f->2	t->6	
g ek	o->1	
g el	l->22	
g em	e->4	o->6	
g en	 ->28	b->1	d->3	h->1	s->1	
g er	 ->8	,->2	h->1	i->2	k->2	
g et	t->20	
g eu	r->1	
g ev	e->1	
g ex	 ->1	a->1	i->1	p->1	
g fa	k->1	r->1	s->2	
g fe	l->1	
g fi	c->3	e->1	n->8	
g fo	r->7	
g fr	a->28	e->4	i->1	ä->1	å->84	
g fu	l->2	n->5	
g fä	l->1	
g få	r->13	t->3	
g fö	l->1	r->296	
g ga	n->1	r->3	v->1	
g ge	 ->4	n->13	r->5	
g gi	c->1	v->2	
g gj	o->5	
g gl	a->2	o->1	ä->9	
g go	d->1	
g gr	a->17	o->1	u->9	
g gä	l->4	r->8	
g gå	r->2	
g gö	r->4	
g ha	 ->4	d->5	n->8	r->138	
g he	d->1	l->11	m->1	n->1	
g hi	e->1	n->1	s->1	t->1	
g hj	ä->3	
g ho	p->54	s->3	t->1	
g hu	r->3	v->1	
g hä	l->2	n->8	r->10	v->5	
g hå	l->15	
g hö	j->1	l->1	r->6	
g i 	"->1	B->2	D->1	E->15	F->1	I->1	K->3	M->1	S->3	T->2	Y->1	a->5	b->4	d->45	e->23	f->24	g->1	h->4	j->2	k->7	m->11	o->2	p->3	r->8	s->22	t->2	u->5	v->9	Ö->2	
g i,	 ->1	
g i.	S->1	
g ia	k->1	
g ih	o->1	
g in	 ->9	d->1	f->16	g->7	k->2	n->9	o->18	r->3	s->18	t->79	v->1	
g ir	r->1	
g iv	ä->1	
g ja	g->2	
g jo	n->1	
g ju	 ->2	r->1	s->2	
g jä	m->3	
g ka	m->1	n->74	p->1	r->2	t->2	
g kl	.->2	a->3	
g kn	a->2	
g ko	l->1	m->64	n->15	p->1	r->1	s->3	
g kr	a->1	i->2	ä->2	
g ku	l->2	n->6	
g kv	a->2	
g kä	n->10	r->1	
g kö	p->1	
g la	d->1	g->9	n->1	r->1	
g le	d->5	g->2	
g li	d->1	g->1	k->2	s->1	t->4	
g ly	f->2	s->5	
g lä	g->4	m->2	n->3	r->1	s->3	x->1	
g lå	n->1	t->2	
g lö	s->6	
g ma	j->1	k->3	n->11	r->2	x->1	
g me	d->76	l->15	n->14	r->11	s->1	
g mi	g->16	l->2	n->8	s->2	
g mo	t->27	
g my	c->13	n->1	
g mä	r->3	
g må	h->1	l->1	n->5	s->34	
g mö	j->2	
g na	i->1	t->6	
g ne	d->3	g->1	
g ni	 ->7	v->7	
g no	g->3	l->1	t->4	
g nr	 ->2	
g nu	 ->7	m->1	
g ny	n->1	s->1	t->1	
g nä	m->7	r->16	s->3	
g nå	g->2	
g nö	d->3	
g ob	e->3	
g oc	h->235	k->29	
g oe	r->1	
g of	 ->1	f->2	t->2	
g ol	j->1	
g om	 ->105	.->1	b->2	e->1	f->1	p->1	s->1	ö->1	
g on	d->1	ö->1	
g or	d->2	i->1	o->1	
g os	v->1	
g pa	r->2	
g pe	k->1	r->10	
g pl	a->1	ä->1	
g po	l->8	s->3	ä->2	
g pr	a->1	e->2	i->1	o->8	
g pu	n->7	
g på	 ->99	,->2	.->2	b->1	g->1	m->5	p->2	s->1	v->3	
g ra	d->1	m->2	p->1	t->1	
g re	a->3	d->15	f->5	g->5	k->4	l->1	s->7	v->1	
g ri	k->4	s->3	
g ro	l->8	
g ru	m->1	
g ry	k->1	
g rä	d->1	k->7	t->3	
g rå	d->5	
g rö	r->4	s->11	
g sa	d->11	g->1	k->2	m->9	t->1	
g se	 ->1	d->3	g->1	i->1	k->3	m->1	n->1	r->13	t->1	
g si	g->5	k->9	m->1	n->3	t->5	
g sj	ä->25	
g sk	a->54	e->1	i->2	r->1	u->124	y->3	ä->1	
g sl	u->2	
g so	c->2	l->2	m->229	
g sp	e->1	r->1	
g st	a->5	o->2	r->7	ä->9	å->5	ö->13	
g su	b->1	
g sv	a->3	
g sy	f->4	m->2	n->1	s->3	
g sä	g->38	k->5	n->1	r->5	t->1	
g så	 ->4	d->1	g->2	l->2	v->2	
g t.	e->1	
g ta	 ->5	c->29	g->4	l->15	n->1	r->6	s->1	
g te	k->2	r->1	
g ti	d->22	l->200	
g to	g->2	l->1	
g tr	a->1	o->117	ä->2	
g tv	e->1	i->3	u->1	å->1	
g ty	c->42	d->5	v->2	
g tä	n->16	v->1	
g un	d->27	
g up	p->57	
g ur	v->1	
g ut	 ->6	a->15	b->4	e->2	f->3	g->7	k->1	m->2	o->1	s->7	t->11	v->2	ö->1	
g va	d->11	k->1	l->1	r->26	
g ve	r->11	t->24	
g vi	 ->11	d->10	l->268	s->6	
g vo	r->1	
g vä	d->2	g->4	l->18	n->7	r->1	x->1	
g vå	g->2	
g yr	k->1	
g yt	t->1	
g Ös	t->2	
g äg	n->2	
g äl	s->1	
g än	 ->3	d->10	n->1	
g är	 ->160	,->2	l->1	o->1	
g äv	e->6	
g å 	P->1	e->1	u->1	
g åk	l->1	
g ås	i->3	t->1	
g åt	 ->21	,->1	e->3	g->5	s->1	
g ök	a->2	n->1	
g ön	s->6	
g öp	p->1	
g öv	e->17	n->1	
g!".	D->1	
g!Ha	n->1	
g!Ja	g->1	
g" a	v->1	
g" o	c->1	
g" s	o->1	
g", 	m->1	o->1	
g".E	u->1	
g".J	a->1	
g".N	ä->1	
g) i	 ->1	n->1	
g) o	c->2	
g), 	t->1	
g).V	i->1	
g)Nä	s->1	
g, B	r->1	
g, I	l->1	
g, O	L->1	
g, a	c->1	n->1	t->9	v->3	
g, b	e->1	l->4	å->2	ö->1	
g, d	e->15	r->1	v->5	ä->3	
g, e	f->15	l->3	n->10	t->5	
g, f	a->3	i->1	o->2	r->8	ö->26	
g, g	e->3	r->2	u->1	ö->1	
g, h	a->5	e->8	å->1	
g, i	 ->11	n->10	r->1	
g, j	u->1	ä->6	
g, k	a->1	l->1	o->3	r->1	u->1	
g, l	e->3	i->3	å->2	
g, m	a->1	e->25	i->5	o->2	å->1	
g, n	u->2	y->1	ä->11	å->1	
g, o	a->1	c->36	m->2	t->1	
g, p	e->1	r->2	å->6	
g, r	ä->1	å->1	
g, s	a->3	j->1	k->4	n->1	o->28	p->3	t->2	ä->4	å->13	
g, t	a->3	i->2	j->1	o->1	r->2	v->1	ä->1	
g, u	p->1	t->16	
g, v	a->5	i->22	o->1	
g, ä	r->6	v->4	
g, å	t->3	
g, ö	v->1	
g-PM	 ->1	
g. D	e->3	
g. E	n->1	
g. F	ö->1	
g. H	ä->1	
g. M	e->1	
g. P	å->1	
g. S	k->1	å->1	
g.(A	p->2	
g.)F	ö->2	
g.)H	e->1	
g.. 	(->2	F->1	
g..(	D->1	
g.Al	l->4	
g.An	d->1	s->1	
g.Ar	b->1	
g.Av	 ->5	s->1	
g.Be	k->1	t->1	
g.Bi	l->1	
g.Br	i->1	
g.Da	l->1	n->1	
g.De	 ->8	n->23	s->2	t->67	
g.Di	s->1	
g.Do	k->1	m->1	
g.Dä	r->10	
g.Ef	f->1	t->3	
g.Em	e->1	
g.En	 ->2	d->1	l->4	
g.Er	i->2	
g.Et	t->1	
g.Eu	r->3	
g.Fl	e->1	
g.Fr	a->1	u->4	å->4	
g.Fö	r->19	
g.Ge	n->4	
g.Gr	u->1	
g.Ha	n->2	
g.He	r->20	
g.Hu	r->2	
g.Hy	c->1	
g.Hä	r->1	
g.Hö	g->1	
g.I 	d->13	e->1	f->1	n->1	s->2	v->2	
g.In	g->2	t->1	
g.Ja	g->62	
g.Ju	s->1	
g.Ka	n->1	t->1	
g.Ko	m->9	n->2	r->1	s->1	
g.Le	d->1	
g.Li	k->1	v->1	
g.Lå	t->3	
g.Ma	l->1	n->7	r->1	
g.Me	d->2	n->7	
g.Mi	n->1	
g.My	n->1	
g.Må	h->1	l->1	n->2	
g.Mö	j->1	
g.Na	t->2	
g.Ni	 ->3	
g.Nu	 ->3	
g.Nä	r->3	
g.Nå	j->1	
g.Oa	v->1	
g.Oc	h->11	
g.Of	t->1	
g.Om	 ->10	
g.PP	E->1	
g.Pa	r->2	
g.Pr	o->2	
g.På	 ->2	
g.Ra	p->1	
g.Re	f->1	t->1	
g.Sa	m->3	
g.Se	d->1	
g.Sk	a->1	u->1	
g.Sl	u->4	
g.Sy	f->1	
g.Så	 ->1	
g.Ta	c->2	
g.Ti	l->3	t->1	
g.Tr	o->1	
g.Un	d->1	g->1	
g.Va	d->4	r->2	
g.Vi	 ->26	l->1	s->2	
g.Vå	r->2	
g.a.	 ->1	
g.Är	 ->3	a->1	
g: D	e->1	
g: d	e->2	i->1	
g: e	t->1	
g: f	ö->1	
g: h	a->1	
g: i	n->1	
g: j	a->1	
g:De	n->1	t->1	
g; d	e->2	
g; e	n->1	
g; f	ö->3	
g; m	i->1	
g; s	l->1	
g?De	n->2	t->2	
g?Dä	r->1	
g?Fi	n->1	
g?Fr	u->1	
g?Fö	r->1	
g?Hu	r->1	
g?Hä	r->1	
g?Ja	g->1	
g?Jo	,->1	
g?Ol	i->1	
g?Ty	c->1	
g?Va	d->1	
g?Är	 ->1	
gNäs	t->1	
ga "	A->1	i->1	
ga -	 ->8	
ga 2	 ->1	
ga 3	7->1	
ga B	e->2	o->1	
ga E	U->2	l->1	u->4	v->1	
ga F	i->1	l->3	r->3	
ga H	a->2	u->1	
ga I	z->1	
ga J	a->1	e->1	o->1	
ga K	o->1	
ga L	i->1	
ga M	u->1	
ga N	a->1	i->1	
ga R	a->1	o->1	
ga S	a->2	v->1	
ga a	d->2	g->2	k->1	l->3	n->19	p->2	r->9	t->121	v->30	
ga b	a->2	e->42	i->12	l->2	o->2	r->8	u->5	ä->1	å->1	
ga c	e->1	h->1	
ga d	a->3	e->46	i->7	o->4	ä->1	å->3	
ga e	f->6	g->1	k->1	l->5	n->11	r->4	t->7	u->2	x->2	
ga f	a->10	e->2	i->4	l->4	o->7	r->108	å->2	ö->91	
ga g	a->3	e->10	i->3	n->1	o->2	r->16	ä->3	å->3	
ga h	a->12	e->3	i->2	o->1	u->6	y->1	ä->6	ö->2	
ga i	 ->28	.->1	a->1	c->1	d->2	f->1	g->1	m->1	n->31	r->1	
ga j	a->2	u->1	
ga k	a->5	e->1	l->2	o->49	r->7	v->4	ä->1	
ga l	a->3	e->2	i->12	o->1	ä->9	ö->4	
ga m	a->4	e->45	i->10	o->6	u->1	y->2	ä->5	å->9	ö->2	
ga n	a->3	e->4	i->3	o->1	r->24	y->6	ä->8	å->10	
ga o	b->1	c->76	e->1	f->2	k->1	l->5	m->94	r->15	s->6	
ga p	a->5	e->2	l->2	o->6	r->19	u->3	å->11	
ga r	a->6	e->38	i->3	o->1	u->18	ä->40	å->9	ö->1	
ga s	a->10	c->1	e->8	i->16	k->15	l->1	m->1	o->52	p->4	t->67	u->2	v->8	y->6	ä->5	å->3	
ga t	a->8	e->7	i->28	j->5	o->2	r->5	u->3	y->2	
ga u	n->5	p->19	t->20	
ga v	a->10	e->7	i->17	r->2	ä->10	å->3	
ga y	t->2	
ga ä	m->13	n->13	r->15	v->1	
ga å	k->1	r->9	s->1	t->15	
ga ö	a->1	n->1	p->2	s->1	v->9	
ga! 	V->1	
ga!D	e->1	
ga!F	r->1	ö->1	
ga!J	a->1	
ga!Ä	v->1	
ga, 	E->1	a->7	b->1	d->4	e->7	f->9	h->5	i->5	k->6	l->2	m->3	n->3	o->16	p->4	r->1	s->5	u->2	v->8	ä->1	å->1	
ga. 	M->2	
ga.(	T->1	
ga.-	 ->1	
ga.A	l->1	n->1	v->2	
ga.D	e->12	ä->1	
ga.E	n->2	t->1	
ga.F	r->1	ö->5	
ga.H	e->5	
ga.I	 ->5	n->1	
ga.J	a->14	
ga.M	a->1	e->5	
ga.N	i->3	
ga.O	c->1	m->2	
ga.P	å->2	
ga.S	o->1	å->1	
ga.T	i->1	
ga.U	t->1	
ga.V	i->12	
ga.Ä	v->1	
ga/h	a->1	
ga: 	"->1	D->1	F->1	N->1	d->1	h->2	o->1	v->3	
ga; 	v->1	
ga?.	 ->1	
ga?D	e->1	
ga?F	ö->1	
gad 	d->1	m->2	o->15	p->1	r->1	s->1	
gad,	 ->1	
gad.	D->1	K->1	M->1	V->1	
gade	 ->31	,->1	.->1	s->7	
gado	,->1	
gage	m->9	r->9	
gagn	 ->3	a->8	
gagå	n->6	
gakt	u->1	
gal 	K->1	b->1	i->1	k->1	o->9	p->3	s->1	t->1	ä->1	
gal,	 ->4	
gala	 ->7	
gale	n->1	
gali	s->1	t->1	
gall	r->1	
galn	a->1	
gals	 ->7	
galt	 ->9	
galu	n->3	
gam 	g->1	
gam,	 ->1	
gaml	a->28	
gamm	a->4	
gan 	-->2	1->1	B->2	D->1	J->1	K->2	L->1	N->1	P->1	S->1	W->3	a->6	c->1	d->3	f->11	g->6	h->2	i->14	j->1	k->3	m->2	n->3	o->104	p->2	r->1	s->15	t->2	u->2	v->5	y->1	ä->16	å->1	
gan"	,->1	
gan,	 ->20	
gan.	D->1	E->1	F->3	H->2	I->1	J->4	K->2	S->2	U->1	V->1	
gan:	 ->5	
gan;	 ->1	
gan?	J->1	
gand	a->3	e->385	
gane	n->5	t->4	
gani	 ->1	,->4	s->61	
gans	 ->1	k->26	v->3	
gant	 ->1	i->5	
gapr	o->1	
gar 	(->3	-->3	E->2	R->1	a->45	b->5	d->12	e->10	f->34	g->5	h->11	i->34	j->6	k->6	m->21	n->4	o->74	p->15	r->1	s->62	t->19	u->5	v->15	ä->16	å->2	ö->7	
gar!	M->1	
gar"	 ->1	
gar)	.->1	
gar,	 ->64	
gar-	 ->1	
gar.	 ->2	)->1	-->1	.->1	B->2	D->20	E->4	F->8	H->4	I->6	J->12	K->3	L->3	M->1	N->1	O->6	P->1	R->2	T->4	U->1	V->12	Ä->1	
gar:	 ->7	
gar;	 ->1	
gar?	J->1	
gara	n->96	
gard	e->2	
gare	 ->241	!->1	"->1	,->27	.->23	:->1	?->1	l->1	n->31	s->10	
gari	e->1	k->15	n->1	
garl	a->2	ä->1	
garm	y->14	
garn	a->286	
gars	 ->5	k->7	
garv	ä->1	
garä	m->1	
gas 	a->5	b->1	d->2	e->4	f->5	i->3	k->2	m->1	p->4	r->1	s->1	t->3	u->4	v->3	ä->1	ö->1	
gas,	 ->8	
gas.	D->1	E->2	J->1	N->1	P->1	R->1	V->3	
gasa	t->1	
gase	r->5	
gask	a->2	
gast	 ->1	,->1	e->54	
gasä	t->19	
gat 	E->2	a->4	e->3	f->4	l->1	m->2	n->1	o->1	r->1	s->4	t->1	
gat,	 ->3	
gat.	D->1	V->1	
gata	 ->1	
gate	l->2	
gati	o->16	v->27	
gato	r->15	
gats	 ->6	.->1	
gau 	f->3	o->1	s->3	
gau,	 ->5	
gau.	E->1	
gauM	e->1	
gaub	e->1	
gaus	 ->3	
gav 	K->1	e->1	h->3	i->1	m->2	n->1	o->1	p->1	s->1	u->1	v->1	
gav,	 ->1	
gava	r->1	
gavs	 ->5	
gbar	 ->2	.->1	a->2	t->10	
gber	o->1	
gbla	d->1	
gbox	n->1	
gbro	 ->1	
gbyg	g->1	
gd a	t->1	v->1	
gd b	a->1	r->1	
gd f	o->1	r->2	ö->2	
gd g	e->1	
gd i	 ->2	n->2	
gd l	ö->1	
gd n	i->1	
gd o	c->3	l->1	m->1	t->1	
gd p	å->2	
gd s	a->1	o->1	
gd y	t->1	
gd ä	n->1	
gd å	t->1	
gd, 	m->1	
gd.D	e->2	
gda 	a->1	f->1	h->2	o->1	r->1	t->1	ä->1	
gda.	V->1	
gde 	"->1	p->1	s->1	v->1	
gden	 ->18	,->3	.->7	s->8	
gder	 ->5	
gdes	 ->1	
gdom	 ->4	,->2	.->1	/->1	a->7	e->4	s->8	
gdpu	n->4	
gdra	g->2	
gdsb	e->1	
gdsk	o->1	
gdso	m->4	
gdsr	e->2	
gdst	u->1	
gdsu	t->1	
gdyr	k->1	
ge E	u->1	
ge F	r->1	u->1	
ge a	k->2	l->3	n->4	r->2	t->4	
ge b	e->1	i->3	u->1	ä->1	å->1	
ge d	e->17	ä->1	å->1	
ge e	n->13	r->7	t->12	
ge f	e->1	ö->3	
ge g	a->1	e->1	r->1	
ge h	a->3	j->2	ö->1	
ge i	 ->2	n->4	
ge j	o->1	
ge k	l->2	o->4	u->1	
ge m	a->2	e->3	i->2	
ge n	u->1	ä->1	å->2	
ge o	c->8	f->1	m->1	r->1	s->8	
ge p	a->3	e->2	i->1	o->1	r->2	å->3	
ge r	a->1	e->3	i->1	o->1	ä->1	å->3	
ge s	e->5	i->4	n->1	o->10	t->2	ä->1	å->2	
ge t	i->2	r->1	y->1	
ge u	n->2	p->2	t->9	
ge v	a->3	e->1	i->3	ä->2	å->1	
ge ä	n->1	r->1	
ge å	t->1	
ge, 	b->1	d->1	m->1	s->1	
ge. 	D->1	
ge.H	e->1	
ge.J	a->2	
ge.O	m->1	
ge.V	å->1	
ge?H	e->1	
gedi	 ->1	.->1	e->2	g->2	
gefä	r->10	
geko	m->1	
gel 	r->1	s->1	ä->2	
gel,	 ->1	
gelb	r->1	u->15	
geli	l->1	
gell	i->1	ö->1	
gelm	e->1	ä->2	
geln	 ->6	s->2	
gelr	ä->2	
gels	e->19	k->10	m->1	y->2	
gelv	e->19	ä->1	
gelä	g->22	n->1	
gema	n->13	
geme	n->386	
gen 	-->7	1->9	2->3	3->4	4->2	7->1	A->2	B->2	E->2	F->1	J->1	K->1	W->1	a->292	b->52	d->25	e->39	f->107	g->35	h->69	i->124	j->3	k->67	l->10	m->73	n->12	o->99	p->44	r->23	s->107	t->75	u->24	v->50	ä->48	å->5	ö->7	
gen!	R->1	
gen"	 ->1	,->2	
gen,	 ->130	
gen.	 ->5	(->1	.->1	A->3	B->1	C->1	D->35	E->4	F->6	G->1	H->12	I->4	J->16	K->4	L->2	M->9	N->1	O->1	P->2	R->1	S->5	T->4	U->2	V->12	Ä->1	
gen:	 ->9	
gen;	 ->3	
gen?	D->4	F->1	H->1	V->1	
genI	 ->1	
gena	 ->1	,->1	n->2	r->3	s->10	v->3	
genb	e->1	
gend	a->1	e->7	o->5	
gene	r->38	t->1	
genf	ö->5	
geng	ä->1	
genh	e->39	
genj	ö->2	
genk	o->1	ä->1	
geno	m->419	
genr	e->1	
gens	 ->88	,->2	e->3	k->24	t->1	v->1	
gent	 ->4	.->1	a->1	e->27	i->22	l->43	u->1	
genu	s->1	
genä	m->1	
geog	r->8	
geos	t->2	
ger 	-->1	1->1	2->1	5->1	E->3	S->1	a->44	b->11	d->23	e->24	f->34	g->4	h->10	i->42	j->12	k->9	l->5	m->20	n->12	o->20	p->15	r->7	s->32	t->22	u->17	v->17	ä->3	ö->1	
ger!	 ->58	D->3	E->1	J->2	V->1	
ger,	 ->30	
ger.	 ->1	A->1	D->2	E->1	F->1	H->2	J->2	N->1	O->2	P->1	T->2	
ger:	 ->6	
ger;	 ->1	
gerM	e->1	
gera	 ->53	!->1	,->5	.->7	d->5	n->18	r->30	s->1	t->10	
gerb	e->1	
gere	x->6	
geri	 ->5	,->5	-->1	.->2	b->4	e->18	k->1	l->1	m->1	n->289	
gerk	r->1	
gerl	i->3	
germ	a->1	
gern	 ->9	,->2	.->3	a->8	s->7	
gerp	o->2	
gers	 ->1	
gerv	r->1	
ges 	a->3	b->1	d->3	e->2	f->1	i->7	k->1	n->2	o->1	p->1	s->1	t->2	u->1	y->1	ä->1	ö->1	
ges,	 ->3	
ges-	 ->1	
ges.	R->1	
gesb	e->1	
gesf	o->1	
gesr	a->2	
gest	 ->1	?->1	u->7	ä->3	
get 	(->2	-->2	1->1	A->1	R->1	a->21	b->5	e->6	f->20	g->10	h->8	i->21	k->10	l->6	m->10	n->2	o->25	p->8	r->3	s->41	t->24	u->5	v->7	y->1	ä->10	ö->2	
get)	 ->1	,->1	.->2	
get,	 ->28	
get.	 ->1	A->1	D->9	E->2	F->4	H->2	I->2	J->8	K->2	L->1	M->5	N->1	O->2	P->2	S->2	T->1	V->1	
get:	 ->1	
get;	 ->1	
get?	V->1	
geta	n->1	r->2	
getb	e->1	
getd	e->1	
gete	c->2	n->15	r->1	
getf	r->2	ö->9	
getk	o->16	r->1	
getm	ä->1	
getp	l->3	o->11	
gets	 ->25	i->1	t->2	y->1	
gett	 ->24	,->1	
getu	t->10	
getå	r->10	
getö	v->1	
gfal	d->15	
gflö	d->1	
gfon	d->1	
gfor	s->20	
gfri	s->1	
gfru	t->1	
gfun	k->1	
gfär	d->1	g->1	
gför	s->5	
gg d	e->1	ä->1	
gg f	a->1	r->1	
gg g	e->1	
gg h	a->2	
gg i	 ->3	n->2	
gg k	u->1	
gg l	å->1	
gg m	a->1	ä->1	
gg o	c->1	
gg p	å->3	
gg s	o->2	
gg t	i->4	
gg u	n->2	p->1	t->1	
gg v	i->1	
gg" 	s->1	
gg, 	e->3	i->1	k->1	m->1	t->1	v->1	
gg.D	ä->1	
gg.F	ö->2	
gg.K	o->1	
gg.M	a->1	
gg.N	u->1	
gg; 	f->1	
gga 	I->1	a->9	b->2	d->4	e->7	f->48	g->1	h->2	i->5	k->3	m->1	n->4	o->6	p->2	r->2	s->8	t->11	u->20	v->7	ö->1	
gga,	 ->1	
ggad	e->3	
ggan	 ->2	d->109	
ggas	 ->11	,->2	.->1	
ggbo	x->1	
ggd 	i->1	p->1	
ggde	 ->1	s->1	
gge 	s->1	
ggel	s->1	
ggen	 ->6	"->1	s->1	
gger	 ->127	,->3	.->2	;->1	
gget	 ->3	,->1	s->2	
gghe	t->6	
ggig	t->3	
ggjo	r->13	
ggli	n->1	
ggna	d->19	
ggni	n->28	
ggor	 ->1	n->1	
ggra	d->1	n->12	
ggre	s->1	
ggs 	f->7	i->3	n->1	p->5	u->2	v->1	
ggs,	 ->1	
ggsb	u->1	
ggsf	r->1	
ggsk	r->1	
ggst	e->1	
ggt 	i->1	p->1	s->1	u->1	
ggts	 ->1	
ggå 	l->1	
ggås	,->1	
ggör	 ->5	a->12	s->4	
gh l	e->1	
gh m	e->1	
gh.V	i->1	
ghet	 ->225	!->1	"->1	,->35	.->40	?->1	e->466	s->82	
ght 	k->1	t->1	
ghts	.->1	
ghål	l->2	
gi -	 ->2	
gi b	e->1	
gi f	ö->5	
gi g	e->1	ö->1	
gi h	a->2	
gi i	 ->1	
gi k	a->1	
gi l	e->1	
gi m	e->1	å->1	
gi o	c->8	
gi s	o->7	
gi t	i->2	
gi, 	d->1	e->1	i->1	k->1	m->1	o->1	
gi-,	 ->1	
gi..	 ->1	
gi.A	l->1	
gi.D	e->1	
gi.E	t->1	u->1	
gi.F	o->1	r->1	
gi.J	a->1	
gi.M	a->1	
gi.V	å->1	
giag	e->1	
gian	v->6	
gibe	s->3	
gice	n->1	
gick	 ->18	,->2	.->2	
gief	f->4	
gien	 ->5	,->3	.->1	?->1	s->1	
gier	 ->11	,->4	.->1	a->1	n->1	
giet	,->1	.->1	
gifo	r->1	
gift	 ->22	!->1	,->2	.->6	:->1	e->59	i->2	s->8	
gifö	r->4	
giga	n->5	
gigg	j->1	
gigt	 ->2	,->1	.->1	
giim	p->1	
gik 	o->1	
gik,	 ->2	
gik.	F->1	H->1	V->1	
gika	p->1	
gike	n->2	
giko	n->1	
gikä	l->37	
gill	a->2	
gilt	i->26	
gime	n->3	
gimi	x->1	
gimy	n->1	
gin 	f->2	k->1	m->1	o->2	s->1	u->1	
gin,	 ->2	
gin.	D->1	S->1	
gina	l->7	
gine	l->1	
gins	 ->1	
ginä	r->1	
gion	 ->12	,->3	.->7	a->89	e->141	
gior	g->2	
gipl	a->1	
gipo	l->1	t->1	
gipr	o->5	
gise	k->4	
gisi	s->70	
gisk	 ->10	a->39	t->17	
gisn	å->1	
giss	l->1	
gist	e->10	r->10	
gisä	k->7	
git 	-->1	a->5	b->3	d->7	e->10	f->5	h->8	i->7	k->1	l->2	m->3	n->4	o->2	p->4	s->8	t->8	u->13	v->3	ä->1	å->1	
git,	 ->2	
git.	F->3	I->1	M->1	
gita	t->1	
giti	m->18	
gits	 ->22	,->2	.->3	
gium	 ->2	.->1	
giva	n->12	r->51	
give	n->5	r->1	s->1	t->25	
givi	t->15	
givl	i->1	
givn	a->5	i->6	
gizi	s->5	
giäk	e->1	
giåt	e->1	
giös	 ->1	a->2	t->1	
gjor	d->41	t->95	
gkra	s->3	
gkul	t->1	
gkör	n->1	
gla 	d->2	m->1	p->4	
glad	 ->20	a->3	d->2	e->5	
glan	d->1	
glar	 ->15	,->3	.->1	
glas	 ->3	.->1	h->1	
gled	a->3	n->2	
gler	 ->39	,->10	.->6	?->1	a->19	i->15	n->36	
gles	a->1	
glew	o->2	
glig	 ->8	,->1	.->1	a->43	e->11	h->4	t->19	
glin	g->2	
glju	d->1	
glob	a->12	
glup	s->1	
gläd	e->19	j->15	s->6	
glän	g->1	
glöm	m->16	s->1	t->4	
gm e	l->1	
gmar	 ->1	
gmat	i->3	
gmet	a->6	
gmär	k->1	
gmäs	t->2	
gmål	,->1	
gn f	ö->3	
gn o	c->1	
gna 	a->9	b->2	d->2	e->2	f->9	g->2	i->9	k->3	l->2	m->8	n->4	o->6	p->6	r->3	s->16	t->1	u->1	v->3	ä->3	å->5	ö->1	
gna,	 ->3	
gna.	D->1	I->1	
gnad	 ->6	.->1	e->14	s->3	
gnal	 ->9	e->5	
gnan	d->1	
gnar	 ->24	,->3	.->4	
gnas	 ->2	.->1	
gnat	 ->5	i->1	s->1	
gne 	f->2	i->1	o->2	s->3	
gne-	A->1	
gnel	s->1	
gnen	 ->2	
gner	.->1	a->2	
gnes	 ->1	
gni,	 ->1	
gnin	g->223	
gnis	k->1	
gnit	u->1	
gniv	å->3	
gnor	e->4	
gnut	t->2	
gnäl	l->1	
go g	r->1	
go s	o->1	
go å	r->1	
god 	a->2	b->1	f->6	i->3	j->1	l->1	m->1	t->6	u->1	v->1	
god.	F->1	
goda	 ->36	.->1	
godk	ä->89	
godo	.->3	s->1	
gods	 ->29	,->1	.->4	;->1	N->1	e->2	
godt	a->38	o->2	y->6	
gofe	m->1	
goge	r->1	
gogi	 ->1	.->2	s->1	
gois	t->2	
golf	e->4	
golv	e->1	
goly	c->1	
gom 	a->1	u->1	ä->2	
gom.	D->1	
gomå	l->3	
gon 	a->15	b->7	c->1	d->4	e->8	f->4	g->7	h->1	i->4	j->2	k->25	l->4	m->5	n->5	o->3	p->5	r->8	s->19	t->7	u->3	v->2	ä->2	å->1	
gon,	 ->5	
gon.	A->1	D->1	H->1	I->1	J->1	V->2	
gonb	l->15	
gond	a->2	e->1	
gons	i->11	t->4	
gont	i->39	
gor 	-->1	F->1	a->10	b->6	d->3	e->4	f->4	g->4	h->6	i->12	k->1	l->1	m->4	o->41	p->3	s->54	t->12	u->2	v->8	ä->5	
gor)	 ->1	
gor,	 ->38	
gor.	 ->1	.->1	D->10	F->4	H->1	J->2	K->2	M->1	N->2	S->1	V->3	
gor:	 ->4	
gor;	 ->1	
gor?	,->1	Ä->1	
gord	n->52	
gori	 ->3	e->5	s->1	
gorl	u->1	
gorn	a->31	
gors	 ->2	
gorö	s->4	
gosk	r->1	
gosl	a->1	
got 	E->1	K->1	W->1	a->22	b->3	d->3	e->3	f->15	h->1	i->4	j->4	k->2	l->6	m->10	o->10	p->5	r->2	s->75	t->4	u->2	v->10	å->1	
got,	 ->2	
got.	A->1	D->2	J->1	S->1	Ä->1	
got?	N->1	
gott	 ->17	.->1	e->1	g->1	
gou 	o->1	
gpla	n->1	t->3	
gpol	i->2	
gra 	-->1	a->24	b->5	d->5	e->7	f->11	g->6	h->2	i->6	k->11	l->1	m->9	n->3	o->7	p->9	r->2	s->20	t->7	u->3	v->7	ä->3	å->8	ö->1	
grad	 ->16	,->1	.->2	e->15	v->3	
graf	 ->1	i->14	r->2	
gram	 ->75	,->17	.->20	?->2	a->1	f->1	m->108	p->11	r->1	u->1	v->1	
gran	 ->5	d->5	n->8	s->55	t->12	
grar	 ->5	a->1	
gras	 ->1	
grat	 ->4	i->28	s->1	u->36	
grav	a->1	e->4	t->1	
gre 	B->1	a->2	b->2	c->1	e->1	f->6	g->4	h->1	i->3	k->8	m->1	n->5	o->4	p->7	r->1	s->11	t->10	u->3	v->4	ä->7	
gre,	 ->1	
gre.	D->1	F->1	I->1	M->1	N->1	R->1	S->1	V->1	Ä->1	
gred	i->2	
grek	e->1	i->6	
grem	s->1	
gren	,->1	a->2	s->1	
grep	 ->1	p->25	
grer	a->18	i->6	
gres	s->3	u->1	
grif	i->1	
grik	e->1	
grin	g->1	
grip	a->37	e->19	i->2	l->6	n->1	s->1	
grit	e->3	
grod	d->1	
grog	r->1	
grot	u->1	
grou	p->1	
grov	 ->1	
grun	d->297	
grup	p->184	
gruv	a->1	
grym	t->1	
gräl	 ->2	,->1	
gräm	e->1	
grän	s->134	
gräv	a->3	e->1	
grå 	v->1	
gråz	o->1	
gröd	o->1	
gröj	a->1	
grön	 ->2	a->14	b->1	t->1	
gröv	s->1	
gs -	,->1	
gs a	l->1	n->1	t->8	v->4	
gs b	o->1	r->1	
gs d	a->1	e->3	i->1	
gs e	m->1	n->2	
gs f	a->2	r->7	y->1	ö->5	
gs g	e->1	
gs h	ä->2	
gs i	 ->6	d->1	g->1	n->3	
gs k	l->2	u->1	
gs m	e->4	å->1	
gs n	u->1	ä->1	
gs o	c->2	m->3	
gs p	o->1	r->1	å->7	
gs r	a->1	e->1	
gs s	i->1	k->4	o->1	t->1	
gs t	i->1	
gs u	n->2	p->3	t->2	
gs v	a->1	e->1	i->2	
gs, 	1->1	a->1	f->1	m->1	u->1	
gs- 	f->1	o->11	
gs.F	ö->1	
gs.J	a->1	
gs.L	å->1	
gsak	t->3	
gsal	t->1	
gsam	 ->2	h->2	m->6	t->3	
gsan	a->1	f->1	l->4	s->2	
gsar	b->6	t->3	
gsav	g->1	t->6	v->1	
gsba	r->2	
gsbe	d->1	h->1	l->1	s->5	t->1	v->4	
gsbi	d->2	l->7	s->2	
gsbo	l->2	r->2	
gsbr	u->6	
gsbu	d->1	
gsce	n->5	
gsch	e->8	
gsde	l->1	
gsdi	r->2	
gsdo	k->1	
gsdr	a->1	
gsek	o->5	t->1	
gsen	 ->2	h->1	
gser	a->1	b->1	
gset	 ->4	a->1	
gsfa	k->1	l->1	r->2	s->5	
gsfe	l->2	
gsfi	e->30	n->1	
gsfl	y->1	
gsfo	n->21	r->1	
gsfr	ä->2	å->14	
gsfu	l->11	n->1	
gsfä	s->1	
gsfö	r->235	
gsgi	v->8	
gsgr	a->3	u->5	
gsha	n->1	
gshe	r->1	
gsho	t->1	
gsid	i->3	k->1	
gsik	t->7	
gsin	d->4	f->1	i->1	s->5	t->1	
gsju	r->2	
gska	p->1	
gskl	a->2	i->1	
gsko	a->2	l->1	m->25	n->135	r->2	s->8	
gskr	a->15	i->1	
gsku	r->1	
gskv	o->1	
gskä	l->2	
gsla	g->1	n->1	
gsli	g->1	n->2	s->47	v->10	
gslo	g->1	
gslä	g->5	n->3	
gslö	s->5	
gsma	j->1	k->1	r->2	
gsme	d->2	k->2	t->3	
gsmi	n->1	
gsmo	d->2	m->1	n->1	t->1	
gsmä	s->4	
gsmå	l->4	
gsmö	j->3	n->1	
gsna	 ->4	,->1	r->1	
gsne	d->1	
gsni	v->5	
gsno	r->1	
gsny	c->1	
gsnä	t->2	
gsom	r->12	
gsor	g->2	
gspa	k->1	n->1	r->2	
gspe	r->3	
gspl	a->17	i->6	
gspo	l->22	
gspr	i->1	o->45	
gspu	n->11	
gspå	f->1	
gsre	f->1	g->7	k->5	p->2	s->8	
gsri	k->15	
gsru	n->1	
gsrä	d->1	t->1	
gsrå	d->3	
gssa	m->2	
gsse	d->1	k->7	
gssi	f->1	t->2	
gssk	a->3	e->3	i->5	r->8	y->3	
gssp	r->1	
gsst	a->2	r->15	å->1	ö->5	
gssy	s->24	
gssä	k->2	l->6	t->8	
gst 	a->3	b->1	f->1	g->1	k->2	o->1	p->2	r->1	t->1	u->1	
gst,	 ->1	
gst.	V->1	
gsta	 ->19	d->1	g->7	n->1	
gste	n->4	x->2	
gsti	d->2	f->127	l->2	
gstj	ä->5	
gstm	ä->2	
gstr	ö->1	
gstä	l->1	t->1	
gsum	m->1	
gsut	r->5	s->1	ö->1	
gsve	r->4	
gsvi	l->3	s->30	
gsvä	n->1	r->5	v->1	
gsvå	g->1	r->1	
gsys	t->2	
gsäg	a->3	
gsän	d->3	
gsär	e->1	
gsät	t->1	
gsår	e->1	
gsåt	g->5	
gsöv	e->1	
gt -	 ->7	
gt 4	0->1	8->1	
gt :	 ->1	
gt D	u->1	
gt E	u->2	
gt G	r->1	
gt I	n->1	
gt K	y->1	
gt R	a->1	
gt S	c->1	
gt T	h->1	
gt a	d->1	l->3	n->5	r->14	s->1	t->197	v->21	
gt b	a->2	e->20	i->4	l->1	o->1	r->4	ä->1	å->1	
gt d	a->1	e->30	i->3	j->1	r->1	ä->2	
gt e	d->1	f->10	g->1	l->4	n->7	r->3	t->4	u->1	x->5	
gt f	a->2	e->3	i->2	l->2	o->2	r->38	u->1	å->1	ö->78	
gt g	e->3	o->40	r->3	ä->1	
gt h	a->15	e->1	i->1	j->1	o->5	u->1	ä->3	å->1	ö->5	
gt i	 ->24	c->1	f->6	n->24	
gt j	a->2	u->1	
gt k	a->4	l->1	n->1	o->16	r->4	v->2	ä->2	
gt l	i->5	ä->7	å->3	
gt m	a->1	e->35	i->38	o->3	y->5	ä->1	å->11	ö->3	
gt n	a->1	e->9	i->1	o->8	ä->6	å->1	
gt o	a->4	b->2	c->59	f->3	m->4	r->6	s->1	t->2	
gt p	a->5	e->1	l->1	o->4	r->19	å->9	
gt r	e->11	u->9	y->1	ä->1	
gt s	a->9	e->4	i->7	j->1	k->15	l->2	n->1	o->27	p->2	t->37	u->1	v->4	y->6	ä->32	å->1	
gt t	a->11	e->2	i->14	o->1	v->1	y->2	ä->1	
gt u	n->6	p->10	r->1	t->9	
gt v	a->6	e->1	i->30	ä->5	å->6	
gt y	t->2	
gt ä	n->2	r->14	v->1	
gt å	t->3	
gt ö	g->1	n->1	v->4	
gt!L	e->1	
gt!M	e->1	
gt, 	a->1	b->2	d->4	e->5	f->6	h->2	i->4	j->3	k->6	l->2	m->5	n->2	o->12	p->1	r->1	s->9	u->3	v->2	ä->3	
gt. 	I->1	
gt.A	r->1	
gt.D	e->11	i->1	
gt.E	f->1	n->1	t->1	
gt.F	r->2	ö->6	
gt.G	e->2	
gt.H	e->4	u->1	
gt.I	 ->1	
gt.J	a->12	
gt.L	å->2	
gt.M	a->1	e->5	i->3	o->1	
gt.N	a->1	ä->1	
gt.O	f->1	m->2	
gt.P	å->1	
gt.S	e->1	o->1	t->2	
gt.U	n->1	
gt.V	a->5	i->9	
gt.Ö	k->1	
gt: 	d->1	
gt; 	d->1	
gt?A	v->1	
gtar	 ->1	
gtek	n->2	
gter	a->8	
gtex	t->2	
gtgå	e->11	
gtid	l->4	s->4	
gton	 ->2	.->1	?->1	s->1	
gtra	n->2	
gts 	-->2	8->1	a->5	b->1	f->17	h->3	i->3	n->1	o->1	t->1	u->2	
gts,	 ->2	
gtvi	s->108	
gtvä	t->4	
guds	 ->2	
gue,	 ->1	
guei	r->1	
guer	 ->2	
gues	a->1	
guld	e->1	
gult	 ->1	
gume	n->17	
gumm	i->1	
guro	,->1	
gust	a->1	
guve	r->1	
gvar	i->6	
gvat	t->1	
gver	k->1	
gynn	a->16	s->3	
gypt	e->2	
gäck	 ->1	
gäld	 ->1	
gäll	a->29	d->11	e->362	n->1	t->2	
gäng	e->1	l->23	
gär 	a->3	b->1	d->1	e->3	o->1	s->1	ö->1	
gär.	V->1	
gära	 ->9	,->1	n->21	s->3	
gärd	 ->13	,->6	.->5	;->1	a->3	e->210	s->10	
gärn	a->32	i->1	
gärs	 ->1	
gärt	 ->7	,->2	.->1	
gäve	s->1	
gå K	i->1	
gå a	n->1	t->1	
gå b	e->2	
gå d	e->2	
gå e	n->3	t->2	
gå f	r->6	ö->3	
gå g	r->2	
gå h	e->1	
gå i	 ->8	g->4	n->15	
gå l	a->1	ä->4	å->1	
gå m	e->3	
gå o	c->2	f->1	
gå p	å->1	
gå s	a->1	n->1	o->2	å->3	
gå t	i->13	
gå u	n->1	t->4	
gå v	i->4	
gå å	t->1	
gå.A	t->1	
gå.D	ä->1	
gå.F	ö->1	
gå.N	ä->1	
gå.O	m->1	
gå.S	o->1	
gå.V	i->1	
gåen	d->101	
gång	 ->109	"->1	,->8	.->13	a->13	e->68	k->1	n->2	s->44	
går 	a->9	b->5	d->15	e->3	f->10	g->2	h->3	i->23	j->2	k->1	l->3	m->7	n->2	o->10	p->4	r->1	s->6	t->17	u->12	v->3	ä->1	å->2	ö->1	
går,	 ->4	
går.	 ->1	D->1	I->1	J->2	V->3	
gård	 ->1	a->4	e->1	
gås 	a->1	i->2	o->1	
gås,	 ->1	
gås:	 ->1	
gått	 ->30	.->3	s->3	
gåvo	r->2	
gömm	a->1	e->2	
gömt	s->1	
gör 	"->1	3->1	8->1	E->1	a->30	b->1	d->56	e->20	f->4	g->5	h->6	i->5	k->2	m->11	n->7	o->4	p->4	r->1	s->8	t->4	u->3	v->10	y->1	ä->4	
gör,	 ->2	
gör.	D->3	E->1	
göra	 ->276	,->7	.->13	?->1	n->58	s->34	
göre	l->5	
göri	n->2	
görl	i->2	
görs	 ->21	,->4	.->3	
h "U	r->1	
h "s	k->1	
h "t	i->1	
h (A	5->1	
h - 	e->1	s->2	
h -o	r->3	
h 0 	p->1	
h 1-	2->1	
h 10	 ->1	0->1	
h 13	8->1	
h 14	 ->1	
h 16	 ->1	
h 17	 ->1	.->1	
h 19	 ->1	4->1	9->11	
h 2 	i->1	
h 2,	 ->1	
h 2.	D->1	
h 20	 ->2	0->1	
h 21	 ->3	
h 22	.->1	
h 25	.->1	
h 27	 ->1	
h 29	 ->1	
h 3.	I->1	
h 30	 ->1	0->1	
h 33	 ->1	
h 34	 ->1	
h 35	.->1	
h 3:	 ->1	
h 4.	J->1	
h 41	 ->2	
h 45	 ->2	,->1	.->1	
h 47	 ->1	
h 48	 ->2	
h 5 	v->1	
h 5.	E->1	
h 53	 ->1	
h 60	-->1	
h 68	 ->1	
h 7 	-->1	f->1	i->1	o->1	
h 7,	 ->2	
h 8 	ä->1	
h 8,	 ->1	
h 82	 ->2	)->1	,->3	
h 86	 ->2	
h 89	 ->1	
h 9 	i->1	m->1	
h 92	/->1	
h 94	 ->1	
h Al	b->1	t->1	
h Am	s->1	
h An	k->1	
h BP	,->1	
h Ba	s->1	
h Be	l->1	
h Br	a->1	o->1	
h Bu	l->1	
h C.	 ->1	
h CE	C->1	
h Ca	u->1	
h Cy	p->1	
h Da	n->2	
h De	 ->1	m->1	
h EL	D->2	
h EU	 ->2	-->1	G->1	
h Ed	i->1	
h El	m->2	
h Em	i->1	
h Er	k->1	
h Et	i->1	
h Eu	r->24	
h FN	:->1	
h FP	Ö->1	
h Fi	n->2	
h Fr	a->10	u->1	
h Ga	l->1	z->1	
h Ge	m->1	
h Go	l->1	
h Gr	a->1	e->1	u->1	
h He	l->1	
h Hi	t->1	
h Hu	h->1	
h II	 ->1	,->1	
h In	d->2	t->2	
h Ir	l->2	
h Is	r->5	
h It	a->1	
h Ja	c->1	
h Jö	r->1	
h Ka	s->1	
h Ki	n->5	r->1	
h Ko	u->1	
h Ku	l->1	
h La	n->3	
h Le	i->5	
h MA	R->1	
h Ma	d->3	
h Me	d->1	
h No	r->1	
h Ny	a->1	
h OL	A->1	
h On	e->1	
h PP	E->1	
h PS	E->2	
h Pa	c->1	k->3	l->4	r->1	
h Pe	t->1	
h Po	r->3	
h Pr	í->1	
h Ra	f->2	p->1	
h Sa	m->10	
h Sc	h->2	
h Si	m->1	
h Sj	ö->1	
h So	c->1	
h Sp	a->1	
h St	o->2	
h Sw	o->1	
h Sy	d->1	r->7	
h Ta	d->1	i->1	m->2	
h Ts	a->1	
h Tu	r->1	
h Ty	s->2	
h Uz	b->1	
h Vi	t->1	
h Vä	s->1	
h Wy	e->1	
h X 	o->1	
h ab	s->1	
h ac	c->1	
h ad	m->1	v->1	
h ag	e->2	
h ak	t->4	
h al	d->2	l->16	
h am	b->4	
h an	a->3	d->27	g->3	n->3	p->2	s->12	t->5	v->3	
h ap	r->1	
h ar	b->14	t->1	
h as	s->1	y->3	
h at	t->150	
h av	 ->14	d->1	g->3	l->1	r->2	s->6	t->3	v->2	
h ba	d->1	g->1	l->3	n->1	r->7	
h be	a->1	d->8	f->7	g->2	h->7	k->4	l->4	m->1	r->3	s->5	t->6	v->4	
h bi	d->6	l->4	
h bl	.->2	a->2	i->3	u->1	
h bo	r->2	s->2	t->1	
h br	a->1	i->2	o->2	u->2	ä->3	å->5	
h bu	d->3	
h by	r->2	
h bä	s->2	t->2	
h bå	t->1	
h bö	r->6	
h ca	l->1	n->1	
h ce	n->6	
h ch	e->1	o->1	
h da	g->2	m->1	t->1	
h de	 ->83	b->2	c->1	l->8	m->10	n->108	r->12	s->35	t->208	
h di	a->1	o->1	r->3	s->4	t->2	
h dj	u->3	ä->1	
h do	m->9	
h dr	a->2	i->2	
h du	k->1	
h dy	r->1	
h dä	r->83	
h då	 ->22	,->1	l->1	
h dö	t->1	
h ef	f->16	t->18	
h eg	e->1	
h ej	 ->1	
h ek	o->22	
h el	e->1	
h en	 ->70	,->1	a->1	d->2	e->2	g->2	h->5	k->1	l->2	s->1	t->2	v->1	
h er	 ->2	.->1	a->2	b->2	f->3	h->1	k->2	s->3	t->1	
h et	i->1	t->32	
h eu	r->9	
h ex	a->2	p->1	t->1	
h fa	k->2	l->2	r->3	s->1	t->5	u->1	
h fe	d->1	l->1	m->1	
h fi	e->1	n->8	r->1	s->2	
h fl	e->8	o->1	y->1	
h fo	d->1	l->2	r->4	
h fr	a->25	e->2	i->6	o->2	u->4	ä->34	å->10	
h fu	l->5	n->2	s->2	
h fy	r->1	s->1	
h fä	l->1	
h få	 ->4	g->1	r->5	t->2	
h fö	l->5	r->163	
h ga	g->1	r->6	
h ge	 ->10	m->6	n->20	o->1	r->3	s->3	
h gi	v->4	
h gj	o->1	
h gl	a->1	o->1	ä->1	
h go	d->1	t->1	
h gr	a->2	u->5	ä->2	ö->1	
h gä	l->1	
h gå	 ->2	r->2	
h gö	r->17	
h ha	 ->2	m->1	n->27	r->16	
h he	l->7	n->4	r->43	
h hi	t->1	
h hj	ä->4	
h ho	b->1	n->1	p->5	t->4	
h hu	m->1	n->1	r->11	s->1	v->1	
h hy	g->1	l->1	
h hä	l->1	r->8	
h hå	l->16	
h hö	g->4	j->2	
h i 	G->1	M->1	N->1	S->1	T->2	a->1	b->1	d->13	e->3	f->5	g->4	h->1	i->1	j->1	k->1	l->1	m->1	n->1	o->1	p->2	r->1	s->16	u->2	v->8	ö->4	
h ib	l->3	
h ic	k->2	
h id	e->2	r->3	
h if	r->1	
h ik	r->1	
h il	l->1	
h im	a->1	m->1	
h in	d->6	f->11	g->7	h->1	i->2	k->1	l->1	n->3	o->7	p->1	r->12	s->12	t->72	v->6	
h ir	l->1	
h is	r->2	
h ja	g->149	
h jo	r->5	
h ju	r->3	s->4	
h jä	m->1	
h ka	b->1	m->1	n->14	p->1	r->2	t->2	
h ki	n->1	
h kl	a->3	o->1	
h kn	u->1	
h ko	h->1	l->2	m->61	n->57	r->5	s->3	
h kr	a->5	e->1	i->6	y->1	ä->4	å->1	
h ku	l->3	n->4	
h kv	a->2	i->8	
h kä	l->1	m->1	r->4	
h kö	r->1	
h la	g->6	n->10	r->1	
h le	d->13	g->1	m->1	v->2	
h li	k->7	t->1	v->3	
h lj	u->1	
h lo	c->1	k->4	s->1	v->3	
h lu	k->1	
h ly	c->3	
h lä	c->1	g->6	m->2	n->1	r->1	t->3	
h lå	n->11	s->1	t->7	
h lö	s->2	
h ma	k->1	n->18	r->1	t->1	
h me	d->122	k->1	l->3	n->2	r->15	t->1	
h mi	g->1	l->18	n->17	s->3	
h mo	d->4	n->6	r->3	t->11	
h mu	s->1	
h my	c->7	n->1	
h mä	n->11	r->1	
h må	h->1	l->6	n->10	s->5	
h mö	j->8	r->1	
h na	t->11	
h ne	d->1	g->1	o->1	p->4	u->1	
h ni	 ->8	v->1	
h no	g->3	r->1	t->1	
h nu	 ->11	
h ny	a->5	e->1	l->3	n->2	t->2	
h nä	m->1	r->14	t->2	
h nå	g->5	
h nö	d->6	
h oa	c->4	
h ob	e->2	
h oc	h->2	k->8	
h od	e->1	
h oe	g->1	k->1	
h of	f->3	t->2	ö->1	
h oj	ä->1	
h ok	l->3	r->1	
h ol	i->5	j->1	y->2	
h om	 ->22	b->2	e->3	f->5	g->3	r->2	s->4	
h on	t->1	
h op	e->1	p->1	
h or	d->3	g->2	i->1	s->1	ä->1	
h os	s->2	t->1	ä->2	
h ot	v->1	
h ou	m->1	n->1	t->1	
h pa	p->1	r->23	s->1	
h pe	k->2	r->7	
h pl	a->1	i->2	
h po	l->15	s->2	
h pr	a->1	e->3	i->8	o->19	ä->1	
h på	 ->22	m->1	p->1	s->2	t->1	v->2	
h ra	p->1	s->4	t->2	
h re	c->1	d->2	f->4	g->34	j->1	k->2	l->3	n->5	p->1	s->11	v->2	
h ri	g->1	k->6	n->1	s->1	
h ro	l->1	m->3	
h ru	t->1	
h rä	d->1	k->1	t->59	
h rå	d->39	
h rö	s->1	
h sa	m->40	n->3	
h se	 ->6	d->9	k->3	l->1	n->1	r->5	t->1	x->3	
h si	f->1	n->3	s->3	t->3	
h sj	u->1	ä->3	ö->2	
h sk	a->14	i->1	o->1	r->1	u->3	y->4	ä->2	ö->4	
h sl	a->1	u->20	ä->3	
h sm	u->1	å->1	
h sn	a->3	å->1	
h so	c->40	l->2	m->92	
h sp	a->1	e->4	r->4	
h st	a->12	i->1	o->3	r->19	ä->7	å->5	ö->14	
h su	c->1	v->4	
h sv	a->4	å->8	
h sy	f->2	n->1	r->1	s->12	
h sä	g->7	k->12	n->1	r->11	t->2	
h så	 ->21	d->4	l->2	s->1	
h sö	d->1	r->1	
h t.	o->1	
h ta	 ->5	c->6	k->1	l->4	n->1	r->1	s->2	
h te	k->2	l->4	
h th	e->1	
h ti	d->3	g->1	l->52	n->2	s->1	t->1	
h tj	o->1	ä->3	
h to	g->1	l->3	p->1	t->1	
h tr	a->9	e->2	o->5	å->2	
h tu	n->1	r->14	s->2	
h tv	å->3	
h ty	d->13	v->1	
h tä	m->1	n->1	p->1	
h un	d->17	g->6	i->2	
h up	p->24	
h ut	a->5	b->4	e->1	f->2	g->4	i->1	l->1	n->2	o->1	r->2	s->4	t->3	v->26	ö->1	
h va	d->10	l->13	n->4	p->3	r->22	
h ve	k->1	m->2	r->9	t->11	
h vi	 ->86	a->1	d->6	k->3	l->13	n->1	s->13	
h vä	d->1	g->2	l->12	n->2	p->1	r->4	x->4	
h vå	l->1	r->11	
h vö	r->1	
h yn	g->1	
h yr	k->1	
h yt	l->1	t->4	
h ÖV	P->1	
h Ös	t->6	
h äg	a->1	n->1	
h än	 ->4	d->5	n->3	
h är	 ->9	e->1	
h äv	e->31	
h å 	a->4	
h åk	l->1	
h ås	a->1	i->1	t->1	
h åt	e->26	g->3	
h ök	a->3	
h öm	s->1	
h ön	s->1	
h öp	p->13	
h ör	e->1	
h ös	t->4	
h öv	e->16	r->4	
h! U	r->1	
h)De	t->1	
h, a	t->1	
h, d	e->1	
h, f	r->1	ö->2	
h, h	e->1	
h, i	 ->1	
h, n	å->1	
h, o	r->1	
h, r	e->1	
h, s	l->1	o->3	
h, t	r->1	
h, u	t->1	
h-Be	h->7	
h-av	t->1	
h.De	t->1	
h.Ef	t->1	
h.Fö	r->1	
h.Ja	g->1	
h.Vi	 ->1	
h/el	l->1	
h: V	e->1	
h?Fr	u->1	
hI o	k->1	
hII.	 ->1	
ha a	n->3	r->1	t->1	
ha b	e->4	r->1	
ha d	e->7	i->1	r->1	ö->1	
ha e	g->1	n->36	r->1	t->17	
ha f	r->3	u->1	ö->2	
ha g	e->2	j->2	r->1	
ha h	a->2	i->1	ö->4	
ha i	 ->1	n->2	
ha k	l->1	o->5	u->2	v->1	ä->1	
ha l	y->3	ä->1	
ha m	a->2	e->2	i->1	o->2	y->2	ö->3	
ha n	e->1	y->1	å->8	
ha o	c->1	f->1	
ha p	r->2	
ha r	ä->2	å->1	
ha s	a->4	e->1	j->1	k->3	t->3	u->1	y->1	
ha t	a->1	i->4	r->1	v->3	y->2	
ha u	n->2	p->1	t->2	
ha v	a->7	e->1	i->3	ä->3	
ha y	t->1	
ha ä	g->1	n->1	
ha å	s->1	
ha ö	n->2	v->1	
ha, 	e->1	
ha.A	l->1	
habi	l->1	
habl	o->1	
hade	 ->84	?->1	
haft	 ->34	,->2	.->1	
hagl	i->2	
haka	t->1	
hall	"->1	
halt	 ->1	
halv	 ->3	a->4	h->1	m->1	o->1	t->5	v->2	å->5	ö->3	
hamb	u->1	
hame	l->1	
hamm	a->1	
hamn	 ->4	.->1	a->28	b->1	e->2	i->1	k->2	
hamp	a->1	
han 	a->6	b->3	d->2	e->1	f->5	g->3	h->22	i->14	j->2	k->7	l->5	m->2	n->3	o->3	p->3	s->12	t->5	u->3	v->6	ä->9	ö->1	
han,	 ->2	
han;	 ->1	
hand	 ->47	,->4	.->3	?->1	a->46	e->36	f->1	i->4	l->348	s->17	u->2	
hang	 ->20	,->6	.->8	e->13	
hank	a->1	
hans	 ->82	e->6	
hant	e->41	v->2	
hape	a->1	
happ	y->1	
har 	-->2	1->2	4->1	A->1	B->1	E->7	G->1	L->2	P->1	S->1	a->85	b->78	c->2	d->97	e->98	f->171	g->92	h->61	i->102	j->39	k->55	l->91	m->67	n->63	o->30	p->37	r->53	s->131	t->72	u->54	v->140	ä->21	å->4	ö->12	
har"	 ->1	
har,	 ->14	
har.	D->1	T->1	
har:	 ->1	
har?	N->1	
hara	d->1	s->1	
hard	 ->1	-->1	
harm	 ->4	-->1	a->1	o->18	
hart	r->1	
has 	b->1	
hast	a->3	i->1	
hat 	o->1	
hate	t->2	
hati	s->1	
hatt	e->1	
haus	s->1	
hav 	f->1	o->1	
hav,	 ->1	
hava	n->1	r->3	
have	n->4	r->7	t->16	
havs	 ->4	,->4	.->4	?->1	f->2	l->1	m->2	o->1	v->1	
he B	a->1	
he R	o->1	
he c	i->1	
he i	m->1	
he o	c->1	
he, 	L->1	
head	-->1	
heat	o->21	
hebr	e->1	
heck	 ->1	
hede	r->3	
hedr	a->5	
heer	 ->3	,->4	J->1	b->3	s->3	
hef 	h->1	
hefe	n->1	r->15	
heik	.->1	h->4	
hejd	a->2	
hekt	a->2	
hel 	b->1	d->6	k->1	p->1	r->2	
hela	 ->105	
helg	e->1	
helh	e->21	j->8	
heli	g->1	
hell	 ->2	e->47	r->6	
helm	s->1	
hels	i->1	t->46	
helt	 ->135	,->1	.->3	ä->4	
hem 	e->1	f->1	o->2	t->1	ä->1	
hem.	 ->1	N->1	
hema	 ->1	
hemb	y->1	
hemf	ö->1	
heml	a->3	i->5	ä->2	ö->5	
hemm	a->9	e->1	
hems	k->5	
hemv	i->1	
hen 	f->3	h->1	i->1	s->1	v->1	
hen,	 ->1	
hen.	F->1	
hen;	 ->1	
heng	e->10	
henn	e->27	
hens	 ->2	
heph	e->3	
her 	i->1	o->1	v->1	
her"	 ->1	
hera	n->1	r->1	
herd	s->3	
here	n->1	
hern	 ->5	,->3	a->2	
hero	i->1	
herr	 ->165	a->45	
hes 	i->1	
het 	-->1	1->1	D->1	R->1	S->1	a->63	b->10	d->12	e->16	f->57	g->3	h->10	i->67	k->10	l->3	m->70	n->6	o->124	p->16	r->5	s->49	t->16	u->7	v->13	ä->19	å->8	
het!	K->1	
het"	 ->3	
het,	 ->116	
het.	 ->4	(->1	A->2	B->1	D->27	E->5	F->8	H->6	I->6	J->12	L->2	M->7	N->6	O->4	P->2	R->2	S->4	T->4	V->10	Å->1	
het:	 ->1	
het;	 ->1	
het?	 ->1	A->1	K->1	N->1	S->1	V->1	
hetJ	a->1	
heta	 ->1	
hete	n->324	r->404	t->1	
hetl	i->36	
hets	 ->2	-->2	a->6	b->3	c->4	e->4	f->26	g->5	k->5	l->3	m->8	n->5	o->4	p->64	r->22	s->9	t->7	u->5	v->2	å->2	
hett	 ->1	a->1	e->1	
heug	e->2	
hez 	t->1	
hhof	e->1	
hiel	 ->1	
hier	a->4	
hies	 ->2	
high	 ->1	
hill	 ->1	
hind	e->34	r->52	
hing	t->3	
hinn	a->2	
hip 	m->1	
hiqu	i->1	
hist	i->2	o->34	
hit 	m->2	o->1	s->1	
hit,	 ->1	
hitt	a->17	i->41	
hjam	o->1	
hjäl	 ->1	p->107	
hjär	t->27	
hler	 ->1	,->1	.->1	s->1	
hne,	 ->1	
hner	 ->3	,->3	s->6	
ho f	ö->1	
ho p	å->1	
ho s	o->1	
ho v	ä->1	
ho. 	D->1	
hobb	y->2	
hoc-	d->1	t->1	
hock	 ->1	a->1	e->2	
hoek	 ->1	
hofe	r->1	
hokl	a->1	
hol,	 ->1	
holk	a->4	
holm	 ->1	,->1	.->1	
hom 	P->3	
homo	f->1	g->2	s->1	
hon 	a->1	f->4	h->4	i->4	j->1	k->2	l->1	p->2	s->4	t->2	u->1	v->1	ä->2	
hono	m->28	
hop 	a->1	d->1	f->1	p->1	s->1	t->1	u->1	ä->1	
hop,	 ->2	
hop.	D->1	I->1	J->1	
hopp	 ->1	a->97	e->1	l->1	n->12	
hord	 ->1	e->1	
hori	s->3	
horm	o->1	
hos 	D->1	E->2	F->1	R->1	a->3	b->2	d->12	e->2	f->3	i->1	k->6	m->4	o->4	p->2	r->1	s->2	t->1	v->2	
hosp	i->1	
hot 	-->1	f->1	m->6	o->1	p->1	s->1	
hota	 ->1	d->6	n->1	r->6	s->4	t->1	
hotb	i->1	
hote	l->1	t->7	
hotf	u->1	
hov 	a->15	i->1	k->1	o->4	s->2	t->8	
hov,	 ->2	
hov.	A->1	H->1	U->1	
hove	n->5	t->34	
hovs	m->5	
how 	t->1	
hren	d->7	
hrey	e->3	
hrko	p->1	
hroe	d->14	
hröd	e->1	
hs i	 ->1	
ht k	a->1	
ht m	e->1	
ht o	c->1	
ht t	i->1	
ht.D	e->1	
htal	a->1	
hter	s->2	
htfö	r->3	
htid	 ->1	
hts.	A->1	
hu o	c->1	
hud 	B->2	
hugg	 ->3	
huld	a->1	
hulz	 ->3	
huma	n->6	
huml	e->1	
humö	r->2	
hun 	s->1	
hund	.->1	r->19	
hur 	E->2	a->5	b->7	d->42	e->3	f->5	g->2	h->4	i->1	k->11	l->9	m->24	n->5	o->2	p->6	r->1	s->26	t->3	u->7	v->31	
hur.	K->1	R->1	
huru	v->14	
hus 	1->1	h->1	o->2	s->1	u->1	
hus,	 ->5	
hus.	E->1	G->1	H->1	
huse	f->3	t->3	
husg	a->4	
hush	å->1	
husl	ä->1	
husö	v->1	
huvu	d->47	
hwar	z->1	
hwei	z->1	
hwit	z->1	
hy o	c->1	
hyck	l->5	
hygi	e->2	
hyll	a->1	n->1	
hypo	t->2	
hyrd	 ->1	
hyre	g->1	
hysa	 ->3	
hyse	r->5	
hyss	e->5	
hyst	e->1	
häft	a->1	i->1	
häle	r->1	
hälf	t->3	
häll	e->42	i->32	s->7	
häls	a->24	n->2	o->8	
hämm	a->4	
hämn	a->1	i->1	
hämt	a->7	n->1	
hän;	 ->1	
händ	a->18	e->61	
hänf	ö->1	
häng	a->6	b->1	e->13	i->2	
häns	e->8	y->72	
hänt	 ->5	.->1	:->1	a->1	
hänv	i->35	
här 	-->6	D->1	a->6	b->9	c->1	d->9	e->3	f->41	g->4	h->6	i->59	k->8	l->5	m->3	n->2	o->14	p->16	r->5	s->18	t->15	u->5	v->11	y->2	ä->8	å->2	ö->2	
här,	 ->14	
här.	 ->1	D->3	E->1	F->1	K->1	V->3	
här;	 ->1	
här?	D->1	
härd	a->2	i->1	l->3	
häre	f->1	
häri	g->2	
härj	a->2	
härl	e->1	
härm	e->3	
härr	ö->4	
härt	i->1	
härv	i->1	
häst	e->1	
häva	 ->3	s->4	
hävd	a->27	v->1	
häve	r->1	
hävs	.->2	
hävt	s->1	
håg 	I->1	a->8	d->3	r->1	s->1	ä->1	
håg.	E->1	
hågo	r->2	
hål 	i->2	
hål,	 ->1	
hål:	 ->1	
håle	n->1	
håll	 ->19	,->5	.->7	:->1	?->1	a->181	b->25	e->121	i->23	n->67	s->22	
hån 	m->1	
håna	r->1	
hård	 ->3	,->1	a->12	n->2	
håre	t->1	
hårk	l->1	
hårt	 ->7	,->1	.->1	
håva	r->1	
hône	-->1	
hög 	a->1	b->1	f->1	g->6	i->1	k->1	n->2	p->2	s->6	
hög,	 ->1	
höga	 ->14	,->1	.->1	k->1	
höge	 ->2	r->30	
högh	e->2	
högl	j->1	
högn	i->3	
högr	a->1	e->19	
högs	k->1	t->28	
högt	 ->9	,->1	.->1	e->2	i->4	
höja	 ->4	n->1	s->1	
höjd	 ->5	e->5	p->2	
höje	r->1	
höjn	i->2	
höjs	 ->1	
höjt	s->1	
höll	 ->14	s->4	
höna	 ->1	
hör 	a->6	b->1	d->2	e->3	f->1	h->6	i->4	j->1	n->3	s->2	t->7	v->2	
hör.	 ->1	
höra	 ->24	,->1	.->2	n->2	r->1	s->2	
hörd	 ->2	.->1	a->1	e->4	
höri	g->19	
hörl	i->1	
hörn	 ->2	s->1	
hört	 ->24	,->1	.->1	s->1	
höst	 ->1	
höva	 ->15	s->1	
hövd	e->2	
höve	r->99	
hövl	i->1	
hövs	 ->20	,->2	.->5	
hövt	 ->2	s->1	
hüss	e->4	
i "g	e->1	
i - 	C->1	a->3	d->1	e->1	j->1	n->1	r->1	s->1	v->1	
i 15	 ->1	
i 19	6->1	9->14	
i 20	 ->1	0->12	
i 55	 ->1	
i 8 	b->1	o->1	
i AB	B->1	
i Ad	a->1	r->1	
i Af	r->3	
i Ak	k->2	
i Al	s->1	
i Am	s->17	
i As	i->1	
i Au	v->1	
i Av	i->1	
i BN	I->1	
i Be	l->2	r->9	
i Bi	s->5	
i Bo	r->1	
i Br	a->2	e->2	y->7	
i Bu	d->1	
i CE	N->1	
i Ca	v->1	
i Ce	n->5	r->1	
i Cu	s->1	
i DD	R->1	
i Da	n->9	
i Du	b->4	
i EC	H->1	
i EG	-->8	
i EK	S->3	
i EM	U->1	
i EU	 ->2	,->1	-->5	:->7	
i Ek	o->1	
i Et	i->1	
i Eu	r->173	
i Fa	c->1	
i Fe	i->1	
i Fi	n->2	
i Fo	l->1	
i Fr	a->11	
i Fö	r->14	
i GU	E->1	
i Ga	z->2	
i Ge	n->2	
i Go	l->2	
i Gr	e->2	u->2	
i Gu	a->1	l->1	
i Ha	i->1	
i He	l->14	
i IC	E->2	
i In	d->1	t->1	
i Ir	l->10	
i Is	r->1	t->1	
i It	a->6	
i Jo	n->1	
i Ka	r->1	u->2	
i Kf	o->1	
i Ki	n->3	
i Ko	s->34	u->1	
i Ky	o->1	
i Kä	r->1	
i Kö	l->1	
i La	m->7	n->4	p->2	
i Le	a->1	
i Li	b->1	i->2	l->1	s->5	
i Lo	m->1	n->4	r->1	
i Lu	t->1	x->4	
i Ma	a->2	c->1	d->2	
i Mc	N->1	
i Me	d->1	l->14	x->1	
i Mi	t->1	
i Mo	n->2	s->1	
i Ne	d->4	w->1	
i No	r->1	
i OL	A->1	
i Om	a->1	
i PP	E->3	
i Pa	d->1	r->1	y->1	
i Pe	k->1	
i Po	r->5	
i Pr	o->1	
i Ra	p->1	
i Ro	m->1	
i Ry	s->2	
i Sa	i->1	n->2	
i Sc	h->4	
i Se	a->3	
i Sh	a->1	e->3	
i Sk	o->2	
i Sr	i->3	
i St	o->11	r->4	
i Sv	e->2	
i Sy	d->2	r->2	
i TV	-->1	
i Ta	d->2	m->14	u->1	
i Te	x->1	
i Th	e->4	y->1	
i Ti	b->5	
i Tu	r->7	
i Ty	s->5	
i UE	N->1	
i US	A->3	
i Ur	b->1	
i Va	n->1	t->1	
i Ve	n->1	
i Vä	r->1	
i Wa	l->3	s->1	
i Wi	e->1	
i Ya	s->1	
i a)	 ->1	
i ab	s->4	
i ac	c->2	
i ag	e->3	
i ai	d->1	
i ak	t->5	
i al	d->1	l->95	
i an	a->3	d->15	l->1	n->5	p->1	s->41	t->1	v->13	
i ar	b->29	t->15	
i at	t->78	
i av	f->1	g->5	h->1	l->1	s->8	t->2	v->6	
i ba	l->1	r->5	
i be	b->1	d->4	f->11	g->4	h->55	k->6	n->1	r->10	s->15	t->24	v->2	
i bi	b->1	d->3	l->12	o->2	
i bl	a->1	e->1	i->5	
i bo	k->1	r->11	
i br	a->1	i->1	o->1	u->2	y->1	ä->1	å->1	
i bu	d->9	
i by	g->1	
i bä	t->2	
i bå	d->3	
i bö	c->1	r->43	
i ce	n->2	
i ci	r->1	
i da	g->166	n->1	t->1	
i de	 ->81	b->10	c->7	l->5	m->4	n->210	r->1	s->28	t->214	
i di	a->2	r->16	s->23	
i do	c->1	k->1	m->4	
i dr	a->1	i->2	
i dä	r->7	
i då	 ->9	
i ef	f->3	t->13	
i eg	e->15	
i ek	o->6	
i em	e->5	
i en	 ->128	a->1	h->1	i->1	k->1	l->28	s->1	
i er	 ->4	a->4	b->1	f->1	k->3	t->7	
i et	t->82	
i eu	r->6	
i ev	e->1	
i ex	a->1	p->2	
i f.	d->1	
i fa	k->6	l->3	r->4	s->4	t->5	
i fe	b->7	m->3	
i fi	c->4	n->3	
i fj	o->2	
i fl	e->7	
i fo	k->1	l->4	r->41	
i fr	a->62	e->8	i->1	o->1	ä->1	å->81	
i fu	l->4	n->2	
i fy	r->2	
i fä	r->3	s->1	
i få	 ->4	r->24	t->5	
i fö	l->3	r->231	
i ga	n->1	r->2	
i ge	 ->4	m->14	n->17	r->7	
i gi	c->1	
i gj	o->6	
i gl	a->2	ä->2	ö->1	
i go	d->13	t->1	
i gr	a->2	u->9	
i gä	l->1	r->2	
i gå	n->6	r->17	
i gö	r->26	
i ha	 ->5	d->11	f->3	m->6	n->16	r->243	v->7	
i he	l->29	m->2	n->1	r->1	
i hi	e->1	s->1	t->5	
i hj	ä->3	
i ho	p->10	
i hu	v->7	
i hy	s->1	
i hä	n->12	r->13	v->2	
i hå	l->10	n->1	r->1	
i hö	g->8	l->1	r->1	s->1	
i i 	E->4	G->2	I->1	L->1	M->1	P->1	S->1	T->1	a->1	d->24	e->5	f->1	g->1	j->1	k->4	m->7	o->1	p->2	s->9	t->1	v->3	Ö->1	å->1	
i ia	k->1	
i ib	l->2	
i ic	k->2	
i ig	e->1	å->1	
i in	b->1	d->1	f->5	g->8	h->1	i->1	k->2	l->11	n->2	o->2	r->2	s->18	t->116	v->1	
i it	a->1	
i ja	g->1	n->1	
i jo	r->1	
i ju	 ->3	l->5	n->6	s->12	
i jä	m->3	
i ka	b->1	l->2	m->21	n->97	p->3	t->1	
i ke	d->1	
i kl	a->8	
i kn	i->1	y->1	
i ko	a->1	m->97	n->27	s->1	
i kr	a->24	i->3	y->1	ä->11	
i ku	l->2	n->9	r->2	
i kv	a->1	ä->4	
i kä	n->13	
i la	d->2	g->13	n->6	
i le	d->3	v->2	
i li	b->1	d->1	k->12	n->5	t->5	v->1	
i lj	u->5	
i lo	v->2	
i ly	c->3	s->3	
i lä	g->8	m->2	n->1	r->1	t->2	
i lå	t->3	
i lö	p->1	s->1	
i ma	j->5	k->1	n->2	r->3	s->1	
i me	d->64	l->2	n->8	r->7	
i mi	g->2	l->6	n->23	s->2	t->18	
i mj	u->1	
i mo	d->1	r->32	t->13	
i my	c->7	n->1	
i mä	n->1	
i må	l->6	n->17	s->145	
i mö	b->1	j->3	
i na	t->7	
i ni	v->4	
i no	r->2	v->5	
i nu	 ->23	l->1	
i ny	a->1	h->1	l->2	
i nä	m->7	r->17	s->1	
i nå	 ->1	g->13	
i nö	d->2	j->1	
i ob	j->1	l->1	
i oc	h->70	k->30	
i of	f->4	t->1	ö->1	
i ok	t->2	
i ol	i->4	j->1	y->1	
i om	 ->6	f->1	r->17	
i on	s->1	
i or	d->7	o->2	
i os	s->10	
i ot	y->1	
i ou	n->1	
i oö	v->1	
i pa	r->40	
i pe	k->1	n->1	r->3	
i pl	a->6	e->4	å->1	ö->1	
i po	l->6	r->2	s->2	
i pr	a->10	e->6	i->12	o->15	
i pu	n->2	
i på	 ->14	b->1	s->1	
i ra	d->2	m->1	p->8	t->2	
i re	a->6	d->11	f->2	g->21	l->2	s->11	t->1	
i ri	k->6	m->1	n->1	s->1	
i ro	p->1	
i ru	l->1	s->2	
i rä	k->4	t->12	
i rå	d->35	
i rö	r->8	s->8	
i sa	d->13	k->2	m->60	t->1	
i se	 ->12	n->2	p->12	r->15	x->1	
i si	d->1	g->19	k->3	n->56	s->2	t->24	
i sj	u->2	ä->28	
i sk	a->74	e->1	i->3	o->2	r->2	u->22	y->3	
i sl	i->2	u->21	ö->1	
i sm	å->2	
i sn	a->11	
i so	c->6	l->1	m->38	r->1	
i sp	e->2	ä->1	
i st	a->5	e->1	i->2	o->12	r->13	y->2	ä->60	å->11	ö->27	
i su	b->1	
i sv	a->3	e->1	å->2	
i sy	d->1	f->8	m->1	n->46	s->5	
i sä	g->9	k->4	m->2	n->1	r->2	t->2	
i så	 ->9	d->7	g->1	l->1	v->1	
i sö	d->1	
i t.	e->2	
i ta	 ->2	c->3	g->3	k->3	l->21	n->2	r->11	
i te	m->1	x->1	
i ti	d->14	l->28	t->1	
i tj	ä->1	
i to	l->3	p->3	r->1	
i tr	a->4	e->5	o->9	ä->2	å->1	
i tv	e->2	i->1	u->3	ä->1	å->5	
i ty	c->7	d->1	s->1	v->2	
i tä	n->6	t->2	
i un	d->13	g->1	i->31	
i up	p->31	
i ur	 ->1	s->1	v->1	
i ut	a->3	b->2	e->1	f->4	g->1	k->1	l->2	n->1	o->1	s->25	t->4	v->11	ö->1	
i va	c->1	d->3	k->1	l->1	n->6	r->37	
i ve	c->1	l->1	m->1	r->18	t->38	
i vi	d->4	k->1	l->85	n->1	s->27	t->13	
i vä	g->3	l->7	n->14	r->12	s->1	
i vå	g->1	r->64	
i yr	k->2	
i yt	t->3	
i zo	n->2	
i ÖV	P->1	
i Ös	t->37	
i äg	a->1	n->4	
i äk	t->1	
i äm	n->3	
i än	 ->1	d->13	n->6	
i är	 ->71	e->1	
i äv	e->6	
i ål	ä->1	
i år	 ->4	,->3	.->4	a->1	t->1	
i ås	t->1	
i åt	a->1	e->7	g->1	m->1	
i ök	a->1	
i ön	s->7	
i öp	p->1	
i ör	e->1	
i ös	t->3	
i öv	e->17	r->5	
i! J	a->1	o->1	
i! U	p->1	
i!He	r->1	
i!Ja	g->1	
i" s	o->1	
i, M	i->1	
i, b	e->1	r->1	
i, d	e->5	å->1	
i, e	f->1	n->3	
i, f	r->3	ö->1	
i, g	i->1	
i, h	e->4	
i, i	n->2	
i, j	a->2	u->1	
i, k	a->2	u->1	
i, l	a->1	i->3	j->1	
i, m	e->9	i->2	
i, n	e->1	ä->1	
i, o	b->1	c->7	m->2	r->1	
i, p	r->1	
i, s	e->1	i->1	k->2	o->5	å->2	
i, t	.->2	i->1	r->1	
i, u	t->2	
i, v	a->1	i->2	
i, ä	n->1	r->1	v->2	
i- o	c->10	
i-, 	t->1	
i-ge	m->1	
i-ir	l->1	
i-ra	s->1	
i.(P	a->1	
i.. 	(->1	
i...	(->1	
i.Al	l->2	
i.An	l->1	
i.Bå	d->1	
i.De	 ->1	n->2	t->8	
i.Dä	r->1	
i.Ef	t->1	
i.En	 ->1	
i.Et	t->1	
i.Eu	r->1	
i.Fo	l->1	r->1	
i.Fr	u->1	
i.Fö	r->1	
i.Ha	i->1	
i.He	r->1	
i.Hu	r->1	
i.Hä	r->1	
i.I 	k->1	
i.Ja	g->3	
i.Ka	n->1	
i.Ku	l->1	
i.Li	k->1	
i.Ma	n->2	
i.Mi	n->1	
i.Nä	r->1	
i.Se	d->1	
i.So	m->1	
i.Så	 ->1	
i.Ut	v->1	
i.Vi	 ->3	d->1	l->1	
i.Vå	r->1	
i: f	r->1	
i; m	a->1	
i? O	c->1	
i?.H	e->1	
ia -	 ->2	
ia B	r->1	
ia E	u->1	
ia P	a->1	
ia R	o->1	
ia a	l->2	t->2	
ia b	i->1	
ia d	a->1	e->2	
ia e	n->1	
ia f	r->1	u->1	
ia h	a->1	
ia i	 ->1	n->1	
ia k	o->1	
ia m	a->1	
ia o	c->2	m->2	
ia r	ö->10	
ia s	a->1	k->1	o->2	t->2	
ia t	i->2	y->1	
ia u	n->1	
ia v	a->3	ä->1	
ia å	t->1	
ia, 	d->1	e->1	o->1	r->1	
ia-R	o->1	
ia.D	e->1	
ia.Ä	n->1	
iage	n->1	
iakt	t->8	
ial 	-->1	b->1	d->2	f->2	i->1	k->1	m->1	n->1	o->6	r->2	s->14	t->4	u->8	
ial,	 ->3	
ial-	 ->1	
ial.	D->2	F->2	J->1	S->1	
iala	 ->78	
ialb	e->2	
iald	e->15	o->1	
iale	n->1	t->3	
ialf	o->17	r->5	ö->6	
iali	n->1	s->41	
ialo	g->31	
ialp	o->4	r->1	
ialt	 ->16	,->1	.->1	
ialu	t->1	
ian 	1->1	
iane	 ->2	,->1	
iano	 ->1	
ians	 ->3	e->4	p->1	
ianv	ä->6	
iari	t->21	
ias 	f->3	o->1	
iasm	 ->3	
iat 	f->1	h->1	
iat.	M->1	
iati	s->4	v->80	
iatä	c->1	
ibak	t->1	
iban	e->1	o->5	
ibbi	g->1	
ibed	r->1	
ibeh	å->11	
ibek	ä->4	
ibel	 ->3	,->1	.->1	t->6	
iber	a->31	i->1	
ibes	p->3	t->2	
ibet	 ->12	"->2	,->3	-->1	.->2	?->1	a->10	
ibi 	n->1	
ibil	i->11	
ibla	 ->3	.->1	n->25	r->2	
ibli	o->2	
ibut	i->1	
ibye	n->1	
ic -	 ->1	
ic B	r->1	
ic i	 ->1	
ical	 ->1	
ican	t->1	
icap	 ->1	
ice 	d->4	f->1	n->1	o->11	t->2	
ice.	A->1	J->1	O->1	S->1	
icek	o->1	v->1	
icen	,->1	s->1	t->1	
icer	a->47	i->10	
icha	r->1	
iche	r->1	
ichi	e->1	
icht	 ->2	.->1	e->2	f->3	
ichy	r->1	
icie	l->7	n->3	
icin	e->1	
icio	 ->1	
icit	.->1	e->2	
ick 	-->1	K->1	a->1	b->3	d->3	e->5	f->2	h->2	i->6	j->5	k->1	m->4	n->3	o->4	s->3	t->3	u->1	v->4	
ick,	 ->3	
ick.	A->1	D->1	H->1	K->1	Ä->1	
icka	 ->6	,->1	d->2	r->3	s->1	t->2	
ickb	a->5	
icke	 ->15	-->19	n->1	r->2	t->11	
ickf	r->1	
ickl	i->1	
ickn	i->1	
icko	r->2	
ickp	r->3	
icks	.->1	i->3	v->1	
icy,	 ->1	
icya	v->1	
icyd	e->1	
icyf	ö->1	
id 1	2->1	
id 7	0->1	
id B	y->3	
id E	G->3	U->1	u->4	
id G	e->1	
id H	a->1	
id K	y->1	
id L	a->1	
id M	e->1	
id P	a->1	
id a	)->1	l->3	n->8	r->1	t->27	v->3	
id b	a->1	e->9	l->2	r->1	ä->1	ö->5	
id c	a->1	
id d	a->1	e->41	o->2	r->1	ä->1	å->3	
id e	f->2	l->1	n->10	t->12	v->1	
id f	a->2	i->2	l->6	r->5	u->1	y->1	å->2	ö->20	
id g	j->2	o->1	r->2	ö->1	
id h	a->15	e->1	i->1	j->1	ä->1	ö->3	
id i	 ->7	n->10	
id j	a->1	o->1	ä->1	
id k	a->5	l->1	o->6	r->2	u->2	ä->1	
id l	a->1	i->1	u->1	ä->2	
id m	a->1	e->9	i->3	o->2	y->1	ä->1	å->2	ö->3	
id n	a->3	o->1	u->1	y->1	ä->2	å->2	
id o	c->7	e->1	f->1	m->7	p->1	r->1	
id p	a->2	l->2	r->3	u->2	å->4	
id r	e->4	ä->2	å->1	
id s	a->3	e->1	i->8	j->2	k->5	l->2	o->4	t->6	y->1	ä->2	å->2	
id t	a->3	e->1	i->8	o->2	r->4	v->2	
id u	n->2	p->3	t->11	
id v	a->6	i->7	å->1	
id y	r->1	
id ä	n->2	r->8	v->1	
id å	r->2	t->3	
id ö	v->2	
id, 	a->2	d->1	e->1	f->1	h->2	i->2	m->1	o->4	p->1	v->3	ä->1	
id..	 ->1	
id.D	e->5	
id.E	n->1	
id.F	ö->1	
id.H	a->1	
id.J	a->1	
id.K	o->1	
id.M	a->1	
id.N	ä->1	
id.O	m->1	
id.S	o->1	
id.T	a->1	i->1	
id.V	i->1	
id: 	d->1	
ida 	E->1	G->1	a->2	b->4	d->11	e->2	f->5	g->1	h->1	i->7	k->5	m->3	n->2	o->2	p->1	r->1	s->6	t->4	u->1	v->3	å->1	
ida,	 ->9	
ida.	D->1	F->1	H->1	I->1	J->1	O->1	V->1	Ä->1	
ida?	I->1	
idag	,->1	
idak	i->2	
idan	 ->43	,->2	.->1	d->15	
idar	e->44	i->31	
idas	 ->1	
idat	 ->1	e->1	l->12	
idd 	b->1	h->1	m->1	o->1	ä->1	
idd.	J->1	
idda	g->13	
idde	l->1	n->1	
ide 	W->1	
idea	l->5	
idee	l->2	
idem	o->1	
iden	 ->76	,->7	.->31	:->1	?->2	s->3	t->30	
ideo	l->5	
ider	 ->48	,->5	.->5	a->8	i->13	s->19	
ides	 ->2	
idga	 ->14	?->1	d->5	r->3	s->13	t->2	
idgn	i->71	
idhå	l->4	
idhö	l->1	
idia	r->21	
idig	 ->7	a->84	h->1	t->78	
idis	k->31	
idit	 ->3	s->1	
idiä	r->1	
idka	r->1	
idla	g->1	n->1	
idli	g->5	
idma	k->1	
idna	p->1	
idni	n->22	
idoe	f->1	
idor	 ->3	.->1	e->2	n->2	
idos	k->2	
idpu	n->10	
idra	 ->35	,->1	g->52	r->20	
idro	g->3	t->4	
ids 	i->1	m->1	p->1	t->1	u->1	ä->1	
ids,	 ->1	
ids-	s->1	
idsa	r->4	
idsb	e->2	
idsd	i->3	u->1	
idsf	r->10	ö->1	
idsg	r->1	
idsi	n->2	
idsm	ä->2	
idso	r->1	
idsp	a->2	e->10	l->5	
idsr	a->5	y->2	
idss	k->1	y->1	
idst	r->1	
idså	l->2	t->1	
idsö	d->1	
idta	 ->33	b->6	g->6	l->1	r->8	s->14	
idto	g->2	
idua	l->1	
idue	l->7	r->1	
idut	s->1	
idé 	-->1	a->2	j->1	k->1	o->1	s->3	ä->1	
idé,	 ->1	
idée	r->8	
idén	 ->13	,->1	
ie C	u->1	
ie R	e->1	
ie a	v->1	
ie o	c->1	
ie, 	h->1	
ie- 	o->1	
ie-s	t->1	
iebe	n->1	s->1	
iebö	r->1	
ieck	 ->1	
ied 	(->1	
ied.	K->1	
iede	p->2	
ieff	e->6	
iefi	n->1	
iefu	s->1	
iekt	i->1	
iel 	v->1	
iela	n->4	
ielf	t->1	
iell	 ->15	,->1	a->61	t->42	
iels	e->7	o->5	
iemi	n->3	
ien 	9->1	a->3	b->1	d->1	e->3	f->3	h->9	i->3	j->1	m->1	n->1	o->21	s->9	t->3	ä->6	
ien,	 ->23	
ien.	D->2	E->1	F->1	H->1	I->1	M->1	O->1	P->1	S->2	U->1	V->1	
ien?	E->1	V->1	
iend	e->1	
ienf	r->1	
ienn	e->1	
iens	 ->10	e->2	k->17	
ient	 ->1	e->10	i->2	l->33	
iepr	o->1	
ier 	-->6	D->1	a->3	e->2	f->13	g->1	h->3	i->1	k->4	m->4	o->21	p->2	r->3	s->17	t->1	u->2	ä->1	ö->1	
ier,	 ->16	
ier.	.->1	A->1	D->4	K->2	L->1	M->2	
iera	 ->16	d->16	r->7	s->11	t->12	
ierb	a->2	
ierd	o->1	
ieri	n->43	
iern	a->44	
iers	 ->2	
ies 	a->1	r->1	v->1	
iesk	i->2	
iesm	i->1	
iest	r->1	
iet 	(->3	D->1	I->1	a->2	d->1	e->2	f->1	h->7	i->3	m->1	n->2	o->7	p->1	r->1	s->4	t->1	v->1	ä->3	
iet"	.->1	
iet)	 ->1	,->2	.->1	
iet,	 ->9	
iet.	A->1	D->2	H->1	M->1	O->1	V->3	
ietn	i->3	
iets	 ->22	
iety	 ->1	
ieur	o->1	
ieäg	a->2	
ifal	l->5	
ifar	t->2	
ifas	c->3	
ifer	a->4	i->1	t->1	
ifes	t->1	
iffe	r->5	
iffr	a->7	o->15	
ific	e->38	i->2	
ifie	r->27	
ifik	 ->3	a->22	t->7	
ifin	-->1	a->1	
ifiq	u->1	
ifol	k->1	
ifon	d->2	
ifor	m->1	
ifrå	g->26	n->35	
ift 	a->3	d->1	e->1	f->3	i->2	k->1	m->1	o->2	p->1	r->1	s->5	t->1	v->1	ä->3	
ift!	H->1	
ift,	 ->2	
ift.	 ->1	A->1	D->1	E->1	J->1	O->1	V->1	
ift:	 ->1	
ifta	 ->4	n->5	r->6	t->1	
ifte	 ->1	,->1	.->1	n->8	r->64	t->3	
ifti	g->3	
iftl	i->8	
iftn	i->113	
ifts	-->1	f->2	l->2	m->1	p->2	s->1	t->1	ä->1	
iful	l->1	
iför	b->1	r->1	s->2	
ig -	 ->1	,->1	
ig E	u->1	
ig O	L->1	
ig a	c->1	l->5	n->10	r->4	s->2	t->63	v->15	
ig b	a->10	e->14	i->1	l->2	o->1	r->3	y->2	ä->2	ö->1	
ig d	a->1	e->35	i->4	j->1	o->2	ä->3	ö->2	
ig e	f->4	k->1	l->5	m->4	n->11	r->1	t->6	u->1	x->2	
ig f	a->1	i->1	o->1	r->29	u->4	å->2	ö->86	
ig g	a->1	e->2	i->2	l->1	r->10	ä->2	ö->2	
ig h	a->10	e->3	i->2	j->3	u->3	ä->5	
ig i	 ->40	.->1	h->1	n->36	v->1	
ig j	o->1	u->3	ä->1	
ig k	a->7	l->1	n->1	o->20	r->1	u->3	v->1	ä->1	
ig l	a->4	e->3	i->1	ä->3	ö->5	
ig m	a->10	e->26	i->4	o->8	y->10	ä->1	å->4	ö->2	
ig n	a->2	e->3	i->3	o->2	u->1	y->1	ä->7	å->1	ö->1	
ig o	b->2	c->53	e->1	f->2	m->40	n->2	r->2	
ig p	a->1	e->4	o->7	r->4	u->7	å->37	
ig r	a->3	e->15	i->3	o->8	u->1	y->1	ä->2	å->2	
ig s	a->8	e->6	i->8	j->11	k->5	l->2	o->11	t->10	u->1	v->1	y->2	ä->9	å->2	
ig t	.->1	a->2	e->2	i->50	o->1	r->1	v->2	y->1	
ig u	n->5	p->7	t->27	
ig v	a->18	e->1	i->6	ä->4	
ig y	r->1	t->1	
ig ä	n->3	r->9	v->2	
ig å	 ->1	k->1	s->3	t->20	
ig ö	k->1	v->9	
ig!"	.->1	
ig!H	a->1	
ig".	E->1	
ig, 	a->4	b->2	d->3	e->4	f->2	g->2	h->5	i->1	l->1	m->4	n->4	o->5	p->1	s->8	u->1	v->3	
ig. 	F->1	S->1	
ig.A	v->1	
ig.B	r->1	
ig.D	e->10	
ig.E	m->1	n->1	r->1	u->1	
ig.G	e->1	r->1	
ig.H	e->2	
ig.I	 ->1	
ig.J	a->13	
ig.K	o->1	
ig.M	a->2	e->2	
ig.N	a->1	
ig.O	c->3	
ig.P	r->1	
ig.S	a->1	
ig.T	a->1	
ig.U	n->1	
ig.V	a->1	i->4	
ig.Ä	r->1	
ig: 	d->2	h->1	
ig; 	d->1	
ig?D	e->1	
ig?H	u->1	
ig?J	o->1	
ig?V	a->1	
iga 	"->1	-->5	3->1	E->4	H->1	a->34	b->55	c->1	d->23	e->20	f->138	g->22	h->14	i->43	k->41	l->25	m->47	n->9	o->85	p->37	r->78	s->111	t->24	u->18	v->22	y->1	ä->22	å->13	ö->9	
iga,	 ->34	
iga.	 ->1	(->1	A->3	D->3	E->1	F->3	H->2	I->4	J->1	M->2	N->2	O->1	P->2	S->1	V->4	
iga/	h->1	
iga;	 ->1	
iga?	F->1	
igad	,->1	.->2	e->8	
igan	d->11	t->5	
igar	 ->4	e->166	
igas	 ->4	,->2	t->52	
igat	 ->8	,->2	.->1	o->14	s->2	
igdo	m->12	
ige 	i->1	o->3	p->1	s->1	
ige.	 ->1	J->1	
igen	 ->482	"->1	,->27	.->12	:->2	a->3	k->1	o->37	s->2	t->4	
iger	 ->2	.->1	a->1	n->1	
iges	 ->1	
iget	 ->5	.->3	s->4	
igga	 ->13	n->10	
igge	r->87	
iggj	o->13	
iggö	r->21	
igh 	l->1	
ighe	t->830	
ight	 ->2	s->1	
ighå	l->2	
igie	r->1	
igin	a->1	e->1	
igit	 ->1	.->1	
igiö	s->4	
igjo	r->1	
igla	n->1	
igli	g->4	
igma	t->1	
igna	 ->1	l->14	
igne	l->1	r->1	
igno	r->4	
igor	ö->4	
igot	t->1	
igou	 ->1	
igra	 ->2	n->2	t->8	
igre	r->1	
igse	k->1	
igsh	e->1	
igss	k->1	
igst	ä->1	
igt 	-->6	:->1	D->1	E->2	G->1	I->1	K->1	R->1	S->1	T->1	a->226	b->29	d->30	e->34	f->94	g->47	h->31	i->41	j->2	k->28	l->15	m->89	n->14	o->80	p->35	r->13	s->137	t->31	u->22	v->45	y->2	ä->16	å->3	ö->5	
igt!	L->1	M->1	
igt,	 ->62	
igt.	A->1	D->11	E->3	F->8	G->2	H->5	I->1	J->11	L->2	M->9	N->2	O->3	P->1	S->3	U->1	V->13	Ö->1	
igt:	 ->1	
igt;	 ->1	
igt?	A->1	
igtv	i->108	
igva	t->1	
igå 	d->1	
igåe	n->4	
igån	g->7	
igås	 ->1	
igör	 ->1	a->4	s->1	
ihan	;->1	d->2	
ihet	 ->44	,->38	.->5	:->1	;->1	e->25	s->2	
ihjä	l->1	
ihop	 ->8	,->1	.->3	
ihär	d->1	
ihåg	 ->15	.->1	
iika	n->3	
iimp	o->1	
iinn	e->1	
iint	r->1	
iis-	J->2	
ij-v	a->1	
ijs 	o->1	
ijs.	(->1	
ik -	 ->2	
ik D	e->1	
ik J	ö->1	
ik a	n->1	v->4	
ik e	g->1	l->2	n->1	t->1	
ik f	i->1	r->1	å->1	ö->16	
ik h	a->3	u->1	ö->1	
ik i	 ->9	n->2	
ik k	a->2	u->1	
ik m	e->5	i->1	o->3	å->3	ö->1	
ik n	ä->3	
ik o	c->28	m->2	r->1	
ik p	o->2	å->3	
ik r	e->1	ö->1	
ik s	a->1	k->1	o->31	t->1	å->1	
ik t	i->1	
ik u	n->1	p->1	t->1	
ik v	a->1	i->2	
ik ä	r->5	
ik å	t->1	
ik ö	v->1	
ik!O	m->1	
ik" 	o->1	
ik, 	d->6	e->2	f->2	h->1	i->2	m->1	n->3	o->1	s->3	t->10	u->1	v->3	
ik- 	o->2	
ik..	(->1	
ik.B	y->1	
ik.D	e->9	ä->1	å->1	
ik.E	n->1	u->1	
ik.F	a->1	r->2	ö->1	
ik.G	e->1	
ik.H	a->2	i->1	ä->1	
ik.I	 ->1	
ik.J	a->1	
ik.M	e->1	
ik.R	e->1	i->1	
ik.T	v->1	
ik.V	i->3	
ik.Ä	v->1	
ik: 	v->1	
ik?H	e->1	
ik?V	a->1	
ika 	E->1	a->11	b->15	d->13	e->8	f->23	g->9	h->6	i->13	k->10	l->10	m->18	n->10	o->6	p->13	r->15	s->22	t->9	u->7	v->17	ä->8	å->4	ö->3	
ika,	 ->9	
ika-	o->1	
ika.	D->1	I->1	J->3	P->1	V->2	
ikab	e->2	
ikad	a->2	
ikaf	r->1	
ikal	 ->3	a->9	e->1	i->6	t->5	y->1	
ikan	 ->1	d->6	e->13	s->11	
ikap	a->1	i->1	p->5	r->1	
ikar	 ->4	e->4	n->5	t->2	
ikas	 ->10	.->2	m->1	t->3	å->4	
ikat	 ->6	,->1	i->18	o->5	
ike 	(->1	-->3	a->3	b->3	d->1	e->4	f->2	g->2	h->2	i->4	k->3	m->4	n->1	o->10	s->7	t->1	v->2	ä->3	
ike,	 ->15	
ike.	 ->1	.->2	D->5	F->3	I->1	J->2	M->1	N->1	O->1	V->3	Ö->1	
ike:	 ->1	
ikeE	n->1	
ikeF	r->1	
ikeN	ä->1	
iked	o->10	
ikel	 ->93	,->2	s->5	
iken	 ->97	,->21	.->28	?->2	H->1	s->19	
iker	 ->25	,->4	.->1	n->12	s->1	
ikes	 ->26	-->4	f->4	h->4	m->9	p->3	
iket	 ->7	,->3	.->2	s->6	
ikgi	l->2	
ikh 	h->1	
ikh-	a->1	
ikh.	D->1	F->1	
ikhe	t->35	
ikis	k->49	t->5	
ikit	 ->1	i->2	
ikla	r->15	
ikle	d->1	
ikli	g->6	
ikme	t->2	
ikna	.->1	n->19	r->2	
ikni	n->44	
iko,	 ->1	
ikol	o->1	
ikom	m->1	r->6	
ikon	t->2	v->1	
ikra	f->4	t->1	v->2	
ikri	k->4	
ikro	f->1	k->2	s->1	
ikry	p->2	
iks 	m->1	
ikso	m->55	
ikst	ä->2	
ikt 	-->2	F->1	a->25	b->4	d->3	e->4	f->5	g->2	h->5	i->4	k->9	l->4	m->5	o->13	p->2	r->1	s->14	v->10	ä->9	ö->1	
ikt,	 ->13	
ikt.	B->1	D->3	I->1	J->1	K->1	O->3	R->1	V->1	
ikt;	 ->1	
ikta	 ->19	,->1	.->1	d->19	n->1	r->9	s->3	t->16	
ikte	,->2	.->1	l->13	n->44	r->31	
iktf	ö->1	
ikti	g->454	o->9	v->1	
iktl	i->78	
iktn	i->55	
iktp	u->2	
ikts	f->3	m->1	p->1	
ikvä	l->4	r->5	
ikäl	l->37	
il -	 ->1	,->1	
il 1	9->1	
il P	o->1	
il e	l->3	n->1	
il f	ö->2	
il g	r->2	
il i	 ->1	
il k	o->1	
il m	e->2	
il n	ä->1	
il o	c->1	
il s	o->5	ä->2	
il u	t->2	
il v	e->1	
il, 	s->1	t->1	
il- 	o->2	
il-D	e->1	
il-R	o->1	
il-p	r->1	
il. 	E->1	
il.D	e->2	
il.J	a->1	
il.L	y->1	
il.T	r->1	
ila 	b->3	s->3	
ilag	a->4	o->2	s->1	
ilan	k->1	
ilar	 ->45	,->14	.->13	?->1	b->1	e->1	n->10	
ilat	e->9	
ilbe	f->2	s->1	
ilbr	a->1	
ild 	a->2	b->3	f->2	i->1	k->3	m->2	o->1	p->1	r->2	t->2	u->2	
ild,	 ->1	
ild.	D->1	F->1	N->1	
ilda	 ->42	d->3	n->5	r->6	s->8	t->3	
ilde	 ->2	,->1	.->1	l->3	n->2	r->2	
ildn	i->66	
ildr	a->6	
iled	a->1	
ileg	e->2	i->4	
ilem	m->3	
ilen	 ->3	,->2	.->2	
iler	a->1	
ilfö	r->2	
ilhe	l->1	
ilia	-->1	
ilie	n->1	
ilig	i->1	
ilik	n->1	
ilin	d->30	
ilis	 ->1	a->1	e->11	m->1	t->1	
ilit	a->2	e->27	ä->6	
ilj 	L->1	
ilja	 ->185	,->2	.->2	d->3	k->4	n->19	r->21	s->9	t->8	
ilje	-->1	d->1	f->2	j->3	l->1	m->1	r->15	s->1	å->1	
iljo	n->65	
iljt	 ->1	
iljö	 ->8	!->1	,->11	-->2	.->6	a->4	b->4	d->2	e->4	f->10	i->1	k->26	l->1	m->15	n->39	o->5	p->14	r->3	s->24	u->1	v->9	
ilka	 ->104	s->2	
ilke	n->55	t->180	
ilko	n->1	
ilky	r->1	
ilkö	p->2	
ill 	"->1	-->2	1->5	2->4	3->2	4->1	5->1	7->3	8->2	9->4	A->1	B->5	C->2	D->1	E->32	F->7	G->2	I->1	K->13	L->2	M->4	N->2	O->1	P->5	R->1	S->7	T->5	V->1	W->4	a->333	b->75	c->1	d->293	e->203	f->165	g->59	h->72	i->41	j->103	k->73	l->19	m->80	n->43	o->77	p->40	r->57	s->214	t->62	u->37	v->92	y->5	Ö->1	ä->21	å->12	ö->5	
ill!	H->1	
ill,	 ->25	
ill.	A->1	D->5	E->1	F->1	H->2	I->2	J->1	R->1	S->1	V->1	
ill:	 ->1	
ill?	D->1	H->1	J->1	
illa	 ->9	,->2	r->1	v->1	
illb	a->52	r->4	
illd	e->12	r->1	
ille	 ->12	g->8	n->7	r->3	s->1	
illf	i->1	o->6	r->27	ä->97	ö->13	
illg	o->1	r->2	ä->21	å->25	
illh	a->43	e->2	ö->8	
illi	!->1	g->27	n->1	
illk	o->70	ä->9	
illm	ä->2	ö->3	
illn	a->44	i->1	ä->6	
illo	b->2	j->2	l->1	r->1	
illr	ä->77	
ills	 ->42	,->2	.->3	?->1	a->33	e->13	k->5	l->1	t->22	v->3	ä->4	
illt	a->3	r->8	
illv	a->1	e->86	i->2	ä->29	
illä	g->20	m->177	
illå	t->55	
ilme	n->1	r->1	
ilmä	r->1	
ilo 	g->1	m->1	o->1	
ilo,	 ->1	
ilob	b->1	
ilom	e->1	
ilos	o->5	
ilot	 ->1	e->1	p->2	
ilov	o->1	
ilpa	r->6	
ilpr	o->1	
ilre	g->1	
ilrä	t->1	
ils 	l->2	
ilse	 ->1	k->1	l->2	
ilsk	a->3	r->2	y->2	ö->1	
ilsp	r->1	
ilst	o->1	
ilt 	E->2	S->2	a->3	b->9	d->7	e->3	f->14	g->5	h->3	i->11	j->2	k->3	l->1	m->11	n->5	o->2	p->8	s->6	t->12	u->4	v->17	ä->2	å->1	
ilt,	 ->1	
ilti	b->1	g->26	l->17	
ilto	n->1	
iltr	e->1	
ilur	e->1	
ilve	r->3	
ilvr	a->6	
iläg	a->1	
ilän	g->1	
ilåt	e->1	
ilön	e->1	
ima 	f->1	i->1	o->2	s->1	
ima,	 ->1	
ima.	H->1	
imag	e->1	i->1	
imal	 ->3	a->4	i->1	t->3	
iman	g->3	
imat	 ->1	.->1	e->7	f->4	p->1	u->1	
imbu	s->1	
imen	 ->1	.->1	s->14	t->1	
imer	a->8	i->1	
imet	e->1	
imib	e->2	
imif	i->1	
imii	n->1	
imik	a->1	o->1	r->2	
imil	ä->1	ö->1	
imin	a->4	e->26	i->1	o->2	ä->3	
imir	e->5	
imis	-->1	t->6	
imit	e->6	i->1	r->5	
imix	e->1	
imiå	l->1	
imli	g->23	
imma	 ->1	r->7	t->1	
imme	 ->5	
immi	g->6	
immu	n->1	
imor	u->1	
impl	e->1	
impo	n->3	p->1	r->6	
imps	o->1	
impu	l->6	
imsa	v->2	
imsb	e->2	
imso	l->1	
imsp	a->1	
imsr	å->2	
imså	t->1	
imt 	i->1	o->2	
imt,	 ->1	
imul	a->6	e->7	
imum	 ->4	
imus	-->1	
imyn	d->1	
imål	,->1	
imög	e->1	
in -	 ->1	
in 1	9->1	
in 2	6->1	
in E	u->1	
in F	r->1	
in a	b->1	k->1	n->7	r->2	t->4	v->4	
in b	a->1	e->9	i->6	l->1	r->2	u->2	
in d	a->2	e->13	j->2	o->1	r->1	
in e	g->10	k->3	n->3	r->2	t->2	x->2	
in f	a->1	o->1	r->19	u->1	y->1	å->1	ö->21	
in g	e->1	l->2	o->1	r->30	
in h	a->6	e->12	u->1	ä->2	ö->2	
in i	 ->33	,->1	n->6	
in k	a->3	o->32	r->1	ä->1	
in l	i->4	ö->1	
in m	a->4	e->20	o->3	å->3	
in n	a->5	u->2	y->1	ä->2	
in o	b->1	c->34	r->6	s->1	
in p	a->1	e->4	l->4	o->4	r->2	å->25	
in r	a->2	e->6	i->2	o->6	ä->5	ö->6	
in s	e->1	i->7	j->2	k->4	l->2	o->18	p->3	t->8	u->1	y->2	ä->2	å->3	
in t	i->4	r->3	u->6	
in u	n->4	p->19	t->7	
in v	a->4	e->1	i->4	u->1	ä->2	å->2	
in w	e->1	
in y	t->1	
in ä	n->1	r->2	
in å	s->12	
in ö	n->4	
in!H	e->1	
in",	 ->1	
in, 	d->1	e->1	f->3	g->2	h->2	m->3	o->7	p->2	r->1	s->5	t->1	u->1	v->2	
in-r	å->3	
in. 	D->1	M->1	
in.A	l->1	
in.B	e->1	
in.C	e->1	
in.D	e->5	ä->1	
in.F	ö->2	
in.H	e->2	
in.I	n->1	
in.J	a->3	
in.L	i->1	å->1	
in.M	e->1	
in.N	ä->1	
in.O	m->2	
in.S	a->1	c->1	t->1	
in.V	a->1	i->4	
in: 	e->1	
in?P	a->1	
ina 	a->10	b->8	d->40	e->18	f->18	g->9	h->7	i->9	j->1	k->29	l->5	m->8	n->3	o->9	p->1	r->16	s->19	t->9	u->10	v->7	y->1	ä->3	å->3	ö->3	
ina,	 ->1	
ina-	I->1	
ina.	H->1	U->1	
inaf	l->1	r->1	
inal	 ->1	e->3	i->5	p->1	v->1	
inan	s->84	
inar	b->1	i->1	
inas	 ->2	
inat	i->8	
inav	i->1	
inba	n->1	
inbe	g->12	
inbj	u->6	ö->1	
inbl	a->14	
inbu	r->1	
inby	g->1	
inci	d->1	p->194	t->8	
ind 	o->1	
inda	 ->3	.->2	n->12	
inde	 ->1	l->18	n->1	r->42	
indf	ä->4	
indi	k->6	r->7	s->1	v->14	
indr	a->53	e->56	ä->2	
indu	s->113	
ine 	d->1	f->1	h->1	n->1	q->2	
ine,	 ->1	
inef	f->3	
inel	l->4	
inen	 ->4	,->3	s->2	t->5	
iner	 ->8	a->17	i->31	n->1	
ines	e->2	i->7	
inet	t->3	
inez	 ->1	
infe	k->2	
infi	l->1	n->2	
infl	y->12	
info	r->92	
infr	a->15	i->1	å->1	
infö	r->164	
ing 	(->6	-->11	1->2	2->2	3->1	6->2	8->2	D->1	E->2	F->1	I->2	T->1	V->1	a->359	b->14	d->12	e->22	f->111	g->10	h->22	i->116	k->23	l->8	m->70	n->10	o->173	p->53	r->6	s->135	t->52	u->12	v->25	ä->40	å->4	ö->2	
ing!	J->1	
ing"	 ->2	,->2	.->1	
ing)	 ->4	.->1	N->1	
ing,	 ->196	
ing-	P->1	
ing.	 ->4	(->1	.->2	A->8	D->65	E->7	F->15	G->2	H->14	I->14	J->29	K->9	L->3	M->13	N->7	O->13	P->5	R->1	S->7	T->3	V->17	Ä->2	
ing:	 ->3	D->1	
ing;	 ->4	
ing?	D->2	H->1	J->1	O->1	T->1	Ä->1	
inga	 ->40	.->1	d->6	l->3	n->8	r->572	s->11	t->4	
ingd	y->1	
inge	l->1	n->901	r->3	t->33	
ingf	l->1	o->21	
ingg	å->2	
ingi	v->6	
ingo	m->4	
ingp	o->2	
ingr	a->2	e->8	i->10	
ings	 ->5	-->12	a->22	b->23	c->13	d->4	e->3	f->320	g->6	h->2	i->11	k->190	l->71	m->27	n->7	o->12	p->94	r->22	s->72	t->14	u->7	v->45	ä->1	å->6	ö->1	
ingt	o->5	v->4	
ingå	 ->8	.->1	e->5	n->1	r->13	t->6	
inhe	m->2	
inho	 ->4	.->1	s->1	
inhä	m->6	
inie	r->17	
inif	r->1	
inim	a->1	e->1	i->19	o->1	u->5	
inin	g->1	
inio	n->4	
inip	e->1	
inir	e->1	
inis	t->99	
init	i->102	u->1	
iniv	å->1	
inje	 ->11	.->2	n->3	r->77	
inke	l->11	
inkl	a->1	u->21	
inko	m->13	n->3	
inkr	i->1	ä->1	
inkt	e->1	i->2	
inkö	p->2	r->1	
inla	n->6	
inle	d->60	t->13	
inli	g->1	
inlä	g->18	m->5	n->5	
inlå	s->1	t->1	
inlö	p->1	
inmä	s->1	
inna	 ->63	,->1	.->1	n->39	s->50	t->1	
inne	 ->9	,->5	.->1	b->116	f->6	h->84	l->1	n->3	r->69	s->3	t->2	v->2	
inni	g->1	n->49	
innl	i->2	
inno	c->24	p->2	r->59	v->6	
inns	 ->321	,->3	.->6	
ino 	i->1	k->1	o->1	
ino,	 ->2	
ino.	J->1	O->1	
inom	 ->283	e->1	
inor	i->22	m->2	n->1	
inos	 ->3	,->2	
inot	t->1	
inpr	ä->1	
inra	 ->11	r->1	s->1	
inre	 ->82	s->4	
inri	k->57	
inry	m->1	
inrä	t->55	
inrå	d->1	
ins 	a->4	d->1	f->1	i->2	j->1	k->2	l->1	p->1	r->1	s->4	t->1	v->1	å->1	
insa	m->8	t->41	
insb	u->1	
inse	 ->13	;->1	e->1	m->3	r->25	
insi	k->4	s->6	
insk	 ->2	a->61	n->16	r->13	
insl	a->6	
insp	e->12	i->3	
inst	 ->28	,->1	a->37	e->8	i->138	m->1	o->27	r->61	s->1	ä->48	
insy	n->13	
int 	b->1	
int-	E->1	
inta	 ->4	g->5	r->4	
inte	 ->1566	!->2	,->13	.->14	:->1	?->2	g->42	l->13	n->13	r->109	t->2	
inti	m->1	
intl	i->10	
into	g->2	l->4	n->1	
intr	e->120	o->6	y->15	ä->28	å->1	
inty	g->4	
intä	k->5	
inuc	 ->1	
inue	r->2	
inus	 ->3	g->2	
inut	 ->3	.->3	e->10	
inva	l->1	n->18	
inve	c->2	n->1	r->7	s->15	
invi	t->1	
invo	l->9	
invä	n->13	
invå	n->9	
inz 	F->2	
inär	 ->1	a->8	e->1	f->1	p->1	
inöv	a->1	
io S	á->1	
io V	a->3	i->1	
io b	e->2	
io f	a->1	ö->3	
io g	r->1	å->2	
io h	a->1	
io l	ä->1	
io m	i->7	å->2	
io p	u->1	
io s	a->1	i->1	k->1	å->1	
io t	i->1	
io u	t->1	
io ä	n->1	
io å	r->7	
io, 	a->1	s->1	t->1	
io-P	l->4	
io.J	a->1	
io.N	ä->1	
io: 	v->1	
io; 	d->1	
iod 	a->2	d->2	f->4	i->4	k->1	o->1	p->2	r->2	s->2	v->1	ä->2	
iod,	 ->5	
iod.	D->1	V->1	
iod?	-->1	
iode	n->39	r->2	
iodi	s->14	
ioek	o->3	
ioel	v->1	
iofe	m->1	
iofö	r->1	
iogr	a->1	
iola	 ->1	
iolo	g->6	
ion 	(->5	-->3	1->5	5->1	A->1	H->1	I->1	P->2	a->25	b->5	d->8	e->4	f->24	g->5	h->8	i->29	j->1	k->9	m->15	n->3	o->53	p->9	r->1	s->64	t->20	u->6	v->7	ä->6	å->2	
ion"	 ->1	
ion)	 ->2	
ion,	 ->48	
ion.	 ->3	1->1	B->1	D->18	E->2	F->5	G->1	H->5	I->6	J->10	K->2	M->3	N->1	O->2	S->5	T->2	U->1	V->11	Å->1	
ion:	 ->3	
ion;	 ->1	
ion?	 ->1	D->1	J->1	K->2	Ä->1	
iona	l->135	
iond	e->2	
ione	l->275	n->1502	r->476	
ioni	s->5	
ionj	ä->1	
ions	 ->2	-->4	a->12	b->2	d->3	f->23	h->9	i->1	k->14	l->12	m->7	n->2	o->1	p->11	r->16	s->17	t->3	u->7	v->1	ä->1	
ionä	r->248	
iopi	e->3	
iopl	a->1	
ior.	D->1	
iorg	a->2	
iori	 ->3	t->36	
ios 	i->1	å->1	
iosf	ä->1	
iosj	u->1	
iosä	k->2	
iot 	i->1	s->1	
iota	l->6	
iote	k->2	
ioti	s->1	
iotu	s->1	
ioxi	d->5	n->2	
ip a	l->1	t->2	
ip e	l->1	n->2	
ip f	ö->1	
ip i	 ->2	n->5	
ip m	e->1	
ip o	c->2	m->2	
ip r	å->1	
ip s	o->4	å->1	
ip ä	r->3	v->1	
ip, 	g->1	m->1	o->1	
ip.J	a->1	
ip.S	j->1	
ip.V	i->2	
ipa 	a->1	d->3	e->2	i->3	m->1	o->2	p->1	r->2	t->2	
ipa,	 ->1	
ipa.	E->1	K->1	
ipan	d->20	
ipar	a->1	
ipas	 ->1	
ipen	 ->73	,->11	.->17	:->2	N->1	d->1	
iper	 ->43	,->4	.->5	:->1	n->10	
ipes	 ->1	
ipet	 ->2	,->1	
ipie	l->8	
ipit	 ->2	
ipla	n->1	
ipli	g->6	n->14	
iplo	m->11	
ipna	 ->1	
ipni	n->9	
ipol	i->4	
ipot	e->1	
ippa	d->3	
ippe	r->2	
ipro	d->3	g->4	
ips 	a->1	
ipsk	ä->1	
ique	 ->1	s->2	
iqui	t->1	
ir E	u->2	
ir a	l->3	n->2	t->4	v->1	
ir b	i->1	r->1	ä->1	
ir d	e->12	i->2	
ir e	n->7	t->3	
ir f	o->1	r->2	ö->3	
ir g	r->1	
ir h	a->1	j->1	o->1	
ir i	 ->2	n->3	
ir j	a->1	u->1	
ir k	o->1	
ir l	a->1	e->1	u->1	ä->2	
ir m	e->4	i->1	y->2	å->1	ö->3	
ir n	a->1	e->1	å->2	ö->1	
ir o	f->1	n->1	t->1	u->1	
ir r	a->1	e->1	ä->1	
ir s	a->2	e->2	k->1	o->1	t->3	v->2	ä->1	å->1	
ir t	i->4	ä->1	
ir u	t->2	
ir v	a->1	e->2	i->1	
ir ä	n->1	
ir å	s->1	
ir ö	v->1	
ir, 	g->1	i->1	
ir: 	O->1	
ira 	R->1	m->1	ä->1	
ira,	 ->2	
ira.	J->1	
irak	e->1	i->1	
irar	 ->1	e->1	n->1	
irat	e->1	
ire 	h->1	
ire,	 ->1	
ire-	A->1	
ire.	D->1	
iref	o->4	
ireg	l->3	
irek	t->257	
irer	.->1	a->3	
irgi	z->5	
irig	e->1	
irka	 ->4	
irke	l->1	s->3	
irkl	a->2	
irku	l->3	
irlä	n->11	
irma	n->1	
irmo	u->1	
iron	i->2	
irra	 ->1	d->2	n->1	t->3	
irre	p->1	
irrg	å->1	
irri	n->8	t->4	
irrv	a->1	
irta	n->1	
is (	P->1	
is -	 ->3	
is A	l->1	
is B	a->1	
is G	o->1	
is M	i->1	
is P	a->1	
is W	u->1	
is a	l->3	n->5	t->13	v->6	
is b	a->2	e->4	r->2	å->1	
is d	e->12	ä->2	
is e	l->2	n->4	t->2	x->1	
is f	i->2	o->2	r->4	u->2	y->1	å->2	ö->8	
is g	e->2	o->3	r->1	ä->1	å->2	
is h	a->10	e->1	j->1	o->1	ä->2	ö->1	
is i	 ->7	l->1	n->20	
is j	u->2	
is k	a->2	e->1	o->5	
is l	a->2	e->1	i->6	o->1	
is m	e->4	i->3	y->1	å->4	
is n	ä->3	
is o	a->1	c->18	m->5	r->1	t->1	
is p	e->2	o->1	r->2	å->10	
is r	a->1	e->1	o->1	ä->1	
is s	a->3	e->1	i->1	j->1	k->11	m->1	o->25	t->4	v->1	ä->2	å->3	
is t	a->1	e->1	i->2	
is u	n->2	p->2	t->4	
is v	a->2	i->8	ä->4	
is ä	n->2	r->15	v->4	
is å	s->1	t->3	
is ö	v->3	
is! 	V->1	
is) 	f->1	
is, 	E->1	a->2	d->4	e->1	i->1	k->2	m->2	n->1	o->3	p->1	s->2	t->1	v->1	
is-J	ø->2	
is-f	ö->1	
is-n	o->1	
is-p	r->1	
is. 	M->1	
is.D	a->1	e->2	å->1	
is.E	f->1	
is.F	ö->2	
is.H	u->1	
is.J	a->2	
is.M	e->1	
is.S	a->1	e->1	
is.V	i->1	
is.Ä	n->1	
is: 	f->1	
is; 	a->1	
is?Ä	r->1	
isa 	(->1	R->1	a->7	b->2	d->4	e->2	f->2	g->1	h->2	i->8	k->1	l->1	m->1	o->3	p->4	s->9	t->10	u->1	v->4	ä->3	
isa,	 ->8	
isa.	.->1	B->1	D->4	E->1	F->1	J->1	K->1	R->1	S->1	U->1	Å->1	
isa?	P->1	
isab	e->1	
isad	e->19	
isak	a->1	
isan	 ->4	.->1	d->2	s->1	
isar	 ->66	,->2	.->1	e->2	
isas	 ->9	,->1	
isat	 ->32	,->1	.->2	i->43	o->1	s->3	
isav	i->1	
isba	r->1	
isbe	s->9	t->1	
isbö	r->7	
isca	y->6	
isce	n->1	
isch	!->1	l->4	
isci	p->14	
isda	g->2	
isdi	k->5	
isdo	m->1	
ise 	G->1	
isee	n->1	
isek	t->8	
isem	i->3	
isen	 ->11	.->4	b->3	s->1	
iser	 ->6	,->1	.->3	a->102	i->89	n->4	
ises	 ->2	
iset	 ->13	.->2	
isfi	s->3	
isfö	r->1	
ish 	P->1	
ishe	t->3	
isio	n->27	
isis	k->70	
isit	i->1	
isiä	r->1	
isk 	-->1	a->19	b->20	c->2	d->14	e->2	f->18	g->8	h->8	i->13	j->5	k->32	l->15	m->15	n->18	o->27	p->26	r->19	s->29	t->9	u->23	v->4	ä->1	å->13	ö->3	
isk,	 ->7	
isk-	i->1	s->1	
isk.	 ->1	D->1	H->2	I->3	J->1	M->1	O->1	V->1	
iska	 ->1341	,->12	.->5	:->1	b->1	d->2	n->6	r->4	s->1	
iskb	e->8	
iske	 ->13	)->2	,->4	.->2	k->1	m->4	n->17	o->2	r->46	s->1	t->8	v->2	
iskf	a->1	r->1	y->1	ö->1	
iskh	a->6	
iskk	a->1	o->2	
iskn	i->1	
isko	f->2	h->3	l->3	r->82	s->1	
iskr	e->1	i->20	
iskt	 ->244	!->1	,->7	.->10	
isku	p->1	s->61	t->81	
iskv	o->2	ä->3	
islä	p->2	
ism 	-->1	e->3	h->1	i->1	m->1	o->18	p->1	s->5	u->1	ä->2	ö->1	
ism,	 ->11	
ism.	D->7	F->1	H->1	I->2	J->1	M->1	N->1	O->2	V->4	
ism?	V->1	
isme	d->2	n->22	r->9	
ismi	s->2	
ismy	n->2	
isni	n->14	v->1	
isnå	l->1	
isol	e->7	
isom	r->1	
ison	t->3	
isor	.->2	i->2	n->1	
ispe	n->1	
ispl	i->1	
ispo	s->3	
isra	e->20	
iss 	b->2	f->5	h->1	i->2	m->8	o->5	p->3	r->1	s->3	t->5	u->2	v->2	å->3	ö->1	
iss,	 ->5	
iss.	D->1	E->1	
issa	 ->141	.->1	b->8	d->2	m->1	r->1	t->1	
issb	r->10	
isse	n->1	r->17	
issf	a->1	o->2	ö->4	
issg	y->7	
issh	e->4	u->1	
issi	o->1151	t->1	
issk	ö->6	
issl	a->1	y->18	ö->1	
issn	ö->3	
isso	 ->5	,->1	
issr	e->2	
isst	 ->7	a->15	e->5	o->1	r->3	y->2	ä->4	
issu	p->2	
issy	s->1	
issä	n->1	
ist 	E->3	P->1	a->6	b->1	f->7	k->2	m->2	n->1	o->3	p->19	s->4	u->1	v->2	ä->2	
ist!	T->1	
ist,	 ->5	
ist.	G->1	
ista	 ->50	,->1	.->6	?->1	N->1	l->2	n->80	s->3	t->2	
istd	e->11	
iste	 ->3	f->1	l->1	n->22	r->157	
istf	l->1	ä->8	
istg	r->3	
isth	a->1	
isti	g->3	k->6	n->2	s->81	
istk	o->1	
istl	i->1	
istn	ä->2	
isto	r->36	
istp	a->5	
istr	a->40	e->11	i->2	
ists	 ->1	e->2	
isty	r->4	
istä	l->2	
istå	 ->1	e->1	n->22	t->1	
isua	l->1	
isue	l->1	
isum	 ->1	
isut	v->1	
isvä	s->1	
isys	t->1	
isäk	e->7	
isär	 ->3	e->1	
it -	 ->2	
it F	P->1	
it a	k->2	l->3	n->2	r->1	t->6	v->2	
it b	e->2	i->2	o->2	ä->1	å->1	
it d	e->9	i->1	ä->3	
it e	f->3	l->1	n->22	r->1	t->12	
it f	a->2	e->2	i->1	l->1	r->15	ö->8	
it g	a->1	o->1	
it h	a->2	u->1	ä->8	ö->7	
it i	 ->8	g->1	n->7	
it k	o->3	ä->2	
it l	a->1	e->3	i->1	o->1	ä->1	å->1	
it m	e->8	i->3	o->2	y->4	ä->1	ö->3	
it n	i->1	y->1	ä->1	å->4	ö->1	
it o	c->4	e->1	f->2	m->2	
it p	e->1	l->1	o->1	r->1	å->8	
it r	i->2	u->1	
it s	e->1	i->12	j->2	k->1	n->1	o->1	p->1	t->8	v->1	y->1	ä->1	å->5	
it t	a->1	i->18	o->1	y->2	
it u	n->6	p->15	t->4	
it v	a->4	i->4	
it ä	n->1	
it å	t->1	
it ö	v->7	
it, 	b->1	e->2	f->1	m->1	o->1	v->1	ä->1	
it-a	n->5	
it.F	r->2	ö->3	
it.I	 ->1	
it.M	e->1	o->1	
it.N	ä->1	
it.P	a->1	
ita 	h->1	i->3	o->3	p->2	s->1	u->1	v->1	ä->1	
ita,	 ->1	
ita.	D->1	M->1	S->1	
itad	e->1	
ital	 ->5	,->1	.->1	e->5	i->20	s->3	
itam	e->8	
itan	,->1	n->14	o->1	s->1	
itar	 ->9	i->4	
itas	,->1	
itat	.->2	i->12	
itau	e->1	
itbo	k->53	
ite 	b->1	e->1	i->1	m->1	s->1	
itel	 ->6	n->1	
iten	 ->20	.->2	
iter	 ->2	,->1	-->1	.->1	a->27	i->37	s->1	
itet	 ->125	!->1	,->35	.->30	:->2	?->3	e->75	s->40	
ithö	r->1	
itia	t->80	
itic	a->1	
itie	-->1	d->2	m->3	r->2	
itik	 ->120	!->1	"->1	,->29	.->25	?->2	e->140	o->6	s->1	
itim	a->7	e->5	i->6	t->3	
itin	 ->1	.->1	
itio	 ->1	n->79	
itis	e->10	h->1	k->247	m->2	
itiv	 ->20	,->1	a->26	l->2	t->36	
itiö	s->12	
itla	n->2	
itle	k->1	r->6	
itli	g->5	
itlä	n->1	
itni	n->1	
itor	i->25	
itra	k->5	
itre	a->1	
itro	v->1	
itru	s->1	t->1	
its 	a->8	b->1	d->1	e->1	f->4	g->1	h->1	i->10	m->4	n->3	o->3	p->4	s->2	t->2	u->7	ä->2	
its,	 ->4	
its.	B->1	D->2	M->1	S->1	
itt 	2->1	a->25	b->12	d->3	e->14	f->16	g->2	h->5	i->8	j->1	k->3	l->19	m->9	o->1	p->10	r->5	s->16	t->10	u->6	v->2	y->5	ä->4	ö->2	
itt,	 ->3	
itt.	M->1	
itta	 ->26	d->1	n->2	r->9	t->2	
itte	n->4	r->23	t->3	
itti	l->44	n->1	s->16	
ittl	i->1	
ittn	a->3	e->2	i->2	
ittr	a->4	i->2	
itts	b->1	r->1	
itté	 ->10	e->4	f->2	n->41	s->2	
itu 	m->20	
itua	t->129	
itud	 ->1	
itue	r->1	
itul	e->2	
itum	.->1	
itut	i->158	
ityd	 ->4	.->1	
itz 	i->1	
itz.	 ->1	
itär	 ->2	a->3	e->1	t->1	
ium 	a->2	b->1	e->1	i->2	m->1	o->3	s->3	
ium!	D->1	
ium,	 ->4	
ium.	A->2	D->1	H->1	L->1	P->1	R->1	S->1	Ä->1	
iuts	k->1	
iv (	K->1	
iv -	 ->3	
iv 9	3->1	4->2	6->5	
iv E	n->1	
iv a	n->3	t->2	v->2	
iv b	a->1	e->1	l->1	
iv d	e->2	i->2	
iv e	f->1	k->2	n->4	
iv f	a->1	r->5	å->2	ö->10	
iv g	e->1	
iv h	a->7	j->1	
iv i	 ->6	m->1	n->7	
iv k	a->3	o->8	v->1	
iv l	a->2	e->1	i->3	ä->1	ö->1	
iv m	e->2	i->2	o->1	å->1	
iv o	a->1	c->9	m->21	p->1	
iv p	o->1	å->7	
iv r	e->1	i->1	o->2	
iv s	a->1	e->2	i->1	k->2	n->1	o->26	t->9	y->3	å->4	
iv t	a->1	i->15	r->1	
iv u	t->3	
iv v	e->1	i->4	ä->1	
iv ä	n->1	r->5	
iv å	t->2	
iv ö	v->1	
iv, 	9->1	a->1	b->1	d->3	e->1	h->1	i->1	j->1	l->1	m->2	n->1	o->5	s->6	t->1	u->1	
iv. 	V->1	
iv..	 ->1	H->1	
iv.A	t->1	v->1	
iv.B	l->1	
iv.D	e->5	å->1	
iv.E	n->1	
iv.F	ö->4	
iv.I	 ->2	n->1	
iv.L	å->1	
iv.M	e->2	
iv.O	m->1	
iv.R	i->1	
iv.S	å->1	
iv.V	i->2	
iv.Y	t->1	
iv: 	F->1	v->1	
iv; 	a->1	
iv?F	ö->1	
iv?N	e->1	
iva 	a->5	b->9	c->1	d->13	e->14	f->9	g->1	h->3	i->7	k->12	l->2	m->3	n->2	o->13	p->10	r->9	s->11	t->11	u->3	v->3	å->4	ö->1	
iva,	 ->4	
iva.	A->1	H->1	V->1	
ivad	e->1	
ivan	d->24	
ivar	e->46	k->1	l->1	n->14	p->1	
ivas	 ->6	,->1	.->2	t->1	
ivat	 ->2	.->1	a->16	e->1	i->3	s->3	
ivav	t->7	
ivbe	t->1	
ivbo	r->1	
ive 	E->1	a->2	b->4	d->4	e->3	f->1	k->4	l->2	m->2	p->3	r->3	s->1	t->2	
ivel	 ->25	,->2	a->3	s->8	
iven	 ->18	,->2	.->1	h->4	s->1	
iver	 ->22	,->1	.->1	a->15	i->4	s->8	
ives	 ->1	
ivet	 ->88	"->1	,->13	.->20	s->10	v->27	
ivfö	r->4	
ivid	 ->2	e->4	u->8	
ivie	n->1	r->1	
ivil	 ->5	-->1	a->3	b->2	e->6	f->2	i->3	l->12	r->1	s->2	t->1	
ivis	e->3	m->1	
ivit	 ->38	.->1	e->39	s->10	
ivkr	a->3	
ivla	 ->1	.->1	d->1	r->5	t->2	
ivli	g->3	s->2	
ivna	 ->9	
ivni	n->11	
ivra	s->1	
ivri	k->1	
ivrä	t->4	
ivs 	a->2	e->2	g->1	i->6	s->1	ö->1	
ivs,	 ->1	
ivs.	D->1	
ivsc	y->3	
ivsd	u->2	
ivsk	r->1	v->5	
ivsm	e->88	i->3	
ivsu	p->1	
ivsv	i->1	
ivt 	-->1	a->11	b->4	d->2	e->1	f->7	h->1	i->8	k->3	m->4	n->1	o->17	p->4	r->4	s->29	t->6	u->2	v->1	y->1	ä->1	å->2	ö->1	
ivt,	 ->7	
ivt.	 ->1	D->2	E->1	I->1	P->1	Ä->1	
iväg	 ->2	,->1	
ivå 	-->1	a->3	d->1	f->5	g->2	h->1	i->4	m->4	n->1	o->7	p->2	s->9	u->3	v->1	ä->2	
ivå,	 ->13	
ivå.	A->1	B->1	D->7	F->1	G->1	H->2	J->4	M->1	N->1	P->1	V->1	
ivå;	 ->1	
ivå?	S->1	
ivåe	r->14	
ivåg	r->3	
ivån	 ->8	.->4	
iwan	 ->1	
ix.D	e->1	
ixas	 ->5	
ixen	 ->1	
ixtr	a->1	
iz e	l->1	
iz f	å->1	ö->1	
iz s	o->1	
iz, 	G->1	t->1	
iz-k	a->1	
izis	t->5	
iäke	r->1	
iär,	 ->1	
iära	 ->1	
iäre	r->4	
iärm	i->10	
iärp	l->1	
iåld	e->1	
iåte	r->1	
ière	 ->1	
ié u	t->1	
iös 	d->1	o->1	s->1	u->1	
iös,	 ->1	
iösa	 ->9	,->1	.->1	r->2	
iöst	 ->6	
j 19	9->3	
j 20	0->1	
j Li	b->1	
j an	g->1	
j at	t->1	
j av	g->1	
j be	r->1	s->1	
j bo	r->1	
j fö	r->3	
j i 	f->1	
j ko	m->1	
j lå	n->1	
j lö	s->1	
j mo	t->1	
j nä	r->1	
j om	 ->1	
j ti	l->1	
j är	 ->1	
j öv	e->1	
j, b	e->1	i->1	
j, d	e->1	
j, h	e->1	
j, j	a->1	
j, m	a->2	
j, n	a->1	
j, o	c->1	m->1	
j, s	k->1	ä->1	
j, ä	v->1	
j-va	n->1	
j.(A	p->1	
j.De	 ->1	
j.Ex	p->1	
j.I 	s->1	
j.Ja	g->1	
j.Rå	d->1	
j.To	n->1	
j.Vi	 ->1	
ja -	 ->3	
ja D	a->1	
ja F	N->1	
ja H	a->2	
ja J	ö->1	
ja M	a->1	
ja a	l->4	n->13	r->4	t->10	v->1	
ja b	e->12	o->1	ö->5	
ja c	h->1	i->1	
ja d	e->47	i->1	
ja e	f->2	k->1	l->2	n->15	r->3	t->4	
ja f	o->2	r->13	u->2	ä->1	ö->21	
ja g	e->4	r->5	ö->10	
ja h	a->8	u->1	ä->2	å->1	ö->2	
ja i	 ->4	n->2	
ja k	l->1	n->1	o->5	r->2	u->2	v->3	ö->1	
ja l	e->1	i->2	o->1	y->1	ä->2	
ja m	e->36	i->4	y->1	
ja n	y->1	ä->3	
ja o	c->7	l->1	m->1	s->8	
ja p	a->1	e->1	r->1	å->10	
ja r	e->3	i->1	ä->3	
ja s	a->3	e->2	i->9	k->1	l->1	o->2	t->5	v->1	y->3	ä->20	
ja t	.->1	a->18	i->14	v->1	ä->1	
ja u	n->5	p->11	r->1	t->6	
ja v	a->4	e->4	i->1	å->2	
ja y	r->1	t->1	
ja Ö	s->1	
ja å	t->6	
ja ö	v->1	
ja, 	d->2	f->1	g->1	h->1	l->1	m->1	p->1	t->2	v->1	
ja..	.->1	
ja.H	e->1	
ja.J	a->2	
ja.K	o->1	
ja.M	i->1	
ja.T	r->1	
ja.V	i->1	
jade	 ->15	s->3	
jag 	-->5	1->1	G->1	a->111	b->36	c->2	d->14	e->24	f->75	g->25	h->78	i->73	j->1	k->57	l->15	m->46	n->23	o->29	p->18	r->23	s->119	t->102	u->30	v->116	ä->40	å->4	ö->1	
jag,	 ->15	
jag.	 ->1	S->1	
jaga	r->2	
jakt	 ->4	i->6	l->14	
jala	 ->2	
jali	s->4	t->1	
jamo	,->1	
jan 	a->11	d->1	e->2	f->5	g->1	h->2	i->3	o->2	p->2	t->1	u->2	
jan,	 ->3	
jana	l->1	
jand	e->77	
janu	a->16	
japa	n->1	
jar 	a->3	b->3	d->4	e->4	f->1	g->1	k->1	m->4	n->1	o->4	p->3	r->2	s->3	t->3	u->1	å->1	
jar.	D->1	M->1	
jarb	a->1	
jard	 ->1	e->14	
jare	 ->4	.->2	n->2	
jarn	a->6	
jas 	a->8	f->8	g->1	i->2	m->1	o->2	s->1	u->1	å->1	
jas,	 ->4	
jas.	H->2	M->2	N->1	V->1	
jat 	-->1	a->2	f->1	h->1	j->1	l->1	m->1	o->1	s->5	t->1	v->1	
jat.	I->1	J->1	
jata	 ->1	
jats	 ->2	,->2	
jd -	 ->1	
jd a	t->1	v->18	
jd g	a->1	
jd m	e->1	
jd p	å->1	
jd s	ä->1	
jd u	t->1	
jd.J	a->1	
jda 	m->7	
jda,	 ->3	
jdas	 ->1	
jdat	 ->1	
jde 	a->1	b->1	d->1	p->1	s->1	u->1	
jden	 ->1	
jder	 ->10	n->9	
jdes	 ->2	
jdos	k->1	
jdpu	n->2	
jdri	k->1	
jdsk	a->2	
jdåt	g->1	
je (	B->1	
je -	 ->1	
je 1	0->1	
je B	a->1	
je E	U->1	u->1	
je a	n->2	s->1	t->1	v->1	
je b	e->3	i->1	o->1	
je d	a->7	e->3	i->1	
je e	n->5	u->2	
je f	a->6	i->1	o->6	r->2	ö->4	
je g	a->1	e->1	r->1	ä->1	å->4	
je h	a->2	
je i	n->3	
je k	o->2	u->1	
je l	a->31	ä->2	
je m	e->14	i->2	å->4	
je n	o->1	
je o	a->1	c->4	
je p	e->1	r->1	u->4	
je r	e->2	i->2	ä->1	
je s	a->2	o->5	t->3	u->1	
je v	i->2	ä->2	
je ä	r->1	
je å	r->10	t->1	
je ö	v->3	
je, 	a->3	v->1	
je- 	o->1	
je.G	e->1	
je.J	a->1	
je: 	u->1	
jebe	f->1	
jebo	l->4	
jebä	l->10	
jede	l->6	
jedo	m->1	
jefa	d->1	
jefö	r->2	
jein	d->3	
jejo	r->3	
jeko	k->1	n->1	
jekt	 ->29	"->1	,->6	.->2	?->2	a->2	e->23	i->3	
jela	n->6	
jeli	n->1	
jels	e->4	
jemä	s->1	
jen 	b->1	h->1	i->1	
jen.	D->1	
jer 	9->1	a->2	b->1	d->4	e->2	f->10	g->2	h->2	i->7	j->1	k->2	l->1	m->6	n->3	o->9	p->2	r->1	s->18	u->2	v->4	ä->1	å->1	
jer"	.->1	
jer,	 ->10	
jer.	D->1	H->1	M->1	V->1	
jer:	 ->1	
jera	d->11	t->5	
jern	a->35	
jesk	a->1	
jest	a->1	
jet 	a->2	
jeta	n->9	
jetr	a->1	u->1	
jett	i->1	o->1	
jeut	s->2	
jevä	c->3	
jeåt	e->1	
jflö	d->1	
jiki	s->5	
jkan	 ->1	
jkon	t->2	
jkot	t->1	
jlig	 ->8	.->2	a->31	e->6	g->12	h->131	t->119	
jnin	g->19	
jobb	 ->2	,->2	
jock	 ->1	a->1	
jol 	o->2	
jol,	 ->1	
jol.	K->1	
jon 	i->1	
jone	r->63	
joni	s->1	
jont	a->1	
jor 	o->1	
jor.	F->1	
jord	 ->1	.->2	a->3	b->64	e->41	m->1	s->1	
jori	t->42	
jorn	a->1	
jort	 ->58	,->8	.->6	o->9	s->23	
jos 	a->1	
jour	n->3	
jovi	s->17	
js a	v->1	
js k	a->1	
js o	c->1	
js t	i->1	
js u	p->2	
js, 	f->1	
js.(	E->1	
jsmå	l->2	
jt i	 ->1	
jt o	s->1	
jt s	i->1	
jt u	t->1	
jt v	i->1	
jts 	t->2	u->1	
jts,	 ->1	
ju E	g->1	
ju M	o->1	
ju a	b->1	l->5	n->1	t->3	v->1	
ju b	a->2	
ju d	e->2	i->1	ä->1	å->1	
ju e	m->1	n->1	
ju f	ö->2	
ju g	å->1	
ju h	ä->1	
ju i	n->11	s->1	
ju l	ä->1	
ju m	e->5	o->1	å->1	
ju o	c->7	f->1	
ju p	a->1	o->1	u->1	å->1	
ju r	e->3	
ju s	a->2	i->1	o->1	t->3	
ju t	i->1	
ju u	t->1	
ju v	i->1	
ju ä	n->2	r->5	
ju, 	o->1	p->1	å->1	
juad	e->1	
jubl	a->1	
juda	 ->15	n->5	r->1	s->2	
judd	a->1	
jude	n->1	r->12	t->4	u->1	
judi	c->1	k->3	s->1	t->1	
judl	i->1	
judn	a->2	i->1	
juge	r->1	
jugo	 ->2	f->1	n->1	
juk.	J->1	
juka	 ->1	,->1	
jukd	o->1	
jukf	ö->1	
jukh	u->7	
jukn	i->2	
jukv	å->3	
jul 	o->1	
julf	e->1	
juli	 ->8	,->2	
julk	l->1	
jund	e->4	
jung	e->2	f->1	
juni	 ->12	
junk	a->4	e->2	i->2	n->1	t->1	
jup 	ö->1	
jupa	 ->5	,->1	d->1	r->1	s->3	t->2	
jupe	t->5	
jupg	å->7	
jupn	i->5	
jups	i->1	
jupt	 ->7	
jur 	o->1	ä->1	
jur,	 ->2	
jur-	 ->2	
jur.	D->1	H->1	
jura	r->1	
jure	n->1	t->1	
jurf	o->4	
juri	d->30	s->17	
jurl	i->2	
jus 	p->1	
jus.	I->1	
juse	t->8	
just	 ->91	,->1	.->2	:->1	e->6	i->10	
juta	 ->9	n->1	s->3	
jute	n->2	r->6	
juti	t->5	
jutn	i->1	
juts	 ->5	
jutt	o->2	
jutv	a->1	
juve	l->2	
jäl 	d->1	
jäl,	 ->1	
jäl.	F->2	
jäle	n->2	
jälp	 ->48	,->2	.->5	a->41	e->5	l->1	s->1	t->3	v->1	
jält	 ->3	
jälv	 ->39	,->5	.->4	a->69	b->5	f->3	h->1	k->21	p->1	s->16	t->5	ä->1	
jämf	ö->16	
jämk	a->2	
jäml	i->13	
jämn	 ->1	,->1	.->1	a->5	i->2	v->1	
jäms	i->1	t->23	
jämt	 ->2	.->1	
jämv	i->2	
jäna	 ->4	d->1	r->16	
jäns	t->123	
jänt	 ->2	a->27	
jära	.->1	
järd	e->11	
järe	r->1	
järn	-->2	a->2	v->15	
järt	a->20	l->7	
järv	 ->1	a->3	h->1	t->2	
jätt	e->21	
jävu	l->2	
jö f	ö->2	
jö i	 ->1	
jö k	a->1	
jö m	o->1	
jö s	a->1	o->1	
jö v	i->1	
jö!D	e->1	
jö, 	f->7	h->1	l->1	s->1	u->1	
jö- 	o->2	
jö.D	e->2	å->1	
jö.M	e->1	
jö.U	n->1	
jö.V	i->1	
jöan	p->1	s->2	
jöav	t->1	
jöbe	l->1	s->2	
jöbr	o->1	
jöd 	f->1	
jöde	p->1	
jödi	r->1	
jöds	 ->1	
jöer	 ->3	n->1	
jöfa	k->1	r->9	
jöfr	å->4	
jöfö	r->4	
jöin	f->1	
jöka	s->1	t->10	
jöko	n->6	
jökr	a->8	
jökv	a->1	
jöla	g->1	
jömi	n->1	
jömä	n->2	s->11	
jömå	l->3	
jön 	e->2	f->1	h->1	i->1	o->6	p->1	s->1	t->1	ä->1	
jön!	D->1	
jön,	 ->9	
jön.	D->3	E->1	F->1	J->1	L->1	M->1	U->1	V->2	
jönk	 ->3	.->1	
jöno	r->2	
jöns	 ->2	
jöom	r->4	
jöov	ä->1	
jöpe	r->1	
jöpo	l->8	
jöpr	o->4	
jöpå	v->1	
jör 	-->2	
jörå	d->1	
jörö	r->2	
jöse	k->1	
jösi	d->1	
jösk	a->2	y->11	ä->2	
jöss	 ->3	)->1	
jöst	e->4	ö->1	
jösy	n->6	
jötr	a->1	
jöut	s->1	
jövä	n->7	r->3	
k - 	d->3	n->1	o->1	v->1	
k De	t->1	
k Jö	r->1	
k Ki	r->1	
k TV	 ->1	
k a 	p->1	
k ag	i->1	
k al	-->1	l->8	
k an	a->1	d->1	g->2	t->2	v->1	
k ar	t->3	
k as	p->1	
k at	t->24	
k av	 ->13	
k ba	k->1	l->2	r->2	s->2	
k be	l->1	r->2	s->4	t->5	
k bi	l->4	
k bl	i->1	o->1	
k bo	j->1	r->1	
k br	o->1	
k by	g->1	r->2	
k bö	j->1	
k ci	v->2	
k da	g->2	
k de	 ->1	b->4	m->2	n->1	t->6	
k di	a->2	m->1	s->4	
k ef	t->3	
k eg	e->1	
k ej	 ->1	
k ek	o->1	
k el	l->4	
k em	e->1	
k en	 ->5	e->1	i->1	
k er	s->1	
k et	a->1	t->1	
k fe	d->1	
k fi	e->1	l->1	n->2	
k fl	a->2	
k fo	n->1	r->2	
k fr	a->2	u->2	ä->1	å->7	
k fy	s->1	
k få	 ->1	r->2	
k fö	r->50	
k ga	v->1	
k ge	m->1	n->3	s->1	
k gj	o->1	
k gl	u->1	
k gr	a->1	u->1	ö->2	
k gä	l->3	
k gå	r->2	
k ha	m->1	n->4	r->12	
k he	l->1	
k hj	ä->2	
k ho	n->2	p->1	
k hu	r->1	v->1	
k hä	n->2	
k hö	r->3	
k i 	A->2	E->2	K->1	L->1	T->2	W->1	a->1	d->1	e->1	f->4	g->1	h->1	k->2	m->1	n->1	o->1	r->1	s->4	u->1	v->2	
k id	e->1	
k im	m->1	
k in	 ->1	d->1	g->1	l->1	o->2	r->3	s->5	t->15	
k ja	g->4	
k jo	r->1	
k ju	 ->2	r->1	s->1	
k jä	m->1	t->1	
k ka	m->1	n->10	r->1	t->3	
k kl	a->1	o->1	
k ko	m->6	n->23	s->1	
k ku	l->3	n->1	r->1	
k kv	i->1	
k kä	n->2	
k la	g->5	
k le	d->2	g->3	
k li	v->5	
k lo	v->1	
k ly	c->1	
k lä	g->1	k->1	n->1	
k lö	s->1	
k ma	k->3	r->2	t->1	
k me	d->13	l->2	n->1	r->1	
k mi	g->1	l->2	n->1	s->1	
k mo	d->2	t->5	
k my	c->2	n->3	
k må	s->6	
k mö	j->2	
k na	t->3	
k ne	d->1	
k ni	v->14	
k nj	u->1	
k nu	 ->1	
k ny	a->1	
k nä	r->5	
k nå	g->3	
k oc	h->72	k->2	
k of	f->4	
k oj	ä->1	
k om	 ->10	s->1	
k op	e->1	
k or	i->1	
k os	s->3	
k pa	r->3	
k pe	r->2	
k pl	a->2	
k po	l->19	ä->1	
k pr	o->5	
k pu	n->1	
k på	 ->13	
k ra	k->1	m->1	s->1	
k re	a->1	f->3	g->3	k->1	n->2	t->1	
k ri	s->1	
k ro	l->5	
k rä	t->1	
k rå	d->1	
k rö	r->2	
k sa	d->2	m->1	
k se	 ->1	g->1	n->1	
k si	g->2	t->3	
k sj	ä->1	
k sk	a->5	u->1	y->1	ö->1	
k sm	i->1	
k sn	a->1	
k so	l->2	m->58	
k st	a->8	r->8	
k sv	å->1	
k sy	n->6	
k sä	g->1	k->1	r->1	
k så	 ->16	d->1	
k te	r->1	
k ti	g->1	l->29	
k tr	a->2	o->1	
k tv	i->1	u->1	
k ty	p->1	
k tä	n->1	
k un	d->3	i->5	
k up	p->6	
k ur	s->1	
k ut	 ->1	a->1	b->2	g->1	m->2	t->1	v->9	
k va	d->1	r->10	
k ve	r->1	
k vi	 ->4	d->4	k->1	l->8	n->1	t->1	
k vä	g->3	r->1	
k än	 ->1	n->1	
k är	 ->12	
k åk	l->13	
k åt	e->1	m->2	
k öv	e->4	n->1	
k!An	d->1	
k!Om	 ->1	
k" -	 ->1	
k" f	ö->1	
k" o	c->1	
k, 1	5->1	
k, R	e->1	
k, a	t->1	
k, b	e->1	
k, d	e->9	v->2	å->2	
k, e	f->2	n->2	x->1	
k, f	i->1	r->6	ö->3	
k, g	o->1	å->1	
k, h	a->1	e->6	ä->1	
k, i	 ->2	n->4	
k, k	o->5	ä->1	
k, m	e->8	o->1	
k, n	e->1	ä->2	å->1	
k, o	c->3	
k, s	a->2	k->1	o->6	å->2	
k, t	i->1	r->12	
k, u	t->1	
k, v	a->2	i->2	ä->1	
k, ä	r->1	
k- e	l->1	
k- o	c->2	
k-br	i->1	
k-da	m->1	
k-fr	a->1	
k-is	r->1	
k-po	s->1	
k-sk	a->1	
k. D	e->1	
k. J	a->1	
k. M	e->1	
k. a	n->1	
k. i	n->1	
k. s	k->1	o->1	
k..(	F->1	
k.At	t->2	
k.Av	g->1	
k.Be	t->1	
k.By	g->1	
k.De	 ->3	n->1	t->16	
k.Dä	r->1	
k.Då	 ->2	
k.En	 ->1	
k.Et	t->1	
k.Eu	r->1	
k.Fa	k->1	
k.Fr	u->1	å->3	
k.Fö	r->1	
k.Ge	n->1	
k.Ha	n->2	
k.He	r->7	
k.Hi	t->1	
k.Hu	r->1	
k.Hä	r->1	
k.I 	b->1	d->1	g->1	
k.In	f->1	
k.Ja	g->7	
k.Ki	n->1	
k.Ko	m->1	
k.Me	n->3	
k.Ni	 ->1	
k.Oc	h->1	
k.Om	 ->1	
k.Re	f->1	
k.Ri	k->1	
k.Sy	r->1	
k.Ta	c->1	
k.Tr	ä->1	
k.Tv	ä->1	
k.Ty	v->1	
k.Va	n->1	
k.Vi	 ->8	l->1	
k.Äv	e->2	
k: g	e->1	
k: v	i->1	
k?He	r->1	
k?Ne	j->1	
k?Re	g->1	
k?Va	d->1	
ka "	s->1	
ka -	 ->4	
ka 1	7->1	
ka 2	5->1	
ka A	h->1	
ka B	a->1	
ka E	U->1	u->5	
ka F	P->1	l->1	
ka G	r->2	
ka K	a->1	o->1	u->1	
ka L	a->1	
ka P	V->1	a->2	o->2	
ka S	c->1	
ka T	V->1	
ka a	b->1	k->3	l->15	m->1	n->19	r->18	s->2	t->37	u->1	v->8	
ka b	a->4	e->50	i->16	l->2	o->1	r->2	u->6	y->4	å->1	ö->2	
ka c	e->3	
ka d	a->1	e->78	i->6	j->2	o->4	u->1	y->2	ä->1	
ka e	f->6	k->9	l->2	m->1	n->14	r->9	t->8	u->2	x->5	
ka f	a->13	i->5	l->3	o->36	r->28	u->2	y->1	å->3	ö->107	
ka g	a->3	e->25	i->3	r->33	ä->2	
ka h	a->14	e->10	i->4	j->1	o->2	u->4	ä->5	å->6	ö->2	
ka i	 ->21	d->1	h->1	m->1	n->96	s->1	
ka j	a->1	o->2	ä->3	
ka k	a->16	i->1	l->3	o->134	r->21	u->18	v->4	y->1	ä->4	
ka l	a->5	e->13	i->16	o->3	ä->17	ö->2	
ka m	a->11	e->49	i->28	o->8	y->19	ä->1	å->20	ö->7	
ka n	a->11	e->1	i->3	o->2	u->1	y->2	ä->7	å->2	ö->2	
ka o	b->1	c->68	e->1	f->6	i->1	k->1	l->1	m->20	n->1	p->2	r->80	s->1	
ka p	a->22	e->7	l->8	o->21	r->37	u->7	å->27	
ka r	a->20	e->72	i->11	u->1	ä->8	å->22	ö->4	
ka s	a->15	c->2	e->6	i->32	j->4	k->21	l->5	o->32	p->4	t->52	v->7	y->14	ä->7	å->3	
ka t	a->5	e->12	i->31	j->2	o->1	r->9	v->1	y->5	ä->1	
ka u	m->1	n->251	p->7	t->39	
ka v	a->24	e->15	i->21	o->3	ä->15	å->7	
ka ä	g->1	m->1	n->8	r->10	v->2	
ka å	k->4	t->28	
ka ö	a->1	g->1	p->1	s->1	v->8	
ka",	 ->1	
ka, 	a->1	b->1	d->2	e->3	f->5	h->3	j->1	k->1	m->4	n->2	o->4	r->1	s->9	t->2	v->3	ä->1	ö->1	
ka-o	l->1	
ka.(	I->1	
ka.B	o->1	
ka.D	e->4	
ka.E	f->1	m->1	n->2	
ka.F	ö->1	
ka.H	e->1	u->1	
ka.I	 ->3	
ka.J	a->5	
ka.L	å->1	
ka.M	e->1	i->1	
ka.O	c->1	
ka.P	å->2	
ka.R	å->1	
ka.T	a->1	
ka.V	a->1	e->1	i->3	
ka.Å	 ->1	
ka: 	"->1	a->1	
ka?"	J->1	
ka?I	 ->1	
kaba	r->1	
kabe	h->1	k->1	l->1	
kabi	n->3	
kad 	a->7	d->1	e->1	f->2	i->2	j->1	k->6	m->1	p->3	r->1	s->9	t->2	u->1	ö->1	
kad.	D->1	
kada	 ->9	!->1	,->1	.->1	d->2	n->3	r->6	t->4	
kade	 ->35	,->1	.->4	e->2	f->1	m->2	s->15	
kadi	n->1	
kadl	i->10	
kadm	i->3	
kado	r->26	
kadr	a->3	
kaff	a->25	e->1	
kafr	å->1	
kagå	n->4	
kaka	d->1	t->1	
kal 	a->1	b->1	f->1	n->2	o->1	p->1	s->3	
kal:	 ->1	
kala	 ->39	.->2	n->2	
kald	j->1	
kale	r->1	
kali	e->5	g->3	s->4	
kall	 ->674	a->38	e->2	t->2	
kalp	a->1	
kalt	 ->5	,->1	.->1	
kalv	 ->1	
kaly	d->1	
kam 	f->1	o->1	
kam!	D->1	
kam,	 ->1	
kaml	i->2	
kamm	a->60	e->1	
kamp	 ->8	a->6	e->16	å->1	
kamr	a->1	
kan 	-->3	A->1	E->3	I->1	a->39	b->46	d->39	e->21	f->80	g->61	h->27	i->79	j->33	k->32	l->28	m->41	n->13	o->32	p->19	r->15	s->60	t->45	u->42	v->76	ä->9	å->12	ö->5	
kan,	 ->6	
kan.	(->1	D->3	O->1	V->2	
kana	d->2	l->9	
kand	a->9	e->360	i->15	
kane	n->6	r->11	
kani	k->1	n->1	s->9	
kano	n->1	
kans	 ->2	k->67	l->2	
kant	 ->3	,->2	.->1	e->1	
kaos	 ->2	
kap 	-->1	a->22	b->2	d->3	e->1	f->3	g->1	h->1	i->7	k->1	m->2	n->1	o->15	s->11	t->1	u->2	v->1	
kap"	 ->1	!->1	,->1	
kap,	 ->16	
kap.	 ->1	D->7	E->1	I->2	J->2	S->1	T->1	V->2	
kap:	 ->1	
kapa	 ->100	c->5	d->5	n->24	r->29	s->13	t->10	
kape	n->125	r->22	t->97	
kapi	t->25	
kapl	i->37	
kapp	 ->1	,->1	.->1	a->3	
kapr	o->1	
kaps	 ->1	-->1	a->2	b->3	d->1	f->1	i->14	k->3	l->3	m->20	n->11	o->1	p->7	r->18	s->4	å->2	
kapt	e->2	
kar 	1->1	F->1	L->1	T->1	a->13	b->4	d->18	e->8	f->14	g->1	h->6	i->15	j->1	k->11	l->2	m->12	n->2	o->10	p->3	r->8	s->18	t->2	u->4	v->16	ä->1	ö->4	
kar,	 ->8	
kar.	D->1	E->1	J->1	M->1	O->1	V->3	
kar:	 ->1	
kara	?->1	k->11	n->6	
kare	 ->30	,->9	.->2	n->13	s->3	u->1	
karg	a->1	
kark	o->2	
karl	a->1	ä->5	
karn	a->52	
karp	t->2	
karr	i->2	
kars	 ->1	
kart	a->3	e->14	l->1	
kas 	a->10	b->1	d->1	e->4	f->6	h->3	i->5	k->3	l->1	m->19	n->2	o->8	p->2	r->1	s->2	t->3	u->3	v->2	ä->4	å->1	ö->3	
kas!	H->1	
kas,	 ->10	
kas.	D->2	F->1	H->3	I->2	J->1	M->1	
kask	a->1	
kasm	u->1	
kass	e->1	o->2	
kast	 ->11	,->1	a->17	e->14	n->1	
kasu	s->3	
kaså	 ->4	
kat 	-->2	9->1	a->7	d->3	e->2	f->4	h->3	i->3	k->2	m->5	o->6	p->5	r->1	s->6	t->1	u->3	y->1	ä->1	
kat,	 ->8	
kat.	D->3	H->3	Ö->1	
kata	l->4	s->88	
kate	g->8	r->2	
kati	o->18	
kato	l->7	r->5	
kats	 ->27	,->1	.->3	?->1	
katt	 ->3	,->2	.->2	a->17	e->32	n->10	
kavi	s->4	
kay 	f->2	h->1	
kay,	 ->3	
kay.	V->1	
kayD	e->1	
kayb	e->1	
kays	 ->2	
kbar	 ->1	a->3	h->5	t->3	
kbed	ö->4	
kbes	t->4	
kbil	d->1	
kbor	r->1	
kbär	a->1	
kdam	m->1	
kdel	 ->5	,->1	.->1	e->1	
kdom	 ->1	
kdör	r->1	
ke (	f->1	
ke -	 ->4	
ke I	t->1	
ke a	g->1	n->1	t->4	
ke b	a->2	e->2	i->1	l->2	
ke d	e->4	y->1	å->1	
ke e	l->3	n->5	t->1	
ke f	i->2	r->1	ö->6	
ke g	e->4	ö->1	
ke h	a->4	
ke i	 ->11	n->10	
ke k	a->1	o->8	u->2	ä->1	
ke l	a->1	e->2	i->2	ä->2	å->1	
ke m	a->1	e->4	i->1	å->2	
ke n	a->1	i->3	
ke o	c->14	f->1	m->5	
ke p	r->3	å->45	
ke r	e->2	ö->1	
ke s	e->1	k->1	n->1	o->8	p->1	ä->2	
ke t	a->1	e->1	i->11	y->1	
ke u	n->1	t->6	
ke v	a->2	i->4	o->2	
ke ä	r->10	v->1	
ke ö	n->1	
ke!Ä	v->1	
ke) 	f->1	o->1	
ke, 	B->1	S->1	b->1	d->3	f->1	g->1	h->3	i->1	k->1	m->1	n->2	o->3	s->1	u->1	v->2	å->1	
ke-a	l->1	v->1	
ke-d	a->1	i->2	
ke-f	o->1	
ke-m	e->1	
ke-s	p->3	t->9	
ke. 	D->1	
ke.-	 ->1	
ke..	 ->1	(->1	
ke.D	e->5	ä->1	
ke.F	r->2	ö->2	
ke.H	e->1	
ke.I	 ->1	
ke.J	a->2	
ke.M	e->2	
ke.N	i->1	
ke.O	m->1	
ke.V	i->4	
ke.Ö	s->1	
ke: 	i->1	
keEn	 ->1	
keFr	u->1	
keNä	s->1	
keba	n->1	
ked 	l->1	o->1	t->1	
ked.	D->1	
keda	 ->2	n->1	t->1	
kede	 ->3	.->1	t->3	
kedj	a->3	o->1	
kedo	m->10	
kefr	i->1	
kefö	r->1	
kegå	n->1	
kekv	o->1	
kel 	-->1	1->16	2->13	3->8	4->8	5->6	6->12	7->8	8->16	9->3	a->3	b->1	f->2	k->2	n->1	o->3	s->3	ä->3	
kel,	 ->4	
kel.	E->1	T->1	V->1	Ä->1	
kel:	 ->2	
kelf	r->2	u->1	
kelm	a->1	
keln	 ->7	,->1	
kelp	r->1	
kelr	i->1	o->1	
kels	e->10	k->1	
kelt	 ->28	i->1	
kelv	ä->2	
keme	d->1	
kemi	k->5	s->2	
kemå	l->3	
kemö	j->4	
ken 	(->1	-->3	1->2	G->1	J->1	K->3	S->2	T->3	a->17	b->7	d->3	e->4	f->36	g->4	h->8	i->30	j->5	k->9	l->4	m->24	n->3	o->23	p->17	r->4	s->26	t->12	u->10	v->5	y->1	Ö->1	ä->4	å->5	ö->1	
ken,	 ->30	
ken.	 ->1	A->1	B->1	D->13	E->3	F->3	H->3	I->1	J->6	K->1	M->2	P->1	S->1	V->1	
ken:	 ->3	
ken?	F->1	J->1	V->1	
kenH	e->1	
kens	 ->30	k->9	
keom	r->2	
kepo	l->1	s->1	
kepp	 ->2	s->6	
keps	i->1	
kept	i->8	
ker 	-->1	C->1	E->1	a->41	b->10	d->23	e->5	f->11	g->4	h->7	i->28	j->16	k->5	m->19	n->7	o->20	p->34	r->6	s->28	t->7	u->7	v->9	ä->6	ö->1	
ker,	 ->13	
ker.	-->1	B->1	D->4	G->1	H->2	M->1	N->1	P->1	V->2	
ker:	 ->2	
kera	 ->2	d->3	n->1	r->18	s->1	t->3	
kere	s->1	
kerh	e->235	
keri	k->1	n->5	p->1	s->2	u->1	
kerl	i->15	
kern	 ->2	a->30	s->1	
kers	 ->2	t->24	
kert	 ->26	!->1	,->2	h->1	
kerä	g->1	t->1	
kes 	a->1	b->1	d->2	f->9	i->2	k->1	n->1	o->3	p->1	r->2	s->2	v->1	
kes-	 ->4	
kesa	r->1	
kese	k->1	t->1	
kesf	r->4	ö->1	
kesh	a->4	
kesi	s->1	
kesk	a->1	v->1	
kesl	a->2	i->2	
kesm	i->9	ä->1	
kesp	o->3	
kest	e->1	
kesu	t->7	
kesv	a->1	
ket 	(->3	-->2	B->1	E->2	G->1	P->1	V->1	a->51	b->22	d->11	e->16	f->44	g->26	h->19	i->35	j->10	k->42	l->29	m->27	n->17	o->38	p->25	r->16	s->104	t->23	u->15	v->92	ä->23	å->2	ö->1	
ket!	(->1	
ket,	 ->35	
ket.	D->2	E->2	I->1	J->1	M->2	N->1	O->1	S->1	V->1	
ket:	 ->1	
ket;	 ->3	
ket?	O->1	
kete	t->3	
keti	n->2	
ketm	a->1	
ketr	y->3	
kets	 ->14	
kett	 ->13	,->1	.->1	
keva	t->2	
kfak	t->1	
kfar	t->7	
kfor	d->1	
kfri	t->2	
kfro	n->1	
kfyl	l->1	
kför	e->8	h->1	s->1	v->1	
kgil	t->2	
kgru	n->31	p->2	
kh h	a->1	
kh-a	v->1	
kh.D	e->1	
kh.F	ö->1	
khan	t->6	
khee	r->14	
khet	 ->30	,->1	.->2	e->8	
khol	m->3	
khus	 ->1	,->2	.->1	e->2	l->1	
khäl	s->9	
ki L	i->2	
ki.D	e->1	
kick	 ->3	.->1	a->12	l->1	
kidn	a->1	
kien	 ->2	,->1	
kiet	 ->27	,->2	.->2	s->4	
kift	e->6	
kig 	s->1	
kigt	 ->4	
kild	 ->17	.->1	a->37	e->4	r->3	
kilj	a->10	e->10	t->1	
kill	i->2	n->45	
kilo	 ->3	,->1	m->1	
kilt	 ->130	
kin 	o->2	s->2	
kin.	D->1	
kine	n->2	r->1	s->9	
king	 ->1	r->3	
kinl	i->1	
kipa	 ->2	n->1	
kipn	i->9	
kire	r->1	
kis 	f->1	i->1	p->1	
kis!	 ->1	
kisb	e->1	
kisk	 ->7	a->57	e->3	
kiss	 ->1	e->3	
kist	a->12	
kit 	a->2	f->1	t->1	
kiti	n->2	
kits	 ->1	
kiv 	l->1	
kive	r->1	
kjut	a->13	e->7	i->5	s->5	v->1	
kkap	i->1	
kki 	L->2	
kkom	m->2	
kkun	n->1	s->1	
kkuy	u->2	
kköy	 ->1	
kl. 	1->17	2->3	
kl.1	2->1	
kla 	a->2	d->2	e->10	f->3	h->1	i->1	k->1	l->1	n->4	o->5	r->1	s->6	t->1	u->1	v->1	ö->1	
kla.	M->1	
klad	 ->2	e->10	
klag	a->79	e->3	l->8	o->4	
klam	 ->2	e->1	
klan	d->43	g->1	
klap	p->2	
klar	 ->25	,->4	.->2	a->83	e->3	g->17	h->12	i->24	l->5	n->12	t->97	
klas	 ->19	.->3	:->1	s->22	t->2	
klat	 ->2	,->1	s->4	
klau	s->6	
klav	e->1	
kled	 ->1	
kler	i->4	n->1	
klet	 ->1	
klib	b->1	
klie	n->1	
klig	 ->38	,->2	.->2	a->97	e->147	h->29	t->70	
klim	a->14	
klin	g->177	
kloa	k->1	
kloc	k->2	
klok	a->2	t->5	
klud	e->4	
kluk	t->1	
klus	i->20	
klyf	t->5	
klyv	e->1	
kläg	g->1	
klös	t->1	
km l	å->1	
km m	i->1	
km, 	t->1	
km.T	r->1	
kmen	i->2	
kmet	e->2	
kmod	e->1	
kna 	d->2	i->1	m->4	s->1	t->1	u->3	v->1	
kna,	 ->1	
kna.	V->1	
knad	 ->9	,->6	.->2	e->158	s->29	
knan	d->20	
knap	p->16	
knar	 ->37	
knas	 ->25	,->3	.->2	
knat	 ->11	,->1	s->7	
knee	x->1	
knel	i->1	
knes	 ->1	
knik	 ->6	e->7	
knin	g->349	
knip	a->1	p->3	
knis	k->36	
kniv	å->1	
knol	o->3	
know	-->1	
knus	s->1	
knut	e->4	n->2	p->1	
knyt	a->5	e->2	n->1	s->1	
knäc	k->2	
ko C	a->5	
ko, 	A->1	
ko.T	y->1	
koal	i->14	
kod 	f->5	h->1	k->1	
kode	n->3	r->3	
kodi	f->2	
koef	f->1	
koff	e->1	
kofi	n->2	
kofö	r->2	
kog 	e->1	f->1	i->1	
koga	r->10	
koge	n->5	
kogr	i->1	
kogs	a->2	b->6	f->1	k->1	o->1	p->1	s->4	u->1	v->1	ä->2	
kogå	r->1	
koha	n->3	
kohe	r->1	
koho	l->1	
koka	 ->1	
koko	r->1	
kol-	 ->1	
kola	 ->2	n->4	
kold	i->5	
kole	n->1	
koli	b->1	v->3	
koll	 ->6	.->3	e->222	i->3	
kolo	g->16	n->1	r->3	s->1	
kom 	-->1	a->1	d->12	e->1	f->7	h->1	i->3	l->1	m->4	n->1	o->3	p->2	r->3	s->1	t->2	u->1	v->1	ö->3	
kom,	 ->1	
kom.	D->1	
koma	n->1	
komb	i->1	
koml	i->9	
komm	a->160	e->822	i->1146	u->32	
komn	a->45	
komp	e->21	l->44	o->4	r->21	
komr	å->10	ö->6	
koms	t->18	
kon 	a->1	
kona	d->1	r->1	
konc	e->40	i->2	
konf	e->172	i->4	l->16	r->1	
kong	r->1	
konj	u->1	
konk	r->57	u->272	
kono	m->286	
kons	e->67	o->3	t->103	u->65	
kont	a->20	e->1	i->7	o->7	r->189	
konv	e->27	
koop	e->1	
kop 	b->1	
kop,	 ->3	
kopi	a->1	e->1	
kopo	u->5	
kopp	l->6	
kor 	-->1	a->2	d->4	e->1	f->21	h->3	i->13	l->2	m->3	n->1	o->6	p->1	s->25	t->5	u->2	v->3	ä->3	
kor,	 ->12	
kor.	B->1	D->4	E->1	G->1	J->1	T->1	Ö->1	
kora	n->1	
kord	 ->1	t->1	
kore	a->1	n->21	
korl	i->2	
korn	a->34	
korr	e->28	i->2	u->9	
kors	 ->15	
kort	 ->55	,->3	.->5	:->1	?->1	a->6	e->20	f->2	n->1	s->4	
kosa	m->1	
kosl	ä->1	
kost	a->9	h->1	n->104	s->2	
kosy	s->4	
koti	k->7	
kott	 ->20	,->2	.->5	e->135	l->5	s->5	
kour	i->1	
kov 	n->1	o->1	
kove	t->1	
kpar	t->10	
kpro	b->1	v->3	
kra 	a->1	d->1	e->12	f->1	g->1	h->1	i->1	k->1	m->1	o->6	p->5	s->4	v->1	ö->1	
krad	 ->1	e->2	
kraf	t->149	
kran	s->1	
krar	 ->4	.->1	e->2	n->3	
kras	.->1	c->3	s->1	t->5	
krat	 ->2	e->24	i->143	t->2	
krav	 ->39	,->4	.->6	?->1	a->1	e->40	
krea	t->3	
kred	i->2	
kreg	e->1	
kren	g->2	
krep	u->3	
krer	a->1	
kret	 ->19	:->1	a->39	e->14	i->2	s->10	
krev	 ->6	s->2	
krid	a->12	e->7	s->2	
krif	t->22	
krig	 ->6	"->1	,->1	.->1	e->12	s->2	
krik	.->1	e->39	t->4	
krim	i->27	
krin	g->55	
kris	 ->7	?->1	e->9	m->2	o->1	s->2	t->13	
krit	a->1	e->21	i->48	
kriv	a->11	b->1	e->25	i->8	n->8	s->8	
kroa	t->1	
kroe	k->5	
krof	i->1	ö->1	
krok	r->2	
krom	 ->1	,->1	a->1	
kron	j->1	
krop	p->1	
kros	s->1	t->1	
krot	.->1	a->10	f->1	n->15	
krov	 ->6	"->1	,->1	.->2	e->3	k->1	s->1	
kry.	D->1	
kryg	g->1	
kryp	h->3	t->2	
krys	s->1	
kryt	e->1	
kräc	k->9	
kräd	d->1	
kräf	t->30	
kräk	t->1	
kräm	d->1	l->1	m->3	
krän	k->29	
kräp	n->1	
krät	t->1	
kräv	a->34	d->4	e->44	s->55	t->2	
krån	g->2	
krön	a->1	
ks a	n->1	v->3	
ks b	e->2	
ks d	e->2	o->1	
ks e	f->1	
ks f	r->1	
ks g	e->1	
ks i	n->1	
ks m	i->2	å->1	
ks n	a->1	
ks o	c->5	m->1	
ks p	a->1	e->1	
ks r	e->1	
ks s	a->1	o->1	t->1	u->1	
ks t	i->2	y->1	
ks u	p->1	t->1	
ks v	a->1	e->1	i->1	
ks ö	v->1	
ks, 	d->1	
ks.D	ä->1	
ks.O	L->1	
ks.P	å->1	
ks.U	t->1	
ks.V	i->1	
ks; 	d->1	
ksak	e->1	
ksam	 ->13	.->1	h->88	m->20	t->7	
ksan	l->1	
ksbo	r->1	
ksbå	d->1	
ksce	n->1	
ksch	e->1	
ksdr	a->3	
ksek	o->1	r->1	
ksfa	l->2	
ksfo	n->1	
ksfr	å->1	
ksil	v->3	
kskö	r->1	
kslo	b->1	
kslu	t->1	
ksod	l->1	
ksom	 ->55	r->2	
kson	 ->2	
kspo	l->6	
kspr	i->1	o->2	
ksre	f->1	g->1	
ksri	s->2	
ksse	k->5	
kssy	n->1	
ksta	n->1	v->1	
ksty	r->1	
kstä	d->1	l->21	
ksva	t->1	
kswa	g->1	
ksäg	n->1	
kså 	"->1	-->2	1->1	E->3	F->1	M->1	a->73	b->28	d->25	e->32	f->43	g->18	h->26	i->37	j->1	k->33	l->2	m->38	n->13	o->11	p->18	r->6	s->48	t->31	u->18	v->35	z->1	ä->20	å->3	ö->3	
kså,	 ->10	
kså.	D->1	I->1	J->1	N->1	P->1	
ksöd	e->1	
kt (	8->2	
kt -	 ->4	,->1	
kt 1	 ->1	,->1	1->1	
kt 2	 ->2	6->1	
kt 4	 ->2	
kt 5	,->1	
kt 6	 ->1	
kt 7	 ->1	
kt D	 ->1	
kt E	U->2	u->4	
kt F	l->1	r->1	
kt K	o->1	
kt M	ü->1	
kt a	b->1	l->1	n->7	r->3	t->46	v->6	
kt b	a->2	e->17	i->12	l->3	r->1	u->1	y->2	ä->1	
kt c	h->1	i->1	
kt d	)->1	a->1	e->12	o->1	r->1	ä->4	
kt e	)->1	f->1	g->2	k->1	l->2	n->4	r->5	t->3	x->2	
kt f	a->4	e->3	i->3	l->1	r->6	u->1	y->1	ä->1	å->5	ö->56	
kt g	e->2	r->3	ä->3	å->2	ö->3	
kt h	a->17	e->1	i->1	u->4	ä->2	å->2	
kt i	 ->14	n->26	s->2	
kt j	u->1	
kt k	a->8	l->3	o->13	u->3	v->1	ä->1	
kt l	a->4	e->2	y->1	ä->4	
kt m	a->4	e->21	i->7	o->6	y->3	å->1	ö->1	
kt n	y->1	ä->5	ö->2	
kt o	c->42	m->15	p->1	r->1	
kt p	a->4	e->3	o->3	å->42	
kt r	a->1	e->3	i->1	ä->2	ö->1	
kt s	a->6	e->10	i->3	k->11	m->1	o->42	p->1	t->16	v->3	y->2	ä->18	å->1	
kt t	a->6	e->1	i->9	o->1	r->1	v->2	
kt u	n->1	p->5	r->3	t->11	
kt v	a->13	e->2	i->19	ä->3	å->1	
kt ä	m->1	n->5	r->17	v->2	
kt å	t->1	
kt ö	g->1	l->1	v->4	
kt!N	ä->1	
kt",	 ->1	
kt, 	"->1	a->1	b->1	d->2	e->5	f->3	g->1	i->1	l->1	m->8	n->2	o->6	r->1	s->4	t->2	u->2	v->4	ä->2	
kt. 	D->1	
kt.(	P->1	
kt.A	l->1	v->1	
kt.B	e->1	o->1	å->2	
kt.D	e->17	i->1	ä->1	å->1	
kt.F	e->1	ö->1	
kt.G	e->1	
kt.H	e->1	
kt.I	 ->3	
kt.J	a->6	
kt.K	o->1	
kt.M	a->4	e->1	i->1	å->1	
kt.N	u->1	å->1	
kt.O	c->1	m->3	
kt.P	r->1	
kt.R	e->1	
kt.S	l->2	
kt.T	a->1	i->1	
kt.U	n->1	
kt.V	a->3	i->2	å->1	
kt.Å	 ->1	
kt: 	J->1	V->1	d->1	u->1	
kt; 	e->1	å->1	
kt?E	u->1	
kt?T	ä->1	
kt?U	t->1	
kta 	a->8	b->12	d->6	e->7	f->4	g->2	h->1	i->3	k->5	m->3	o->4	p->4	r->7	s->14	t->1	u->7	v->2	
kta,	 ->2	
kta.	F->1	J->3	
ktab	e->2	i->1	
ktad	 ->6	.->2	e->14	m->2	
ktag	a->1	
ktai	n->2	
ktak	e->2	u->1	
ktal	a->1	
ktan	 ->5	d->6	s->7	
ktar	 ->22	,->1	.->2	e->13	n->6	
ktas	 ->18	.->1	
ktat	 ->13	,->2	.->1	o->1	s->6	u->2	
ktba	l->2	r->3	
ktbe	f->2	
ktde	l->1	
ktdi	k->1	
kte 	E->1	J->1	a->5	d->2	e->1	i->2	j->1	k->1	m->2	o->2	p->1	s->8	t->2	u->1	v->1	
kte,	 ->3	
kte.	F->1	M->1	
ktel	s->13	
kten	 ->146	,->16	.->29	s->4	
kter	 ->109	,->20	.->21	:->2	?->2	a->40	i->3	n->31	t->2	
ktes	 ->5	
ktet	 ->14	,->1	s->1	
ktfa	r->1	
ktfö	r->2	
ktha	v->1	
kthe	t->1	
kthå	l->1	
ktie	b->1	ä->2	
ktig	 ->86	,->7	.->11	?->1	a->153	h->65	t->168	
ktik	 ->1	,->1	e->10	
ktin	g->14	n->1	v->1	
ktio	n->124	
ktis	k->74	
ktiv	 ->121	,->15	.->14	:->2	?->2	a->56	e->110	f->3	i->40	t->52	
ktko	n->1	
ktli	g->18	n->74	
ktlö	s->3	
ktme	d->2	
ktmi	s->1	
ktni	n->55	
ktob	e->8	
ktor	 ->14	,->5	.->5	a->18	e->33	h->1	i->7	n->49	p->1	s->4	
ktpu	n->2	
ktra	 ->1	
ktri	c->1	
ktro	n->9	
ktru	m->2	
kts 	a->1	e->2	i->1	l->1	o->2	u->3	ö->1	
kts!	F->1	
ktsa	n->3	
ktsb	a->1	
ktsf	o->1	ö->3	
ktsm	e->1	
ktsp	l->1	r->1	
ktta	 ->3	g->1	r->1	s->3	
ktua	l->1	
ktue	l->34	
ktum	 ->64	,->1	.->2	e->1	
ktur	 ->15	,->4	.->3	b->1	e->52	f->58	m->1	n->1	p->12	r->1	s->3	u->2	å->1	
ktyg	 ->6	?->1	s->1	
ktyr	.->1	
ktär	 ->4	,->1	.->1	e->3	
ktör	 ->1	,->1	e->20	s->1	
kubi	k->2	
kugg	a->2	b->1	
kula	 ->1	.->1	t->5	
kuld	a->1	b->1	e->1	
kule	r->2	
kuli	s->1	
kull	 ->13	,->2	.->3	e->486	k->1	
kulo	r->1	
kult	u->121	
kulä	r->1	
kume	n->46	
kumu	l->2	
kund	,->1	e->30	v->1	ä->1	
kung	a->15	
kunn	a->255	i->6	
kuns	k->17	
kupa	n->1	t->1	
kupe	r->3	
kupp	g->1	
kur 	f->1	
kura	r->1	
kurr	e->285	
kurs	 ->4	,->1	.->1	e->10	ä->1	
kus 	f->1	s->1	
kus.	D->1	
kuse	r->3	
kuss	i->61	
kust	 ->1	b->1	e->20	l->2	m->3	o->2	r->1	v->1	
kuta	 ->2	b->3	n->2	
kute	r->78	
kuum	 ->1	t->1	
kuyu	 ->2	
kva,	 ->1	
kval	d->2	i->51	
kvan	t->7	
kvar	 ->19	,->2	.->2	;->1	h->3	s->8	
kvat	 ->3	a->2	i->1	
kven	s->46	t->16	
kves	t->3	
kvic	k->3	
kvid	d->3	
kvin	n->59	
kvis	t->1	
kvot	 ->4	!->1	,->1	e->10	
kväl	 ->4	l->10	
kväm	l->15	t->1	
kvär	d->11	t->7	
kväv	a->2	
kvår	d->3	
ky f	ö->1	
kydd	 ->34	)->1	,->3	.->6	a->31	e->18	s->16	
kyfa	l->1	
kyhö	g->1	
kyla	.->1	n->1	
kyld	i->29	
kyli	g->1	
kyll	a->3	e->1	s->1	
kymm	e->6	
kymr	a->10	
kymt	s->1	
kynd	a->11	s->4	
kyrk	o->1	
kyvä	r->1	
käl 	-->2	6->1	a->2	b->1	d->1	e->1	f->4	h->3	i->4	n->1	o->2	s->6	t->5	ä->2	
käl,	 ->1	
käl.	A->1	D->1	F->1	J->1	
käle	n->3	t->9	
käli	g->1	
käll	a->8	o->39	
kämd	a->1	
kämm	a->2	
kämn	e->1	
kämp	a->34	n->12	
kämt	s->1	
känd	 ->5	,->2	.->1	a->12	e->20	
känk	a->2	
känn	a->69	e->78	s->4	
käns	l->43	
känt	 ->19	,->2	s->8	
kär 	n->1	p->1	
kära	 ->53	
käre	 ->1	
kärl	 ->1	e->2	
kärn	a->4	e->8	f->2	i->3	k->21	p->4	s->4	t->2	v->8	
kärp	a->8	n->1	t->2	
kärs	 ->1	
kåda	d->2	r->1	
kådl	i->6	
kådn	i->1	
kåle	n->1	
kår,	 ->1	
kåt 	i->2	
kåts	t->1	
köks	b->1	
köl 	n->1	
köl,	 ->1	
köla	r->1	
köld	b->1	g->1	
köne	n->3	
könh	e->1	
köns	g->1	k->5	
köp 	a->2	
köpa	r->4	
köpe	r->1	
köpk	r->1	
köps	b->1	l->1	
köpt	 ->1	
kör 	ö->1	
kör.	K->1	
köra	 ->3	s->1	
körd	 ->1	a->1	e->1	
körn	i->2	
körs	 ->2	p->1	
kört	 ->3	
köt 	9->1	l->1	
köta	 ->6	s->1	
köte	r->1	
köts	 ->2	.->1	e->5	
kött	 ->5	e->2	k->1	s->3	
kövl	a->1	
köy 	-->1	
l "M	i->1	
l (B	r->1	
l (k	o->2	
l - 	d->3	f->1	n->2	o->1	r->1	s->2	u->2	ö->1	
l -,	 ->1	
l 1 	i->1	o->2	u->1	
l 1,	 ->2	
l 1-	o->4	r->5	s->2	
l 1.	J->1	
l 10	 ->1	5->1	
l 11	0->1	
l 12	 ->1	,->1	
l 13	 ->4	.->1	
l 14	3->1	
l 15	 ->1	8->3	
l 16	)->1	
l 19	3->1	5->1	9->2	
l 2 	-->1	0->1	b->1	e->1	o->1	s->1	
l 2,	 ->1	4->1	6->1	
l 2-	o->2	s->1	
l 2.	1->1	2->1	M->1	
l 22	6->1	
l 25	 ->1	5->4	
l 28	0->5	
l 29	9->2	
l 3 	0->1	
l 3.	1->1	8->1	
l 30	 ->2	
l 33	 ->2	
l 37	 ->1	.->1	
l 39	 ->1	
l 4 	c->1	i->4	p->1	
l 4.	2->1	
l 42	 ->1	
l 48	 ->2	
l 5 	g->1	
l 5.	4->1	
l 50	 ->2	,->1	
l 52	 ->1	
l 56	,->1	
l 5b	 ->1	.->1	
l 6 	i->6	o->3	
l 6,	 ->1	
l 6.	S->1	
l 62	 ->1	
l 67	 ->1	
l 7 	i->6	n->1	
l 7,	 ->1	4->1	
l 70	0->1	
l 75	 ->1	
l 77	 ->1	
l 81	 ->1	.->9	
l 82	,->1	.->1	
l 83	 ->1	
l 85	 ->1	
l 87	.->2	
l 88	 ->2	
l 9 	m->1	
l 9.	1->1	
l 91	 ->1	
l 94	 ->2	,->1	
l 95	 ->1	
l Al	b->1	
l Ba	r->1	s->1	
l Bo	u->2	
l Br	y->2	
l Ch	i->1	
l Co	n->1	u->1	
l De	n->1	
l Di	m->1	
l EG	 ->1	-->2	
l EU	 ->2	-->1	.->1	:->2	
l Ef	t->1	
l Eu	r->25	
l Fr	a->3	
l Fö	r->4	
l Ge	n->1	
l Gr	e->1	
l He	i->1	
l Hi	l->1	
l In	t->2	
l Ir	l->1	
l Ka	n->1	r->1	u->1	
l Ki	n->1	r->2	
l Ko	s->9	u->1	
l Ku	l->1	
l Lo	r->2	
l Mc	N->1	
l Mi	c->1	
l Mo	r->2	
l Ni	e->2	
l Ny	a->1	
l OL	F->1	
l PP	E->1	
l Pa	l->1	t->2	
l Pe	a->1	
l Po	l->1	
l Pu	r->1	
l Ra	p->1	
l Ri	o->1	
l Sc	h->1	
l Sh	e->1	
l So	l->3	
l St	.->1	r->1	
l Sy	r->1	
l Th	e->1	
l Ti	b->1	
l Tr	e->1	
l Ty	s->2	
l Ul	s->1	
l Ve	r->1	
l Wa	l->1	s->1	
l Wi	l->1	
l Wu	r->1	
l ab	s->1	
l ac	c->1	
l ag	e->1	
l al	d->2	l->35	
l an	d->5	f->1	g->1	l->1	m->2	n->1	p->1	s->12	t->3	v->11	
l ap	p->1	
l ar	b->8	m->1	t->5	
l at	t->300	
l av	 ->132	,->1	g->2	k->1	l->1	m->1	s->9	t->2	v->3	
l ba	c->1	g->1	l->1	n->2	r->11	s->1	
l be	 ->6	d->5	f->4	g->7	h->10	k->1	m->1	r->5	s->13	t->37	v->5	
l bi	b->3	d->5	l->5	
l bl	a->1	i->23	o->2	
l bo	r->3	t->3	
l br	a->1	i->2	o->1	ä->1	ö->1	
l bu	d->1	
l by	g->2	
l bä	r->3	s->1	t->2	
l bå	d->2	
l bö	d->1	r->13	
l ca	 ->1	
l ce	n->1	
l ci	t->2	
l co	r->1	
l da	g->1	
l de	 ->71	b->4	c->1	f->1	l->15	m->11	n->90	r->5	s->13	t->88	
l di	a->3	r->17	s->8	
l do	c->2	m->2	
l dr	a->2	i->1	y->1	
l du	m->3	
l dä	r->17	
l då	 ->3	?->1	
l ef	f->2	t->4	
l eg	e->3	
l ek	o->3	
l el	l->7	
l em	e->2	i->1	
l en	 ->108	b->1	d->3	e->2	k->1	l->1	t->1	
l er	 ->3	,->4	:->1	b->1	f->1	h->1	i->2	s->1	t->1	
l et	t->32	
l eu	r->3	
l ex	e->45	i->1	
l fa	l->3	m->1	r->1	s->2	t->7	
l fe	b->1	l->2	
l fi	c->1	n->6	s->1	
l fl	e->1	y->2	
l fo	n->3	r->10	
l fr	a->10	e->2	i->4	u->1	ä->8	å->31	
l fu	l->5	n->9	
l fy	l->2	
l fä	r->1	s->1	
l få	 ->10	n->1	r->2	
l fö	l->24	r->198	
l ga	g->3	m->2	n->1	r->2	
l ge	 ->10	m->8	n->17	s->2	t->1	
l gi	s->1	
l gl	ä->1	
l go	d->10	
l gr	a->8	u->13	
l gä	l->8	r->7	
l gå	 ->10	.->1	n->2	
l gö	r->25	
l ha	 ->39	.->1	m->1	n->22	r->17	v->14	
l he	d->1	l->4	m->2	n->1	r->4	
l hi	n->5	
l hj	ä->6	
l ho	n->1	p->1	
l hu	m->1	r->5	
l hy	c->1	
l hä	l->1	n->3	r->5	
l hå	l->2	
l hö	g->4	r->3	
l i 	1->1	A->1	D->1	E->4	F->1	M->1	V->1	a->6	d->16	e->2	f->8	g->3	i->1	k->1	l->2	m->5	n->1	o->2	p->1	s->9	t->1	u->2	v->7	ä->1	
l ic	k->1	
l id	é->1	
l in	 ->1	b->2	d->5	f->7	g->4	l->5	n->3	o->9	r->5	s->7	t->60	v->1	ö->1	
l is	r->1	
l ja	g->108	n->1	
l jo	r->1	
l ju	 ->4	l->1	s->1	
l jä	m->2	
l ka	l->1	m->3	n->13	s->1	t->1	
l kl	a->4	
l kn	y->1	
l ko	d->1	l->5	m->56	n->22	r->3	s->1	
l kr	a->1	i->3	ä->2	
l ku	l->1	n->57	
l kv	e->1	i->4	ä->1	
l kä	n->1	r->2	
l kö	k->1	
l la	g->1	n->2	
l le	d->5	t->1	
l li	g->7	k->2	v->5	
l lu	c->1	
l ly	c->3	d->1	f->1	s->2	
l lä	g->4	m->6	n->2	r->1	s->1	t->2	
l lå	t->3	
l lö	p->1	s->2	
l ma	j->2	k->5	n->11	r->5	
l me	d->46	l->10	n->2	r->4	t->1	
l mi	d->1	g->3	l->1	n->18	s->1	t->2	
l mo	b->1	t->6	
l mu	s->1	
l my	c->5	n->3	
l mä	n->1	r->1	
l må	l->3	n->6	s->7	
l mö	j->4	t->2	
l na	c->4	t->10	
l ni	 ->5	v->11	
l no	g->1	r->1	
l nu	 ->4	
l ny	 ->2	a->4	l->1	t->6	
l nä	m->4	r->10	s->4	
l nå	 ->1	g->11	
l nö	d->2	
l oa	c->1	
l oc	h->127	k->27	
l oe	n->1	
l of	f->2	ö->1	
l oi	g->1	
l oj	ä->1	
l ol	i->3	y->3	
l om	 ->30	,->1	f->9	l->1	r->4	s->2	v->2	
l op	t->1	
l or	d->3	g->2	o->3	ä->1	
l os	s->4	
l oä	n->2	
l pa	r->10	s->1	
l pe	l->1	n->4	r->6	
l pi	l->1	
l pl	a->5	
l po	l->6	s->2	
l pr	a->1	e->7	i->7	o->9	
l pu	n->2	
l på	 ->35	,->1	.->1	l->1	m->1	p->3	s->2	t->1	v->1	
l ra	d->1	m->2	t->1	
l re	d->6	f->1	g->14	k->4	p->1	s->11	t->1	v->2	
l ri	k->5	s->2	
l ro	l->4	
l ry	m->1	
l rä	c->4	k->1	t->18	
l rå	d->20	
l rö	r->3	s->1	
l sa	k->4	m->19	n->1	t->1	
l se	 ->15	r->1	s->2	t->1	
l si	g->4	m->1	n->14	s->12	t->9	
l sj	ä->3	ö->4	
l sk	a->17	e->4	i->5	j->2	o->3	r->1	u->6	y->7	ö->2	
l sl	u->15	å->2	
l sm	å->2	
l sn	a->1	
l so	c->4	l->3	m->105	
l sp	e->3	ä->1	
l st	a->9	e->1	i->1	o->13	r->6	y->1	ä->5	å->42	ö->3	
l su	b->4	s->1	v->1	
l sv	a->3	å->1	
l sy	n->2	s->5	
l sä	g->39	k->10	n->2	r->4	t->2	
l så	 ->4	d->2	
l sö	r->1	
l ta	 ->17	c->21	l->12	s->3	
l te	n->1	r->1	x->1	
l ti	d->3	l->40	t->2	
l to	l->2	t->1	
l tr	a->2	e->4	o->5	y->3	ä->4	
l tu	r->1	
l tv	i->1	ä->1	å->6	
l ty	c->2	d->1	
l tä	c->1	n->1	
l u-	l->1	
l un	d->16	i->3	
l up	p->24	
l ur	 ->4	s->1	v->1	
l ut	a->9	b->2	f->7	g->3	n->1	o->1	r->2	s->12	t->8	v->10	ö->2	
l va	d->10	l->1	n->1	p->1	r->47	
l ve	r->15	t->9	
l vi	 ->40	a->1	c->1	d->10	k->1	l->7	s->11	
l vo	l->1	n->3	r->2	
l vä	g->1	l->2	n->2	r->1	s->1	
l vå	r->16	
l yr	k->2	
l yt	t->3	
l Ös	t->1	
l äg	n->1	
l än	 ->8	d->15	
l är	 ->40	?->1	
l äv	e->6	
l åk	l->2	
l år	 ->2	
l ås	i->1	t->2	
l åt	 ->1	a->2	e->14	g->3	s->1	t->1	
l ök	a->5	n->1	
l ön	s->1	
l öp	p->3	
l ös	t->1	
l öv	e->20	
l! I	n->1	
l! J	a->1	
l!He	r->1	
l!Hä	r->1	
l!Ja	g->1	
l!Me	n->1	
l!Ti	l->1	
l" m	e->1	
l" o	c->1	
l", 	s->1	v->1	
l".I	 ->1	
l'ea	u->1	
l, A	n->1	
l, R	e->1	
l, T	y->1	
l, a	n->1	t->5	v->2	
l, b	e->1	
l, d	e->4	i->1	v->1	ä->2	å->1	
l, e	f->3	l->2	r->1	t->2	u->1	
l, f	o->1	r->2	ö->5	
l, g	e->1	r->1	
l, h	a->4	u->1	ä->1	
l, i	 ->7	n->1	
l, j	a->1	u->2	
l, k	a->1	o->3	u->1	
l, l	a->1	i->1	ä->1	
l, m	e->19	o->1	
l, n	a->1	i->1	ä->5	å->2	
l, o	c->30	m->2	
l, p	o->1	r->1	å->1	
l, r	e->1	ä->1	ö->1	
l, s	i->1	o->15	å->6	ö->1	
l, t	i->1	o->2	å->1	
l, u	n->1	t->4	
l, v	a->4	i->7	
l, ä	n->1	v->3	
l, å	n->1	t->2	
l, ö	v->1	
l- o	c->18	
l-2-	o->1	
l-De	l->1	
l-Fi	n->3	
l-He	i->1	
l-I)	;->1	
l-II	)->1	
l-Ro	b->1	
l-Sh	a->1	e->5	
l-Sy	r->1	
l-fö	r->1	
l-pr	o->1	
l-so	c->2	
l. 1	1->6	2->6	3->1	5->2	7->1	9->1	
l. 2	0->1	1->2	
l. D	e->1	
l. E	n->1	
l. J	a->1	
l. o	c->1	
l.12	.->1	
l.Al	l->1	
l.An	g->1	
l.Av	s->1	
l.Be	t->1	
l.Bi	l->1	
l.Bä	s->1	
l.De	 ->2	n->7	s->1	t->34	
l.Dä	r->3	
l.EU	-->1	
l.Ef	t->1	
l.En	l->3	
l.Et	t->3	
l.Eu	r->2	
l.Fi	n->2	
l.Fr	a->1	u->3	å->1	
l.Fö	r->8	
l.Ge	n->1	
l.Ha	r->1	
l.He	r->8	
l.Hu	r->1	
l.Hä	r->1	
l.I 	A->1	d->1	e->1	f->2	o->1	s->1	u->1	
l.In	g->1	t->1	
l.Ja	 ->1	g->21	
l.Ka	n->1	
l.Ko	m->3	s->1	
l.Ku	l->1	
l.Kä	r->1	
l.Ly	n->1	
l.Ma	r->1	
l.Me	d->1	n->8	
l.Mi	n->1	
l.Må	l->1	
l.Nä	r->4	
l.Om	 ->1	
l.Or	k->1	
l.Pe	r->1	
l.Pr	o->1	
l.På	 ->1	
l.Re	s->1	
l.Sa	m->3	n->1	
l.Sc	h->1	
l.Sj	ä->1	
l.Sm	å->1	
l.So	m->1	
l.St	r->1	
l.Så	 ->3	s->1	
l.Ta	n->1	
l.Tr	o->1	
l.Tv	å->1	
l.Tä	n->1	
l.Ut	m->1	
l.Vi	 ->23	
l.Vo	n->1	
l.Vå	r->1	
l.a.	 ->27	
l.Än	 ->1	d->1	
l.Är	 ->1	
l.Äv	e->1	
l: "	h->1	
l: E	u->1	
l: F	i->1	
l: O	s->1	
l: U	n->1	
l: V	e->1	i->1	
l: a	t->1	
l: d	e->1	
l: e	n->1	
l: j	a->1	
l: p	r->1	
l; a	t->1	
l; f	ö->1	
l; i	 ->1	
l?. 	(->1	
l?Da	g->1	
l?El	l->1	
l?Hu	r->1	
l?Ja	g->2	
l?Ko	l->1	
lFin	a->1	
la -	 ->2	
la 9	0->1	
la A	l->1	
la B	a->1	
la E	U->4	u->20	
la F	ö->1	
la H	i->1	
la K	o->2	
la L	o->1	
la M	e->1	
la P	a->1	
la S	u->1	
la U	C->1	
la a	g->1	k->3	l->5	n->16	r->5	s->9	t->32	v->16	
la b	a->3	e->30	i->14	l->2	o->4	r->3	u->2	ö->3	
la d	e->133	i->17	o->6	r->1	ö->1	
la e	f->2	g->2	k->7	l->10	m->2	n->37	r->9	t->8	u->7	v->2	x->1	
la f	a->26	i->4	l->2	o->17	r->33	u->1	å->2	ö->43	
la g	e->6	i->2	l->1	o->3	r->13	å->1	
la h	a->19	e->1	i->2	j->2	o->5	u->3	ä->1	å->1	ö->5	
la i	 ->10	d->5	g->1	n->41	s->1	
la j	o->3	u->2	ä->2	
la k	a->9	l->5	n->2	o->47	r->6	v->3	ä->1	ö->1	
la l	a->6	e->5	i->7	o->1	ä->7	ö->4	
la m	a->11	e->40	i->16	o->4	u->1	y->32	ä->3	å->4	ö->5	
la n	a->1	e->2	i->9	o->2	u->1	y->3	ä->4	å->1	ö->1	
la o	b->3	c->61	d->1	f->1	j->1	l->5	m->72	p->3	r->7	s->5	
la p	a->24	e->3	l->2	o->15	r->23	u->1	å->7	
la r	a->4	e->35	i->3	o->1	u->1	ä->16	ö->3	
la s	a->24	e->3	i->42	j->5	k->27	l->4	n->1	o->17	p->6	t->29	u->2	v->1	y->8	ä->5	å->4	
la t	a->3	e->3	i->20	j->11	o->3	r->10	y->2	ä->1	
la u	n->11	p->11	r->1	t->31	
la v	a->6	e->10	i->13	ä->11	å->10	
la ä	n->4	r->5	
la å	 ->1	k->2	r->2	s->1	t->10	
la ö	n->1	p->1	s->1	v->5	
la!H	e->1	
la" 	s->1	v->1	
la".	B->1	H->1	
la";	 ->1	
la, 	a->1	c->1	d->1	f->1	h->2	i->2	k->1	l->1	m->1	n->2	o->3	p->1	r->2	s->3	v->1	ä->1	
la.B	i->1	
la.D	e->11	ä->1	
la.H	e->2	
la.I	 ->1	
la.J	a->3	
la.K	o->1	
la.M	e->2	
la.N	ä->1	
la.S	m->1	
la.V	i->4	
la.Ö	v->1	
la:F	ö->1	
la?A	v->1	
la?D	e->3	
laam	s->1	
labo	r->3	
lace	r->17	
laci	o->15	
lad 	a->12	e->1	f->2	h->1	i->1	l->1	m->2	o->1	p->1	r->2	s->2	ö->4	
lad,	 ->1	
lada	 ->3	k->1	
ladd	a->1	e->2	
lade	 ->83	s->17	
lafr	a->1	
lag 	-->2	1->18	2->7	3->5	4->8	5->2	6->2	a->14	b->9	d->3	e->4	f->35	g->7	h->15	i->23	j->1	k->7	l->1	m->3	n->4	o->35	p->2	r->3	s->64	t->60	u->2	v->5	ä->4	å->1	ö->1	
lag,	 ->40	
lag.	 ->1	)->3	.->1	B->1	D->9	F->5	H->4	I->2	J->6	K->1	L->1	M->2	P->1	S->1	T->1	U->1	V->4	
lag;	 ->1	
lag?	D->1	F->2	
laga	 ->8	!->1	.->2	d->2	n->10	r->73	t->1	
lagd	 ->4	,->1	a->7	
lage	l->3	n->83	r->2	t->71	
lagf	ö->5	
lagg	 ->6	,->7	.->5	;->1	a->5	e->2	n->1	o->1	
lagi	t->16	
lagl	i->18	
lagn	a->16	i->17	
lago	m->4	r->5	s->1	
lagr	a->2	e->1	
lags	 ->15	d->1	f->1	k->1	t->128	
lagt	 ->46	,->1	e->2	s->26	
lai 	L->7	
lak 	s->1	
lakt	a->1	i->24	
lam 	f->2	l->1	
lam,	 ->1	
lame	n->600	r->2	
lamo	d->2	
lamp	o->1	
lams	k->4	
lamt	 ->1	
lan 	1->6	8->2	C->2	D->1	E->10	G->1	H->1	I->9	P->3	S->3	a->5	b->2	c->1	d->32	e->8	f->20	g->2	h->2	i->1	k->18	l->6	m->16	n->4	o->9	p->8	r->19	s->15	t->2	u->8	v->7	Ö->1	ä->2	
lan"	 ->1	.->1	
lan,	 ->6	
lan.	 ->1	D->2	E->1	I->2	J->1	S->1	U->1	V->1	
lan:	 ->1	
lan?	H->1	
lanN	ä->1	
lana	 ->2	,->2	
lanc	a->1	
land	 ->196	)->1	,->31	.->29	a->18	e->286	n->10	s->69	v->2	
lane	n->13	r->85	t->3	
lang	,->1	e->7	
lanh	ö->4	
lank	e->1	l->1	o->1	t->1	
lanl	i->1	
lann	i->1	
lans	 ->16	,->2	e->22	l->1	t->7	v->1	å->1	ö->1	
lant	a->1	e->7	i->2	k->1	l->1	o->1	
lanö	s->19	
lapp	a->1	h->3	j->1	s->1	v->2	
lar 	"->1	-->4	2->1	a->25	b->4	d->31	e->7	f->24	g->2	h->6	i->30	j->4	k->4	l->2	m->26	n->6	o->114	p->10	r->5	s->39	t->6	u->7	v->10	ä->8	å->1	
lar,	 ->30	
lar.	B->1	D->10	E->1	F->2	I->4	J->7	K->1	M->2	V->4	
lar:	 ->1	
lar;	 ->1	
lar?	K->1	N->1	
lara	 ->36	,->1	.->2	d->5	r->29	s->5	t->5	
larb	e->1	
lare	 ->32	,->8	.->3	n->14	
larf	o->1	ä->1	
larg	ö->17	
larh	e->12	
lari	n->24	s->3	
larl	a->3	ä->2	
larm	r->2	s->2	
larn	 ->2	a->60	
lars	 ->2	t->1	
lart	 ->86	,->2	.->1	:->1	e->7	i->2	
larv	e->1	
lary	 ->1	
las 	a->7	b->1	d->3	e->10	h->1	i->16	k->2	l->1	m->3	n->2	o->11	p->9	s->6	t->9	u->8	v->4	y->2	ö->1	
las,	 ->8	
las.	B->1	D->4	K->2	T->1	
las:	 ->1	
lash	u->1	
lasi	a->2	e->4	
lasp	e->1	
lass	 ->2	a->1	e->3	i->15	p->1	
last	 ->5	!->1	,->2	-->1	.->1	a->6	e->6	i->1	n->6	
lat 	"->2	B->1	a->9	d->3	e->5	f->5	g->3	h->3	i->4	k->1	m->1	n->2	o->9	p->1	s->4	u->3	v->1	ö->1	
lat,	 ->5	
lat.	H->1	I->1	V->1	
late	r->14	
lath	 ->3	,->1	
lati	o->19	v->15	
latl	a->1	
lato	n->1	r->2	
lats	 ->35	,->7	.->4	e->19	
latt	a->1	
laud	e->1	
laus	u->6	
laut	r->2	
lava	n->2	r->2	
lave	r->1	
lavi	e->1	
lavt	a->1	
law,	 ->1	
law.	M->1	
laya	b->1	
laye	d->2	
lbac	è->1	
lbak	a->51	s->1	
lban	 ->1	e->5	i->1	k->8	s->4	
lbar	 ->20	a->6	h->2	t->19	
lbef	o->2	
lbel	o->1	
lber	t->1	ä->1	
lbes	 ->2	l->1	t->5	
lbil	d->1	
lblo	c->1	
lbor	d->3	
lbra	n->1	
lbri	g->1	n->4	
lbro	t->1	
lbun	d->15	
lbyr	å->1	
ld W	i->1	
ld a	v->3	
ld b	e->3	o->1	
ld f	r->5	u->1	
ld i	 ->2	n->2	
ld k	l->1	o->2	u->1	
ld m	a->1	e->1	i->1	
ld o	c->2	
ld p	a->1	e->1	o->1	u->1	å->1	
ld r	e->2	o->1	
ld s	o->1	
ld t	a->1	i->1	o->1	
ld u	p->2	
ld ä	r->1	
ld å	t->1	
ld, 	d->2	k->1	m->3	o->3	s->1	
ld.D	e->1	
ld.F	ö->1	
ld.J	a->2	
ld.N	u->1	
lda 	b->1	d->3	e->4	f->9	i->6	k->2	l->2	m->7	n->1	o->2	p->5	r->6	s->10	t->4	v->2	ä->1	å->3	
lda,	 ->5	
lda.	D->1	E->1	H->1	J->2	Ä->1	
lda?	F->1	
ldad	e->3	
ldag	e->1	
ldan	d->6	
ldar	 ->6	
ldas	 ->6	,->1	.->1	?->1	t->1	
ldat	 ->1	e->2	s->2	
ldbe	l->1	s->1	
lde 	B->1	K->1	a->1	d->5	e->4	f->4	h->1	j->1	m->1	n->2	o->1	t->1	u->1	å->1	
lde,	 ->1	
lde.	E->1	
ldel	a->13	e->23	n->3	t->3	
ldem	o->16	
lden	 ->27	,->9	.->4	:->1	?->1	s->4	
lder	 ->7	.->3	d->2	n->3	
ldes	 ->11	.->1	
ldet	 ->1	,->1	
ldez	,->1	-->2	
ldgr	ä->1	
ldhe	t->23	
ldig	 ->3	a->14	e->1	h->15	t->21	
ldio	x->5	
ldir	e->17	
ldis	t->1	
ldju	r->1	
ldni	n->66	
ldom	s->1	
ldra	 ->3	d->3	g->1	r->1	t->2	
ldre	 ->5	,->1	.->1	
ldri	g->32	
ldsa	m->3	
ldsd	e->1	
ldse	k->1	
ldsf	r->1	
ldsh	a->6	
ldsk	r->6	
ldsl	i->1	
ldsm	a->1	
ldsn	i->1	
ldso	m->1	
ldsu	t->1	
ldta	 ->1	g->1	
le -	 ->1	
le E	u->3	
le K	i->1	
le a	l->3	n->3	t->18	v->1	
le b	a->3	e->9	i->1	l->5	é->1	ö->2	
le d	e->28	o->3	ä->8	å->2	
le e	l->1	m->1	n->5	v->1	
le f	a->1	i->2	r->4	å->4	ö->20	
le g	e->2	o->1	r->1	ä->7	å->1	ö->5	
le h	a->18	e->1	ä->4	
le i	 ->6	n->20	
le j	a->44	
le k	a->1	o->6	r->2	u->56	ä->1	
le l	e->4	ä->1	
le m	a->2	e->2	o->1	
le n	a->1	i->1	u->1	ä->1	
le o	c->12	f->1	l->1	
le p	a->3	l->1	o->1	å->2	
le r	e->2	ä->1	å->1	ö->1	
le s	a->1	e->1	j->1	k->5	l->2	o->4	p->1	t->3	v->1	ä->4	å->6	ö->1	
le t	.->1	a->5	i->5	r->1	v->2	
le u	n->3	p->4	r->3	t->6	
le v	a->37	e->2	i->81	ä->3	
le ä	n->1	r->2	v->1	
le å	t->2	
le ö	n->2	
le, 	o->3	
le-d	e->2	
le.J	a->1	
le.V	i->1	
led 	i->1	m->1	
leda	 ->57	,->1	m->154	n->14	r->14	s->6	
ledd	a->3	e->20	
lede	r->40	s->44	
ledi	g->1	
ledn	i->74	
leds	 ->5	e->2	t->2	
lefa	n->1	
lefo	n->1	
lega	 ->36	!->4	,->3	.->1	d->2	l->22	n->16	s->2	t->19	
lege	.->1	?->1	r->131	
legi	e->5	t->18	u->3	
lego	r->4	
leha	n->3	
leid	o->2	
lejd	a->1	o->1	
leka	s->1	
leke	n->2	r->1	
leko	m->3	n->4	
leks	a->1	
lekt	e->3	i->16	r->10	u->3	y->1	
lele	r->3	
lell	a->2	t->3	
lels	e->9	
lem 	-->1	a->2	d->2	e->3	f->3	h->3	i->13	k->2	m->12	n->4	o->7	p->1	s->17	u->1	v->3	ä->4	ö->1	
lem,	 ->14	
lem.	 ->1	.->1	A->1	D->6	F->1	H->2	I->1	J->3	M->1	P->1	S->2	V->3	
lem:	 ->1	
lem;	 ->2	
lem?	M->1	
lema	t->5	
leme	n->37	t->48	
lemi	k->1	
leml	ä->1	
lemm	a->17	
lemo	m->3	
lems	k->2	l->36	r->1	s->284	
len 	B->1	E->1	a->27	b->7	d->3	e->4	f->16	g->2	h->8	i->33	k->5	m->9	n->2	o->13	p->2	s->18	t->6	u->6	v->3	ä->4	å->3	ö->1	
len"	 ->2	,->1	
len,	 ->32	
len.	 ->1	A->1	D->10	E->1	H->3	I->2	J->3	K->3	M->5	R->1	S->2	T->1	U->1	V->4	
len?	Ä->1	
lenF	r->2	
lena	 ->4	,->1	r->5	
lenn	i->7	
lens	 ->11	k->1	
lent	i->1	
lenu	m->5	
lenÄ	r->1	
lenä	t->1	
leot	e->1	
ler 	-->3	2->1	7->1	8->1	9->1	A->3	D->1	E->8	F->4	I->1	J->1	L->1	M->1	N->1	P->2	R->2	S->5	T->3	U->2	a->73	b->31	c->2	d->114	e->66	f->98	g->22	h->21	i->70	j->5	k->44	l->23	m->66	n->20	o->61	p->42	r->16	s->86	t->32	u->20	v->37	Ö->2	ä->21	å->8	ö->7	
ler,	 ->20	
ler-	r->1	
ler.	A->1	D->6	E->1	F->3	H->2	J->3	K->1	M->2	O->1	R->1	Ä->1	
ler;	 ->1	
ler?	P->1	
lera	 ->119	"->1	,->1	.->1	d->12	n->12	r->20	s->21	t->10	
lere	r->7	
leri	 ->4	e->1	n->25	
lerk	ä->3	
lerm	o->1	
lern	a->52	
lers	 ->2	t->1	u->3	
lert	a->6	i->67	
lerå	r->12	
les 	G->1	a->2	e->2	f->8	h->2	i->1	j->1	k->1	n->4	p->1	r->6	s->6	t->1	u->2	
les.	H->1	V->1	
les;	 ->1	
lesa	 ->1	m->5	r->1	
lese	 ->1	
lesk	a->1	
lesm	a->1	ä->1	
lesn	å->4	
lest	a->25	i->22	
lesä	t->2	
let 	-->1	A->1	E->1	T->1	V->2	a->15	b->4	d->3	e->7	f->41	g->4	h->11	i->26	j->1	k->6	l->3	m->22	n->2	o->20	p->1	r->6	s->14	t->14	u->2	v->6	Ö->1	ä->10	å->1	ö->1	
let!	P->1	
let,	 ->31	
let.	 ->1	)->1	A->2	D->11	F->1	H->2	I->2	J->7	K->1	N->1	O->1	S->2	T->1	U->1	V->4	
let:	 ->1	
leta	r->1	
lets	 ->6	
lett	 ->14	e->13	s->10	
leum	 ->1	
leur	o->3	
lev 	a->3	d->2	f->2	i->2	k->1	o->3	t->1	u->1	
leva	 ->17	,->1	?->1	n->12	
levd	e->2	
leve	b->1	l->2	r->20	
levi	s->1	
levn	a->12	
levs	 ->3	
levt	 ->4	
lewo	o->2	
lex 	f->1	
lex.	J->1	
lexa	,->1	n->2	
lexi	b->27	
lext	 ->1	
lez 	o->1	
lf H	i->2	
lf-M	a->2	
lfab	e->1	
lfed	e->1	
lfen	 ->2	.->2	
lfer	i->1	
lfin	g->1	
lfkr	i->1	
lfog	a->6	
lfon	d->15	
lfor	d->3	
lfra	m->3	
lfre	d->27	
lfri	h->2	
lfrå	g->9	
lfst	r->3	
lfte	 ->1	n->3	
lfun	k->2	n->1	
lfäl	l->97	
lfär	d->9	
lfån	g->4	
lföl	j->3	
lför	 ->3	.->1	a->2	b->4	e->7	f->2	l->4	s->14	v->2	
lgad	o->1	
lgar	i->1	
lgem	e->1	
lgen	 ->1	
lger	i->1	
lgie	n->9	
lgis	k->8	
lgiv	n->1	
lgjo	r->1	
lgod	o->1	
lgri	p->2	
lgru	n->2	
lgän	g->21	
lgån	g->25	
lgåv	o->1	
lgör	a->2	
lhan	d->43	
lhav	a->1	e->1	s->2	
lhel	m->1	
lhet	 ->11	,->7	.->1	?->1	e->1	s->3	
lhjä	r->8	
lhoe	k->1	
lhör	 ->4	a->3	i->1	
li -	 ->1	
li 1	9->4	
li 2	0->3	
li a	k->1	l->2	n->2	t->4	v->2	
li b	e->3	r->1	ä->1	
li d	e->3	o->2	
li e	f->2	n->18	t->11	
li f	l->2	r->1	ä->1	ö->9	
li g	a->1	
li h	a->1	e->1	
li j	u->1	
li k	l->3	o->1	
li l	e->1	i->2	ä->1	
li m	e->11	i->2	y->5	ö->3	
li n	ä->1	å->2	ö->2	
li o	b->1	m->1	t->1	
li p	l->1	r->2	
li r	i->1	
li s	l->1	t->3	u->1	v->1	y->1	ä->1	å->1	
li t	v->3	
li u	n->1	
li v	a->1	e->2	å->1	
li ä	m->1	
li ö	v->2	
li!J	a->1	
li, 	e->1	m->1	o->1	
li.U	t->1	
lia-	R->1	
lian	s->7	
liba	k->1	n->1	
libb	i->1	
libe	r->29	
libi	 ->1	
lic 	-->1	
lica	n->1	
lice	n->1	r->16	
lici	e->2	t->2	
lick	 ->4	,->1	.->2	a->2	b->5	e->10	o->1	
licy	,->1	a->1	d->1	f->1	
lida	 ->1	n->2	r->30	
lide	r->10	
lidi	t->3	
lien	 ->12	,->5	.->2	s->18	t->1	
lier	 ->4	a->1	n->1	
lies	t->1	
lifi	c->14	k->1	
lig 	a->11	b->9	d->14	e->7	f->30	g->8	h->9	i->14	j->2	k->19	l->7	m->13	n->8	o->23	p->9	r->15	s->28	t->14	u->20	v->2	y->1	å->2	ö->2	
lig!	H->1	
lig,	 ->13	
lig.	 ->2	D->2	G->2	J->4	O->3	V->2	
lig:	 ->2	
lig?	D->1	H->1	
liga	 ->633	,->18	.->18	/->1	;->1	?->1	d->1	n->5	r->67	s->10	t->16	
lige	n->481	
ligg	a->23	e->86	j->12	ö->21	
ligh	e->333	å->2	
ligi	e->1	ö->4	
ligs	e->1	
ligt	 ->641	!->2	,->30	.->55	:->1	;->1	v->101	
liho	p->1	
lik 	h->1	m->1	p->2	
lik.	D->1	
lik:	 ->1	
lika	 ->165	,->1	.->3	b->1	d->2	l->1	n->6	r->5	s->2	
like	n->11	r->4	
likg	i->2	
likh	e->35	
likn	a->21	i->44	
likr	i->3	
liks	o->47	t->2	
likt	 ->16	,->1	.->2	a->4	e->28	f->1	i->5	
likv	ä->8	
lill	a->4	f->1	i->1	
lima	n->3	t->14	
lime	n->1	
limi	n->6	
lims	o->1	
lin 	1->1	b->1	f->2	i->1	n->1	o->4	s->1	u->1	
lin,	 ->3	
lin.	L->1	O->1	
lina	r->1	
linb	a->1	
lind	a->3	r->4	u->56	
line	 ->1	r->3	
linf	r->1	
ling	 ->100	,->25	.->29	a->76	e->89	s->121	
lini	s->2	
linj	e->93	
link	o->2	
lino	r->1	
linr	i->5	å->1	
lins	b->1	
lint	 ->1	o->1	r->1	
linä	r->4	
liot	e->2	
lipp	e->2	
lir 	E->2	a->10	b->3	d->14	e->10	f->6	g->1	h->3	i->5	j->2	k->1	l->5	m->11	n->5	o->4	r->3	s->13	t->5	u->2	v->4	ä->1	å->1	ö->1	
lir,	 ->2	
lir:	 ->1	
lira	r->1	
lirt	a->1	
lis 	f->1	
lis,	 ->1	
lis.	V->1	
lis;	 ->1	
lisa	b->1	k->1	t->1	
lise	n->5	r->80	
lisi	o->3	ä->1	
lisk	 ->4	,->1	.->1	a->18	e->1	t->1	
lism	 ->7	.->3	?->1	e->3	y->2	
liss	a->1	e->1	t->1	
list	a->63	e->27	g->3	i->37	k->1	p->5	s->1	
lisv	ä->1	
lit 	-->1	a->2	b->1	e->3	f->2	h->1	i->1	m->1	o->2	p->2	s->4	t->1	ö->1	
lit,	 ->1	
lita	 ->5	d->1	n->1	r->13	t->7	
lite	 ->5	n->22	r->3	t->107	
liti	c->1	k->309	o->14	s->223	
litl	i->5	
lits	 ->4	.->2	
litt	e->8	r->4	
litä	r->6	
liv 	f->2	i->1	k->1	o->2	s->2	t->1	
liv,	 ->4	
liv.	A->1	D->1	I->1	M->1	V->1	
liva	 ->3	d->1	n->8	s->6	t->4	
live	t->25	
livi	e->1	t->26	
livs	c->3	d->2	k->6	m->88	u->1	v->1	
lixt	r->1	
lj L	i->1	
lj o	m->1	
lj ö	v->1	
lj, 	o->1	ä->1	
lj.V	i->1	
lja 	-->1	F->1	H->1	M->1	a->16	b->18	c->1	d->6	e->12	f->23	g->17	h->13	i->2	k->4	l->3	m->1	n->3	o->5	p->8	r->5	s->30	t->25	u->21	v->9	y->1	ö->1	
lja,	 ->5	
lja.	.->1	J->1	M->1	T->1	
ljad	e->3	
ljak	t->18	
ljan	 ->12	,->1	a->1	d->46	
ljar	 ->5	.->1	b->1	d->15	e->7	n->6	
ljas	 ->12	,->1	.->3	
ljat	 ->5	s->3	
ljd 	a->18	
ljd.	J->1	
ljde	 ->3	r->16	s->2	
ljdr	i->1	
ljds	k->2	
ljdå	t->1	
lje-	 ->1	
ljeb	e->1	o->4	ä->10	
ljed	o->1	
ljef	a->1	ö->2	
ljei	n->3	
ljej	o->3	
ljek	o->2	
ljel	i->1	s->3	
ljem	ä->1	
ljer	 ->38	,->4	.->1	a->16	n->4	
ljes	k->1	t->1	
ljet	a->9	r->2	
ljeu	t->2	
ljeå	t->1	
ljfl	ö->1	
ljko	n->2	
ljni	n->13	
ljon	 ->1	e->63	t->1	
ljs 	a->1	k->1	u->2	
ljs,	 ->1	
ljt 	i->1	u->1	v->1	
ljts	 ->2	
ljud	d->1	e->1	l->1	
ljug	e->1	
ljus	 ->1	.->1	e->8	
ljö 	f->2	i->1	k->1	m->1	s->2	v->1	
ljö!	D->1	
ljö,	 ->11	
ljö-	 ->2	
ljö.	D->3	M->1	U->1	V->1	
ljöa	n->3	v->1	
ljöb	e->3	r->1	
ljöd	e->1	i->1	
ljöe	r->4	
ljöf	a->2	r->4	ö->4	
ljöi	n->1	
ljök	a->11	o->6	r->8	v->1	
ljöl	a->1	
ljöm	i->1	ä->11	å->3	
ljön	 ->15	!->1	,->9	.->10	o->2	s->2	
ljöo	m->4	v->1	
ljöp	e->1	o->8	r->4	å->1	
ljör	å->1	ö->2	
ljös	e->1	i->1	k->15	t->1	y->6	
ljöu	t->1	
ljöv	ä->9	
lk a	t->1	
lk b	l->1	o->1	
lk h	a->1	
lk i	 ->2	
lk o	c->2	
lk r	e->1	
lk s	k->1	o->2	
lk t	v->1	
lk u	p->1	
lk, 	d->1	
lk.A	t->1	
lk.D	e->1	
lk.M	e->1	
lk.O	c->1	
lk.V	i->4	
lka 	a->1	b->2	d->8	e->3	f->9	g->5	i->2	j->1	k->16	l->4	m->6	n->2	o->4	p->4	r->1	s->11	t->3	u->4	v->5	ä->9	å->7	ö->1	
lkad	e->1	
lkan	 ->3	.->4	
lkar	 ->3	n->2	
lkas	 ->6	,->1	.->1	t->2	
lkat	s->1	
lkem	i->1	
lken	 ->56	,->1	s->4	
lkes	t->1	
lket	 ->185	,->1	.->1	:->1	i->2	s->4	
lkfr	o->1	
lkgr	u->2	
lkhä	l->9	
lkla	p->1	r->2	
lkli	g->1	n->1	
lkni	n->57	
lkoh	o->1	
lkom	l->5	m->11	n->42	r->6	s->3	
lkon	s->1	v->1	
lkor	 ->29	,->5	.->7	a->1	e->21	l->2	
lkpa	r->10	
lkre	g->1	p->3	t->4	
lkri	t->1	
lkrä	t->1	
lks 	f->1	s->2	
lkst	y->1	
lksw	a->1	
lksä	g->1	
lkur	s->1	
lkva	l->2	
lkvo	t->1	
lkyr	k->1	
lkän	d->2	n->9	t->1	
lköp	a->2	
ll "	M->1	
ll -	 ->3	
ll 1	0->1	5->1	9->3	
ll 2	 ->1	,->2	5->1	
ll 3	 ->1	0->1	
ll 4	 ->1	
ll 5	0->1	
ll 7	,->1	0->1	5->1	7->1	
ll 8	3->1	5->1	
ll 9	 ->1	1->1	4->2	
ll A	l->1	
ll B	a->1	o->2	r->2	
ll C	h->1	o->1	
ll D	i->1	
ll E	G->3	U->6	f->1	u->25	
ll F	r->3	ö->4	
ll G	e->1	r->1	
ll I	r->1	
ll K	a->2	i->3	o->9	u->1	
ll L	o->2	
ll M	c->1	i->1	o->2	
ll N	i->2	
ll O	L->1	
ll P	P->1	a->3	u->1	
ll R	a->1	
ll S	c->1	o->3	t->2	y->1	
ll T	h->1	i->1	r->1	y->2	
ll V	e->1	
ll W	a->2	i->1	u->1	
ll a	b->1	c->1	g->1	l->34	n->33	p->1	r->13	t->275	v->38	
ll b	a->17	e->79	i->7	l->25	o->6	r->5	u->1	y->2	ä->5	å->2	ö->12	
ll c	a->1	e->1	i->2	
ll d	a->1	e->281	i->28	o->4	r->3	u->1	ä->16	å->3	
ll e	f->3	g->3	k->2	l->3	m->3	n->111	r->15	t->31	u->3	x->46	
ll f	a->10	e->3	i->7	l->3	o->11	r->41	u->13	y->2	ä->2	å->11	ö->152	
ll g	a->7	e->32	i->1	l->1	o->10	r->19	ä->14	å->12	ö->23	
ll h	a->82	e->11	i->3	j->5	o->2	u->5	ä->5	å->2	ö->7	
ll i	 ->34	c->1	d->1	n->82	s->1	
ll j	a->108	o->1	u->6	ä->2	
ll k	a->11	l->4	n->1	o->82	r->6	u->57	v->1	ä->2	ö->1	
ll l	a->3	e->5	i->12	u->1	y->7	ä->12	å->3	ö->1	
ll m	a->20	e->30	i->25	o->5	u->1	y->7	ä->1	å->10	ö->5	
ll n	a->14	i->10	o->1	u->3	y->11	ä->13	å->11	ö->2	
ll o	a->1	c->71	e->1	f->2	i->1	j->1	l->6	m->23	p->1	r->8	s->4	ä->2	
ll p	a->10	e->8	i->1	l->2	o->5	r->19	u->2	å->13	
ll r	a->2	e->33	i->5	o->1	y->1	ä->20	å->20	ö->2	
ll s	a->13	e->17	i->35	j->6	k->38	l->17	m->2	n->1	o->34	p->4	t->73	u->6	v->2	y->6	ä->49	å->5	ö->1	
ll t	a->53	e->3	i->21	o->2	r->14	u->1	v->8	y->2	ä->2	
ll u	-->1	n->14	p->19	r->2	t->37	
ll v	a->55	e->18	i->67	o->3	ä->7	å->15	
ll y	r->2	t->3	
ll Ö	s->1	
ll ä	g->1	n->18	r->13	v->5	
ll å	k->1	r->2	s->2	t->19	
ll ö	k->6	n->1	p->3	s->1	v->15	
ll!H	e->1	
ll!J	a->1	
ll",	 ->2	
ll".	I->1	
ll, 	a->3	b->1	d->3	e->3	f->3	h->3	i->4	j->2	k->1	m->8	n->4	o->12	p->1	r->1	s->8	t->1	u->3	v->5	ä->3	å->2	
ll- 	o->4	
ll. 	D->1	o->1	
ll.A	n->1	v->1	
ll.B	i->1	
ll.D	e->21	ä->1	
ll.E	n->2	t->1	
ll.F	i->2	r->1	ö->2	
ll.H	a->1	e->3	ä->1	
ll.I	 ->4	n->1	
ll.J	a->11	
ll.K	o->3	
ll.M	e->2	å->1	
ll.O	m->1	r->1	
ll.P	r->1	å->1	
ll.R	e->1	
ll.S	a->1	m->1	o->1	å->2	
ll.T	a->1	ä->1	
ll.U	t->1	
ll.V	i->8	o->1	å->1	
ll.Ä	n->1	
ll: 	"->1	e->1	j->1	
ll?.	 ->1	
ll?D	a->1	
ll?H	u->1	
ll?J	a->1	
ll?K	o->1	
lla 	-->1	A->1	E->4	F->1	H->1	P->1	a->61	b->39	d->110	e->45	f->84	g->14	h->31	i->32	j->6	k->47	l->20	m->69	n->18	o->55	p->47	r->50	s->100	t->35	u->23	v->31	ä->5	å->10	ö->5	
lla!	H->1	
lla,	 ->13	
lla.	D->6	H->1	J->1	V->2	
lla:	F->1	
llad	 ->5	e->5	
llam	t->1	
llan	 ->194	"->1	,->3	.->2	d->145	l->1	n->1	s->7	t->2	ö->19	
llar	 ->16	,->3	.->1	;->1	e->5	n->4	
llas	 ->41	,->4	.->2	t->1	
llat	 ->5	
llav	a->1	
llba	k->52	r->26	
llbe	s->1	
llbi	l->1	
llbo	r->3	
llbr	i->4	
lld 	a->1	b->1	p->2	t->1	
llda	 ->11	,->4	.->6	s->2	
llde	 ->21	l->36	s->9	
lldh	e->23	
lldr	a->1	
lle 	-->1	E->3	K->1	a->25	b->20	d->41	e->8	f->31	g->17	h->23	i->26	j->44	k->66	l->5	m->5	n->4	o->12	p->5	r->5	s->30	t->14	u->16	v->123	ä->3	å->2	ö->2	
lle,	 ->3	
lle.	J->1	
lleg	a->71	e->127	i->4	o->4	
lleh	a->3	
llek	t->13	
llel	e->3	l->5	s->9	
llen	 ->65	"->1	,->10	.->19	a->6	n->7	s->2	Ä->1	
ller	 ->945	,->6	.->10	;->1	a->35	k->3	n->5	t->67	
lles	 ->6	a->5	
llet	 ->137	!->1	,->17	.->28	:->1	s->3	
lleu	r->2	
llfi	n->1	
llfo	g->6	
llfr	e->27	
llfu	n->1	
llfä	l->97	r->1	
llfö	l->3	r->17	
llgj	o->1	
llgo	d->1	
llgr	i->2	
llgä	n->21	
llgå	n->25	v->1	
llgö	r->1	
llha	n->43	
llhe	t->3	
llhö	r->8	
lli 	h->1	
lli!	J->1	
llia	n->7	
llib	e->1	
llie	r->1	
llig	 ->9	a->22	e->5	h->25	s->1	t->26	
llih	o->1	
llin	d->1	g->1	
llis	e->2	i->3	
llit	 ->21	,->1	e->1	s->6	
lliv	e->1	
llka	s->1	
llkl	a->2	
llko	m->11	r->64	
llkä	n->9	
llma	k->1	
llmo	s->1	
llmy	n->2	
llmä	n->125	r->1	t->2	
llmö	j->2	s->1	t->3	
llna	,->1	d->44	
llni	n->140	s->1	
llnä	r->6	
llo 	g->1	i->1	o->1	r->1	å->1	
llob	b->2	
lloj	a->2	
llok	e->1	
llol	j->1	
llom	r->1	
llor	 ->18	,->5	.->12	g->1	n->5	
llpo	l->1	
llra	 ->9	n->1	
llre	 ->6	
llri	n->1	s->1	
llrä	c->75	t->6	
lls 	C->1	a->7	b->3	d->4	e->1	f->1	h->13	i->17	k->1	m->2	n->1	o->2	p->5	s->7	t->4	u->3	v->7	ä->3	å->2	ö->1	
lls,	 ->4	
lls.	D->3	F->1	H->1	N->1	T->1	U->1	Y->1	
lls?	V->1	
llsa	m->32	t->3	
llsb	e->1	
llse	 ->13	k->3	
llsf	ö->1	
llsh	a->1	
llsi	d->1	
llsk	a->9	o->1	r->2	t->1	y->1	
llsl	i->1	u->1	ö->1	
llsm	e->1	ä->3	
llso	m->1	
llsr	i->2	
llss	e->1	t->3	
llst	i->7	o->3	r->4	u->1	ä->41	å->22	
llsv	a->3	i->1	ä->1	
llsy	n->2	s->3	
llsä	m->1	t->4	
llt 	-->1	1->1	a->23	b->12	d->42	e->6	f->38	g->8	h->2	i->28	k->19	l->1	m->17	n->7	o->19	p->13	r->4	s->56	t->7	u->20	v->15	y->1	ä->9	å->1	ö->3	
llt,	 ->17	
llt.	D->5	H->1	M->2	V->2	
llt:	 ->1	
llt;	 ->1	
llta	 ->1	g->1	l->1	
lltf	l->1	ö->39	
llti	d->77	h->1	n->5	
lltj	ä->3	
lltm	e->1	
lltr	o->1	ä->7	
llts	 ->9	:->1	a->1	e->3	å->63	
llut	i->1	s->14	
llva	l->1	r->74	
llve	r->87	
llvi	d->1	l->1	
llvä	g->8	n->1	r->2	x->20	
lly 	f->1	
lly!	 ->1	
lly.	A->1	
llyb	e->1	
llys	 ->1	
llyw	o->1	
lläg	g->18	n->2	
lläm	p->177	
llän	d->2	
llån	g->4	
llåt	 ->10	a->13	e->20	l->3	n->6	s->3	
llös	a->1	n->1	
lm d	e->1	
lm, 	h->1	
lm.H	e->1	
lmaj	o->1	
lmak	t->1	
lman	 ->7	!->242	,->157	:->1	n->11	s->9	
lmar	 ->2	
lmas	t->1	
lmed	e->2	v->1	
lmen	 ->1	t->2	
lmer	 ->1	
lmos	o->1	
lmsh	a->1	
lmyn	d->2	
lmän	 ->18	g->1	h->47	n->42	t->17	
lmär	k->2	
lmäs	s->2	
lmät	a->1	e->1	
lmåe	n->2	
lmöj	l->2	
lmös	s->1	
lmöt	e->3	
ln "	u->1	
ln a	t->1	
ln f	ö->3	
ln i	 ->2	
ln k	o->1	
ln m	e->1	
ln o	c->2	m->1	
ln t	i->5	
ln ä	r->2	
ln, 	d->1	h->1	
ln.D	e->1	
lna 	k->1	
lna,	 ->1	
lnad	 ->10	:->1	e->33	
lnin	g->212	
lnis	c->1	
lns 	l->2	
lnär	m->6	
lo g	o->1	å->1	
lo i	 ->1	
lo m	å->1	
lo o	c->3	
lo r	e->1	
lo å	t->1	
lo, 	W->1	s->2	
loak	l->1	
loba	l->12	
lobb	y->10	
lock	a->6	b->1	e->3	
lod 	t->2	
lode	n->2	
lodl	a->1	
log 	a->2	b->2	e->3	f->1	i->3	m->10	o->1	s->5	t->1	v->1	ä->1	å->1	
log,	 ->2	
log.	D->1	F->2	H->1	J->2	N->1	
loge	 ->1	,->1	n->8	
logi	 ->3	k->8	n->1	s->33	
logs	 ->4	
loja	l->7	
lok 	o->1	
loka	 ->1	l->44	s->1	
loke	r->1	
lokt	 ->5	
lola	d->1	
lolj	a->1	
loma	t->11	
lome	t->1	
lomm	a->1	o->2	
lomr	å->1	
loms	t->3	
lomä	s->1	
lona	p->2	
loni	a->1	
lonm	ä->1	
looi	j->1	
lopp	 ->7	,->1	.->1	e->12	
lor 	f->2	h->3	i->2	k->1	m->2	o->7	s->2	t->2	v->2	ä->2	
lor,	 ->6	
lor.	D->4	F->1	H->1	J->2	M->2	O->1	V->1	Ä->1	
lora	 ->4	d->5	r->4	t->8	
lore	n->19	
lorg	a->1	
lorn	a->5	
lors	 ->2	.->1	
los 	f->1	o->4	
losi	o->1	v->1	
loso	f->5	
loss	 ->1	a->1	n->1	
lot 	i->1	
lote	n->1	
lotp	r->2	
lott	 ->2	a->8	o->1	s->1	
lov 	a->1	i->1	
lova	 ->2	d->4	k->1	r->1	t->7	
love	n->1	
lovo	 ->1	r->2	
lovv	ä->2	
lovy	t->1	
loyd	s->1	
lp a	t->1	v->26	
lp d	e->1	
lp f	r->3	ö->3	
lp n	i->1	
lp o	c->2	
lp p	å->1	
lp s	k->1	o->1	
lp t	i->5	
lp v	i->2	
lp ö	v->1	
lp, 	d->1	m->1	
lp.D	e->1	
lp.H	ä->1	
lp.I	 ->1	
lp.J	a->1	
lp.V	i->1	
lpa 	W->1	a->1	d->5	f->2	g->1	h->1	i->1	k->2	l->1	m->8	o->3	p->1	s->2	t->7	v->1	
lpan	d->3	
lpar	e->1	k->6	l->1	
lpat	r->1	
lpe 	p->1	
lpen	 ->4	
lper	 ->1	n->1	
lpes	 ->1	
lpla	n->1	
lpli	g->1	
lpol	i->45	
lpro	b->1	d->2	g->1	
lps.	J->1	
lpt 	t->1	
lpta	.->1	
lpte	 ->1	
lpun	k->2	
lpvi	l->1	
lra 	b->2	f->1	h->1	s->3	v->2	
lran	d->1	
lrap	p->1	
lre 	H->1	a->1	b->1	h->1	s->1	v->1	
lreg	e->1	l->4	
lres	u->4	
lrik	a->4	t->1	
lrin	g->1	
lris	k->1	
lrol	l->1	
lrum	 ->1	
lryc	k->1	
lräc	k->75	
lräk	e->1	n->1	
lrät	t->11	
ls C	E->1	
ls a	l->3	n->2	r->3	t->4	v->5	
ls b	a->1	e->2	l->1	
ls d	e->3	r->1	ä->1	
ls e	n->1	x->1	
ls f	a->2	i->1	r->1	u->1	ö->3	
ls g	a->1	
ls h	a->11	e->1	u->1	ä->1	
ls i	 ->7	l->1	n->12	
ls k	o->1	u->1	v->1	
ls l	i->2	
ls m	e->3	i->3	ä->2	å->1	
ls n	å->1	
ls o	c->4	l->1	r->2	
ls p	r->4	å->5	
ls s	a->2	e->1	k->4	o->3	t->1	
ls t	i->6	r->1	v->1	
ls u	p->1	t->3	
ls v	a->4	i->3	ä->2	
ls ä	n->1	r->2	
ls å	r->2	s->1	t->3	
ls ö	v->1	
ls, 	f->1	g->1	o->1	p->1	
ls- 	o->1	
ls.D	e->4	
ls.F	ö->1	
ls.H	a->1	
ls.N	u->1	
ls.T	a->1	
ls.U	n->1	
ls.Y	t->1	
ls?V	i->1	
lsa 	k->1	o->11	p->1	s->1	t->1	
lsa,	 ->3	
lsa.	H->1	
lsac	e->3	
lsam	h->1	m->31	
lsan	 ->1	,->2	.->1	
lsar	 ->1	
lsat	s->1	t->3	
lsav	g->1	
lsbe	d->1	
lsbu	r->1	
lsdo	m->1	
lsdr	ä->1	
lse 	-->3	a->27	b->1	d->2	e->1	f->16	g->3	h->3	i->5	j->3	k->5	m->15	n->4	o->17	p->2	r->1	s->20	t->2	u->1	v->1	ä->3	ö->4	
lse,	 ->12	
lse-	 ->1	
lse.	B->1	D->5	E->2	J->3	K->1	L->1	M->2	N->1	S->2	V->2	
lsea	k->1	
lseb	y->1	
lsef	u->11	
lseh	i->1	
lsek	o->5	r->2	t->6	
lsel	e->2	ö->3	
lsem	ö->1	
lsen	 ->41	,->3	.->5	l->2	s->4	
lseo	m->1	
lser	 ->88	!->1	,->19	.->13	:->1	i->1	n->52	s->1	
lseu	t->1	
lsev	i->2	
lsex	p->1	
lsfa	l->1	s->1	
lsfl	o->2	
lsfr	å->2	
lsfö	r->2	
lsha	n->2	
lshi	n->1	
lsid	i->1	
lsig	n->1	
lsik	e->1	
lsin	d->2	g->20	
lsit	u->1	
lsk-	f->1	
lska	 ->14	.->1	:->1	n->2	p->9	r->1	t->3	
lske	n->1	
lski	f->1	
lskn	i->1	
lsko	m->1	n->2	t->1	
lskr	i->4	o->4	
lskt	 ->2	.->1	
lsku	l->1	
lskv	a->1	
lsky	d->4	n->1	
lskö	p->1	
lsla	g->5	
lsli	g->1	
lslo	g->1	
lslu	t->1	
lslö	s->2	
lsme	d->1	
lsmy	n->9	
lsmä	n->2	s->4	
lsni	n->2	
lsny	h->1	
lso-	 ->1	
lsoc	i->1	
lsoe	f->1	
lsom	g->1	r->2	
lson	 ->4	.->1	
lsor	e->1	g->3	i->1	
lsos	k->1	
lsov	å->3	
lspa	r->1	
lspl	a->2	
lspo	l->2	
lspr	i->1	o->3	
lspu	n->6	
lsri	k->2	
lsru	h->2	n->1	
lsse	k->1	r->1	
lssi	d->1	
lssj	ö->1	
lsst	i->1	r->3	ö->1	
lssy	s->1	
lssä	k->43	
lst 	a->2	b->1	f->1	h->1	i->6	k->1	l->1	m->3	n->1	p->2	r->1	s->7	t->2	u->1	v->4	ä->1	
lst,	 ->7	
lst.	 ->1	A->1	D->1	F->1	V->1	
lsta	t->7	
lste	r->1	
lsth	o->3	
lsti	l->9	
lsto	l->4	r->41	
lstr	u->1	ö->4	
lstu	d->1	
lstv	i->1	
lstä	n->41	
lstå	n->28	
lstö	d->2	
lsum	m->1	
lsut	a->3	s->1	
lsva	r->4	
lsvi	l->1	
lsvä	r->1	s->1	
lsyn	.->1	t->2	
lsys	t->6	
lsäm	n->1	
lsät	t->123	
lsök	a->6	
lt -	 ->2	
lt 1	8->1	
lt 2	7->1	
lt 7	0->1	
lt 9	5->1	
lt E	U->4	
lt S	t->1	u->1	
lt a	b->1	d->1	k->1	l->1	n->14	r->1	t->22	v->6	
lt b	e->12	i->1	l->2	o->1	r->1	u->2	ä->1	ö->3	
lt d	e->48	i->1	o->1	r->2	ä->2	
lt e	f->3	k->1	l->1	n->25	r->2	t->5	
lt f	a->4	e->1	i->6	l->3	o->1	r->7	ä->1	å->1	ö->42	
lt g	e->5	i->1	l->1	o->5	y->1	ä->3	
lt h	a->9	e->1	ä->2	
lt i	 ->33	l->1	m->1	n->24	
lt j	o->1	u->1	
lt k	a->4	l->16	o->20	r->1	u->2	ä->4	
lt l	i->1	o->1	y->1	ä->1	
lt m	e->22	i->4	o->2	y->1	ä->1	å->3	
lt n	a->1	o->3	y->3	ä->8	å->2	ö->3	
lt o	a->3	c->31	f->2	l->1	m->8	r->4	s->3	t->1	v->1	
lt p	a->2	l->4	o->2	r->3	u->2	å->16	
lt r	a->1	e->2	i->7	ä->8	
lt s	a->12	e->13	i->4	j->2	k->8	n->1	o->10	p->1	t->16	v->2	y->1	ä->15	å->1	ö->1	
lt t	a->2	i->16	r->3	v->1	y->4	
lt u	n->4	p->9	r->1	t->17	
lt v	a->8	i->20	ä->5	å->4	
lt y	t->1	
lt ä	n->4	r->9	v->1	
lt å	t->3	v->1	
lt ö	p->1	v->11	
lt, 	a->1	b->2	d->1	e->1	f->2	j->1	m->3	o->6	s->1	t->1	u->1	v->2	ä->1	å->1	
lt. 	D->1	
lt.D	e->10	
lt.E	n->1	
lt.H	e->2	ä->1	
lt.I	 ->1	
lt.J	a->2	
lt.M	a->1	e->1	
lt.O	m->1	
lt.U	n->1	
lt.V	a->3	i->3	
lt: 	a->1	
lt; 	d->2	
lt?J	a->1	
lta 	f->1	i->13	o->3	p->2	s->1	u->1	ä->2	ö->2	
lta,	 ->3	
ltag	a->25	i->6	
ltak	t->1	
ltal	a->1	i->2	
ltar	 ->10	e->1	
ltas	 ->1	
ltat	 ->31	,->6	.->10	:->1	?->2	e->44	i->3	l->1	t->7	ö->6	
ltba	s->1	
lte 	k->1	v->1	
lte,	 ->2	
lten	 ->7	!->2	,->1	.->4	a->1	b->4	e->18	s->3	
lter	 ->2	a->8	n->12	
ltes	i->3	
ltet	 ->5	"->1	.->3	
ltfl	e->1	
ltfö	r->39	
lthe	n->6	t->2	
ltib	e->1	
ltid	 ->74	,->2	.->1	a->1	e->1	s->1	
ltie	t->3	
ltig	 ->3	a->7	h->12	t->4	
ltih	o->1	
ltil	a->1	l->17	
ltim	a->1	
ltin	a->5	g->5	
ltis	k->1	
ltjä	m->3	
ltme	r->1	
ltni	n->48	
ltog	 ->2	
lton	.->1	
ltra	f->1	l->1	p->1	
ltre	r->1	
ltro	 ->1	
lträ	d->7	
lts 	-->1	a->1	f->1	i->2	m->1	o->2	p->1	s->1	t->1	u->1	ä->1	
lts.	K->1	
lts:	 ->1	
ltsa	m->1	
ltse	d->3	
ltsi	t->1	
ltså	 ->61	,->2	
ltur	 ->41	,->11	-->1	.->3	?->1	a->8	e->64	f->1	h->1	o->1	p->8	s->5	u->1	
ltäc	k->4	
luck	a->3	o->2	
ludd	i->2	
lude	r->4	
luft	b->1	o->1	
lufö	r->1	
lugn	 ->1	a->5	
luka	r->2	s->1	
lukt	 ->1	a->1	
lump	 ->3	.->1	
lumr	a->1	
lunc	h->1	
lund	a->14	r->1	
lunt	a->4	o->1	
lups	k->1	
lura	l->1	s->1	t->1	
lure	s->1	
lus 	a->1	t->1	
lusi	v->20	
luss	a->2	
lust	 ->1	.->1	b->1	e->7	
lut 	-->1	8->2	9->1	a->7	b->6	d->1	e->2	f->10	g->1	h->4	i->16	k->3	l->4	m->3	n->11	o->26	p->11	r->1	s->16	t->2	u->4	v->3	ä->4	å->1	
lut,	 ->14	
lut.	 ->1	D->3	F->1	I->1	N->2	O->1	S->1	T->1	V->1	
lut;	 ->1	
luta	 ->44	,->5	d->30	f->10	n->32	p->1	r->9	s->10	t->14	u->3	
lutb	e->2	i->3	
lute	n->15	r->8	t->55	
lutf	ö->9	
lutg	i->8	
luth	a->1	e->1	
luti	o->101	t->4	
lutk	o->1	
lutl	i->72	
lutn	a->15	i->40	
lutp	e->1	
lutr	e->3	
luts	 ->1	a->55	c->1	f->12	k->14	p->4	r->1	t->1	
lutv	e->3	
lutä	n->5	
lux,	 ->1	
lv a	n->1	r->1	t->3	
lv b	e->1	i->1	
lv d	a->1	
lv f	r->2	ö->3	
lv g	o->1	
lv h	a->2	ö->1	
lv i	 ->3	
lv k	o->1	
lv m	e->2	
lv o	c->3	
lv s	a->1	e->1	k->1	o->3	ä->1	
lv t	a->1	i->2	
lv u	n->1	t->1	
lv v	a->1	e->1	
lv ä	r->3	
lv å	r->1	
lv, 	h->3	m->2	
lv.D	e->1	
lv.J	a->1	
lv.K	o->1	
lv.V	i->1	
lva 	E->1	a->2	b->5	d->3	f->1	h->1	i->1	k->6	l->1	m->1	o->4	r->1	s->5	t->3	u->1	v->28	ä->2	å->2	
lva,	 ->3	
lva.	D->1	L->1	N->1	O->1	V->1	
lval	.->1	
lvan	d->1	
lvar	 ->6	,->1	.->4	e->1	l->62	
lvbe	s->3	
lvbi	o->1	
lvbä	r->1	
lver	 ->2	,->1	a->9	k->113	s->1	
lvet	 ->1	
lvfa	l->2	
lvfö	r->1	
lvhj	ä->2	
lvid	a->1	
lvil	l->1	
lvin	i->1	
lvis	 ->38	,->2	
lvkl	a->20	
lvko	s->1	
lvmi	l->1	
lvni	n->3	
lvof	f->1	
lvol	y->1	
lvpl	å->1	
lvra	k->6	
lvst	y->7	ä->8	
lvsä	k->1	
lvt 	d->1	h->2	k->1	s->1	å->2	
lvti	d->1	m->2	
lvvä	g->2	
lväg	a->8	g->3	
lvän	d->1	n->1	t->1	
lvär	d->2	
lväx	t->20	
lvår	 ->1	e->2	s->2	
lvö,	 ->1	
lvö.	D->1	
lvön	 ->1	
ly f	ö->1	
ly å	t->1	
ly! 	G->1	
ly, 	k->2	
ly.A	n->1	
ly.V	i->1	
lybe	t->1	
lyck	a->85	l->9	o->17	s->9	ö->5	
lyda	 ->2	n->1	
lyde	l->2	r->3	
lyft	 ->2	a->6	e->2	o->3	
lyg,	 ->1	
lyga	 ->1	n->1	
lygb	l->1	
lyge	r->1	t->1	
lygk	r->1	
lygn	i->1	
lygp	l->4	
lygs	a->4	
lygt	r->2	
lykt	a->1	e->3	i->13	
lym 	a->1	o->1	
lyme	n->1	r->1	
lymp	i->2	
lyr 	f->1	
lys 	-->1	a->16	b->1	f->2	g->1	i->1	j->1	o->2	s->1	v->1	
lys,	 ->4	
lys.	D->2	F->1	G->1	H->1	
lys?	D->1	I->1	
lysa	 ->5	n->4	t->2	
lyse	n->5	r->18	
lysn	i->4	
lyss	n->29	
lyst	 ->2	
lyta	n->12	
lyte	l->1	
lytt	 ->1	.->1	a->11	n->4	
lyve	r->1	
lywo	o->1	
lz e	n->1	
lz s	a->2	
lzen	.->1	
lzma	n->2	
läck	a->3	e->1	o->1	t->3	
läde	r->22	
lädj	a->8	e->7	
läds	 ->6	
läga	r->1	
läge	 ->9	,->1	.->2	n->15	r->1	s->3	t->19	
lägg	 ->20	,->1	.->1	a->180	e->43	n->27	s->21	
lägl	i->1	
lägn	a->8	
lägr	e->11	
lägs	e->6	n->5	t->1	
läka	r->5	
läke	m->1	
läkt	a->3	e->1	i->1	
lämn	a->81	i->5	
lämp	a->100	l->60	n->68	
länd	a->4	e->185	s->26	
läng	a->1	d->4	e->35	n->3	r->62	s->2	t->1	
länk	a->2	
länn	i->1	
länt	.->1	
läpa	d->1	
läpp	 ->2	,->1	.->1	a->6	e->5	h->1	s->1	t->3	
lär 	e->1	
lära	 ->7	r->2	
lärd	e->1	o->7	
lärl	i->1	
läro	a->1	s->1	
lärt	 ->3	
läs 	t->1	u->1	y->1	
läsa	 ->3	
läsb	a->2	
läse	r->6	
läsf	r->1	
läsk	u->1	
läsn	i->2	
läst	 ->4	a->1	e->1	
lät 	d->1	m->1	s->3	
lätt	 ->9	.->2	a->39	f->1	i->2	n->1	v->2	
läxa	n->1	t->1	
läxo	r->1	
lå E	u->1	
lå a	t->6	
lå b	a->1	
lå e	l->1	n->3	
lå f	a->6	
lå i	h->1	
lå k	o->4	
lå m	e->2	
lå n	å->1	
lå p	r->1	
lå r	å->1	
lå s	a->1	i->1	
lå v	a->2	e->1	i->1	
låda	 ->1	
låde	f->1	r->11	
låen	d->1	
låg 	a->1	d->1	h->1	i->1	n->2	t->1	
låga	 ->5	
låge	r->1	
lågt	 ->2	
låna	n->1	
lånb	o->1	
lång	 ->34	,->1	.->1	a->10	d->1	f->2	r->1	s->13	t->52	v->6	
låni	n->1	
lår 	B->1	a->7	d->3	e->6	f->1	i->4	j->4	k->2	m->2	n->1	r->1	s->2	t->1	v->6	ä->2	
lår"	.->1	
lår.	 ->1	M->1	
lår?	S->1	
lås 	a->3	b->2	d->2	e->1	g->2	i->11	m->1	p->1	t->2	
lås.	D->1	
låse	r->3	
låss	 ->1	
låst	 ->1	a->2	
låt 	e->1	m->15	o->8	
låta	 ->41	n->3	s->6	
låte	n->6	r->23	t->1	
låti	t->3	
låtl	i->5	
låtn	a->6	
låts	 ->4	a->2	
léch	a->1	
löde	n->1	t->2	
lödi	g->1	
löft	e->11	
löja	d->1	n->1	r->3	s->1	
löje	v->3	
lökm	o->1	
lömm	a->14	e->2	
löms	k->1	
lömt	 ->4	
lön 	f->1	
löna	r->1	s->1	
löne	-->1	a->1	r->1	
löns	a->5	
lönt	 ->1	a->3	
löpa	 ->2	n->6	
löpe	r->10	
löpt	 ->5	e->2	
lörd	a->1	
lös 	-->1	d->1	e->1	k->1	s->1	
lös.	D->1	
lösa	 ->38	,->3	.->3	r->1	s->6	
löse	r->4	s->1	
lösg	ö->1	
lösh	e->44	
lösn	i->52	
lösr	y->1	
löst	 ->10	,->1	a->6	e->1	s->1	
löt 	a->1	d->1	v->1	
löts	l->4	
lövs	k->1	
løn,	 ->2	
m "E	q->1	u->1	
m "K	u->1	v->1	
m "n	å->1	
m "o	r->1	
m "v	a->1	
m "ö	p->1	
m - 	K->1	a->4	e->1	i->1	k->1	m->2	o->3	p->1	s->2	t->1	v->2	
m 1 	0->1	
m 15	0->1	
m 16	 ->1	
m 19	8->1	9->2	
m 20	 ->3	
m 28	 ->1	
m 3-	l->2	
m 31	4->1	
m 35	 ->2	0->1	
m 40	 ->2	0->1	
m 45	 ->1	
m 50	 ->1	
m 5b	-->1	
m 6,	0->1	
m 80	 ->1	
m Ag	u->1	
m Ah	e->1	
m Al	a->1	p->1	
m Am	o->1	s->2	
m Ap	a->1	
m At	l->1	
m BS	E->1	
m Ba	r->1	
m Be	l->1	r->5	
m Bl	a->1	
m Bo	w->1	
m Br	i->1	y->1	
m CE	N->1	
m Ce	y->1	
m Co	c->1	x->1	
m Da	 ->1	l->1	n->2	
m De	 ->1	t->1	
m Di	m->1	
m Du	t->1	
m EG	-->3	
m EM	U->1	
m EU	 ->11	,->1	-->2	.->3	:->3	
m Eh	u->1	
m El	l->1	
m Er	i->1	
m Et	i->1	
m Eu	r->73	
m FB	I->1	
m FP	Ö->1	
m Fl	o->1	
m Fr	a->2	
m Fö	r->4	
m GU	S->1	
m Ga	l->1	
m Ge	n->2	
m Go	l->1	o->1	
m Gr	e->2	
m Ha	i->3	t->2	
m He	d->1	
m Hi	t->1	
m IN	T->1	
m In	d->1	
m Ir	l->1	
m Is	r->1	
m It	a->2	
m Jo	n->2	
m Jö	r->2	
m Ka	u->1	
m Ko	s->4	u->1	
m La	n->6	
m Li	b->1	
m Ll	o->1	
m Ma	l->1	r->1	
m Mc	C->1	N->1	
m Ne	d->1	
m Of	f->1	
m PP	E->1	
m Pa	k->1	l->1	y->1	
m Po	r->1	w->3	
m Pr	o->1	
m Ra	c->1	
m Ri	c->1	
m Ro	t->1	
m SE	K->1	
m Sc	h->3	
m Se	i->2	
m Sj	ä->1	
m Sk	o->1	
m Sp	e->1	
m Sy	r->1	
m Ta	m->1	
m Th	e->3	
m Ti	b->2	
m To	r->1	t->1	
m Tu	r->4	
m Vä	r->1	
m Wa	l->2	
m Wi	e->1	
m a 	p->1	
m ab	s->2	
m ac	c->1	
m ad	v->2	
m ag	e->3	r->1	
m al	d->1	l->57	t->1	
m am	b->1	e->1	
m an	d->10	f->2	g->3	k->1	l->2	n->2	o->1	s->25	t->13	v->8	
m ap	p->1	
m ar	b->17	g->1	m->1	r->1	t->2	
m as	y->5	
m at	t->398	
m av	 ->53	,->1	f->2	g->7	k->2	l->2	s->10	t->1	v->2	
m b)	 ->1	
m ba	k->2	l->1	n->1	r->3	
m be	a->2	d->8	f->9	g->7	h->30	k->10	l->1	m->1	o->1	r->15	s->28	t->20	v->6	
m bi	d->7	l->2	n->1	o->1	t->1	
m bl	.->2	a->2	e->2	i->4	y->1	
m bo	r->12	s->2	t->1	
m br	i->3	o->4	u->1	y->2	å->3	
m bu	d->4	
m by	g->1	r->1	
m bä	r->5	t->2	
m bå	d->5	
m bö	c->1	r->14	t->1	
m c)	 ->1	
m ca	n->1	
m ce	n->1	
m ch	a->1	o->1	
m co	r->2	
m da	g->8	m->1	
m de	 ->161	,->1	b->3	c->1	f->3	l->7	m->6	n->149	r->3	s->36	t->296	
m di	a->1	f->1	k->1	o->1	p->1	r->7	s->8	
m dj	ä->1	
m do	g->1	m->5	
m dr	a->12	i->3	y->1	
m du	 ->1	b->1	
m dy	k->1	
m dä	r->12	
m då	 ->6	l->2	
m dö	d->1	e->1	l->1	m->1	
m ef	f->3	t->10	
m eg	e->5	n->1	
m ej	 ->1	
m ek	o->5	
m el	-->4	e->1	l->5	
m em	e->1	o->17	
m en	 ->184	b->1	d->6	e->5	h->1	l->4	o->1	s->3	
m er	 ->3	a->4	f->1	k->1	s->1	t->5	ö->1	
m et	c->1	t->125	
m eu	r->10	
m ex	 ->1	a->2	c->2	e->9	p->1	
m fa	d->1	k->3	l->7	r->1	s->11	t->9	
m fe	m->2	
m fi	c->1	n->39	s->4	
m fj	o->1	
m fl	a->1	e->6	y->5	
m fo	d->1	l->2	n->1	r->18	s->1	
m fr	a->29	e->6	i->8	u->2	ä->1	å->19	
m fu	l->1	n->4	s->1	
m fy	l->1	r->1	
m fä	l->1	r->1	
m få	r->6	t->3	
m fö	l->8	r->287	
m ga	m->1	r->5	v->1	
m ge	 ->2	m->19	n->14	r->10	s->4	t->1	
m gi	c->1	l->2	v->1	
m gj	o->10	
m gl	o->1	
m go	d->8	
m gr	a->2	i->2	u->13	ä->2	
m gä	l->22	
m gå	n->1	r->9	t->2	
m gö	m->1	r->36	
m ha	 ->1	d->4	m->3	n->42	r->152	s->1	v->2	
m he	d->1	l->52	r->3	t->1	
m hi	n->2	t->12	
m hj	ä->6	
m ho	b->1	n->10	t->3	
m hu	m->2	r->32	
m hy	s->1	
m hä	l->2	n->18	r->18	v->4	
m hå	l->8	r->1	
m hö	g->4	r->3	
m i 	B->2	C->1	E->2	G->1	H->1	N->1	T->4	U->1	a->2	b->3	d->34	e->4	f->18	g->1	h->7	k->1	l->1	m->15	n->2	o->3	p->7	r->4	s->20	t->3	u->1	v->7	Ö->1	å->1	ö->1	
m ic	k->4	
m id	é->1	
m if	a->1	r->1	
m ig	e->1	
m ih	å->1	
m in	 ->1	b->1	d->6	f->18	g->11	i->2	k->1	l->9	n->29	o->8	r->7	s->4	t->108	v->3	
m is	r->1	
m ja	g->136	
m jo	r->6	
m ju	 ->5	s->9	
m jä	m->2	r->1	
m ka	m->1	n->58	p->4	r->5	
m ke	m->1	
m kl	a->2	
m ko	a->1	d->1	l->4	m->146	n->32	r->10	s->6	
m kr	a->3	i->6	ä->18	
m ku	l->7	n->1	r->1	
m kv	a->1	i->1	
m kä	n->6	r->6	
m kö	p->1	r->1	
m la	d->4	g->15	n->2	
m le	d->30	g->1	t->1	v->6	
m li	b->2	g->16	k->5	t->2	v->16	
m lj	u->1	
m lo	k->1	
m ly	c->2	d->1	f->1	k->1	s->1	
m lä	c->1	g->8	k->1	m->11	n->5	t->1	
m lå	g->2	n->2	
m lö	p->1	s->4	
m ma	i->1	j->2	k->1	n->98	r->5	x->1	
m me	d->68	l->3	n->5	r->7	s->1	
m mi	l->9	n->19	s->4	t->1	
m mo	d->3	t->13	
m mu	s->1	
m my	c->9	n->8	
m mä	n->13	r->1	
m må	h->1	l->2	n->5	s->32	
m mö	j->52	
m na	r->1	t->9	z->3	
m ne	d->2	g->1	k->1	
m ni	 ->64	,->5	.->1	o->1	
m no	r->2	
m nu	 ->25	m->1	
m ny	 ->1	a->2	l->2	s->1	t->1	
m nä	m->5	r->11	s->1	
m nå	g->30	
m nö	d->1	t->1	
m oa	c->1	
m ob	e->2	
m oc	h->72	k->20	
m of	f->3	t->4	
m og	e->1	
m ol	i->3	j->2	y->1	
m om	 ->41	b->1	e->1	f->5	l->1	r->10	s->1	ö->1	
m on	ö->1	
m or	d->11	i->1	o->2	s->3	
m os	s->4	
m ot	i->1	
m pa	r->25	
m pe	k->2	n->2	r->3	
m pl	a->4	
m po	l->6	s->1	ä->1	
m pr	a->2	e->3	i->7	o->11	
m pu	b->1	m->1	n->2	
m på	 ->52	.->1	g->1	m->1	p->1	t->2	v->8	
m ra	d->1	m->52	p->1	s->2	t->1	
m re	d->35	f->9	g->25	k->1	l->8	p->1	s->16	t->1	v->2	
m ri	k->5	m->2	s->8	
m ro	l->1	
m ru	l->2	s->1	
m ry	g->1	s->1	
m rä	c->1	k->1	t->14	
m rå	d->36	
m rö	r->13	s->3	v->1	
m s.	k->1	
m sa	d->3	g->4	k->7	m->35	n->1	t->2	
m sc	h->1	
m se	d->5	g->3	k->2	n->1	r->5	x->1	
m si	n->6	t->8	
m sj	u->2	ä->1	ö->1	
m sk	a->79	e->12	i->3	j->1	o->5	r->7	u->27	y->5	ö->1	
m sl	o->1	u->7	
m sm	å->3	
m sn	a->2	e->1	
m so	c->2	l->1	m->132	
m sp	e->9	o->1	r->3	
m st	a->15	e->1	i->1	o->2	r->11	y->3	ä->14	å->27	ö->15	
m su	b->4	
m sv	a->3	
m sy	f->9	n->2	s->10	
m sä	g->2	k->17	r->3	t->1	
m så	 ->19	d->8	l->1	t->1	
m sö	k->1	r->2	
m t.	e->2	o->1	
m ta	g->2	l->6	n->2	r->6	s->5	x->1	
m ti	b->1	d->12	l->112	o->1	
m tj	ä->3	
m to	g->5	l->5	
m tr	a->17	e->6	o->2	ä->5	
m tu	r->1	
m tv	e->1	å->5	
m ty	c->2	d->5	n->1	s->1	v->2	
m tä	c->2	n->1	p->1	
m un	d->20	i->22	
m up	p->36	
m ur	 ->2	s->7	
m ut	 ->1	.->1	a->7	b->5	d->1	e->1	f->7	g->11	i->1	j->1	l->2	m->2	n->1	r->2	s->12	t->14	v->13	ö->1	
m va	d->16	g->1	l->4	n->4	r->40	
m ve	d->1	l->1	m->2	r->20	t->5	
m vi	 ->280	,->3	?->1	a->1	d->13	k->2	l->39	n->1	s->24	t->5	
m vo	n->3	r->2	
m vr	ä->1	
m vu	x->1	
m vä	c->3	g->4	l->4	n->2	r->1	s->1	
m vå	r->19	
m yr	k->1	
m yt	t->4	
m Ös	t->4	
m äg	e->2	n->1	t->1	
m än	 ->6	d->17	n->4	t->3	
m är	 ->191	,->1	
m ät	e->1	
m äv	e->15	
m åk	l->1	t->1	
m ål	a->1	i->1	
m år	 ->8	,->1	.->2	e->5	s->2	
m ås	a->1	i->1	t->1	y->4	
m åt	e->17	g->7	m->1	
m öa	r->1	
m ök	a->3	n->1	
m öm	s->1	
m ön	s->1	
m öp	p->7	
m ör	o->1	
m ös	t->2	
m öv	e->23	r->1	
m!De	n->1	t->1	
m!Me	n->1	
m!Tr	o->1	
m".D	e->1	
m) o	m->1	
m); 	a->1	
m, K	u->1	
m, a	l->2	n->2	t->4	v->1	
m, b	l->1	å->1	ö->2	
m, d	e->11	ä->1	å->1	
m, e	f->5	n->3	t->1	x->1	
m, f	i->1	r->3	ö->3	
m, g	e->1	r->1	
m, h	a->3	e->2	u->1	
m, i	 ->5	d->1	n->1	
m, j	a->1	u->2	
m, k	a->2	r->1	v->1	
m, l	e->1	
m, m	e->12	
m, n	a->1	i->1	ä->2	å->1	
m, o	c->20	m->1	p->1	r->1	
m, p	r->1	å->4	
m, r	e->1	
m, s	a->1	e->1	o->7	p->1	ä->2	å->5	
m, t	i->1	r->1	
m, u	p->1	t->8	
m, v	a->3	e->1	i->9	
m, ä	n->1	r->3	v->5	
m, å	t->1	
m- o	c->1	
m-el	-->1	
m. D	e->1	ä->1	å->1	
m. H	o->1	u->1	
m. M	a->1	
m. a	v->2	
m. d	e->1	
m. i	 ->1	
m. ä	n->1	r->1	
m.(A	p->1	
m., 	d->1	
m.. 	F->1	
m..(	F->1	
m.Al	l->1	
m.At	t->1	
m.Av	 ->1	b->1	s->1	
m.Be	t->1	
m.Bu	d->1	
m.De	 ->5	n->7	s->2	t->24	
m.Dä	r->5	
m.EG	-->1	
m.EK	S->1	
m.En	 ->1	
m.Eu	r->1	
m.Ex	p->1	
m.Fr	u->5	
m.Fö	r->3	
m.Ge	n->2	
m.Gö	r->1	
m.He	r->10	
m.Hu	r->2	
m.I 	d->2	n->1	r->1	
m.In	f->1	o->1	
m.Ja	g->17	
m.Ko	m->1	s->1	
m.Ku	l->1	
m.Lå	t->1	
m.Ma	n->1	
m.Me	d->3	n->9	
m.Må	n->1	
m.Na	t->1	
m.Ne	j->1	
m.Ni	 ->1	
m.Nu	 ->1	
m.Nä	r->3	
m.Nå	g->1	
m.OM	R->1	
m.Oc	h->4	
m.Om	 ->2	
m.Pr	o->2	
m.Re	f->1	s->1	
m.Rå	d->1	
m.Sa	m->1	
m.Sl	u->2	
m.So	m->2	
m.St	a->2	
m.Sy	f->1	
m.Så	 ->1	
m.Ti	l->1	
m.Tr	o->1	
m.Ty	v->1	
m.Ur	 ->1	
m.Va	d->1	
m.Ve	m->1	
m.Vi	 ->16	d->2	l->1	
m.m.	O->1	
m.Än	d->1	
m.Är	 ->1	
m/ri	k->1	
m: A	s->1	
m: N	ä->1	
m: d	e->2	u->1	
m: e	n->1	
m: p	a->1	
m; d	e->2	
m?De	t->1	
m?Ja	g->1	
m?Me	n->1	
m?Vi	l->2	
mI. 	f->1	
ma -	 ->2	
ma 1	6->1	
ma B	r->1	
ma E	u->1	
ma H	a->2	
ma M	a->1	
ma a	l->2	m->1	n->2	r->3	t->15	v->2	
ma b	e->5	i->2	o->4	r->1	ä->1	
ma d	a->1	e->22	i->1	r->1	
ma e	n->6	r->1	t->3	u->2	
ma f	a->1	i->1	r->11	ö->17	
ma g	r->1	ä->2	å->1	
ma h	a->3	i->2	o->1	u->1	ä->3	å->1	ö->1	
ma i	 ->12	.->2	f->2	g->1	h->14	n->15	v->1	
ma j	o->5	
ma k	a->2	l->1	o->7	r->5	u->2	ä->1	
ma l	a->2	i->1	ä->1	å->2	ö->1	
ma m	a->3	e->17	i->1	o->2	ä->1	å->5	ö->2	
ma n	a->1	i->1	ä->4	å->3	
ma o	c->4	m->7	r->5	s->1	
ma p	a->1	e->2	o->5	r->6	u->1	å->9	
ma r	e->9	i->5	o->1	ä->2	
ma s	a->13	i->3	k->4	l->1	n->1	o->10	t->55	u->1	v->2	y->2	ä->18	å->1	
ma t	e->1	i->12	y->2	
ma u	n->1	p->2	t->12	
ma v	a->6	i->5	ä->1	å->2	
ma ä	r->3	
ma å	r->2	s->1	t->2	
ma ö	v->9	
ma, 	a->1	d->3	f->2	m->1	o->1	s->1	u->1	
ma.D	e->1	
ma.H	e->2	
ma.J	a->4	
ma.O	m->1	r->1	
ma.V	i->1	
ma: 	a->1	u->1	
mace	u->1	
mad 	o->1	
made	 ->9	s->1	
maff	ä->1	
mage	 ->1	r->1	
magh	 ->1	
magi	n->1	
magn	a->1	i->1	
mago	g->4	
mail	 ->1	
main	s->7	
maj 	1->3	2->1	f->1	
maj,	 ->1	
maj.	J->1	T->1	
majo	r->41	
mako	l->1	
makr	o->6	
makt	 ->15	,->2	.->5	b->4	d->2	e->8	f->1	h->2	k->1	l->3	m->3	
makä	m->1	
mal 	b->2	e->2	f->1	p->1	s->1	
mala	 ->6	y->1	
mali	s->4	t->1	
malt	 ->5	.->3	e->3	
man 	"->1	E->1	F->1	I->2	R->1	a->35	b->31	d->25	e->13	f->30	g->20	h->40	i->88	j->5	k->40	l->16	m->36	n->15	o->23	p->14	r->14	s->87	t->32	u->17	v->38	y->1	ä->15	å->6	ö->7	
man!	 ->224	A->1	D->2	E->2	J->6	M->1	S->1	T->2	U->1	V->2	
man,	 ->171	
man.	D->1	H->1	K->1	M->1	S->1	
man:	 ->1	
mana	 ->13	d->2	r->32	s->4	t->3	
manb	i->1	l->2	o->1	r->1	u->1	
mand	a->23	e->80	i->1	r->1	
mane	n->8	r->1	
manf	a->14	ö->1	
mang	 ->11	,->1	.->4	e->4	
manh	a->47	ä->1	å->53	
mani	f->1	n->28	s->3	t->2	
manj	ä->1	
mank	a->9	o->3	
manl	a->1	i->1	ä->1	
mann	 ->2	,->1	-->1	a->2	e->24	i->2	
mano	 ->2	
mans	 ->32	,->3	.->1	;->1	a->3	k->9	l->7	m->1	t->6	v->1	ä->5	
mant	r->38	
manö	v->1	
mapl	a->1	
mar 	B->2	P->1	R->1	a->2	e->2	f->5	i->7	k->2	n->3	o->9	p->2	s->5	t->1	u->1	ö->2	
mar!	 ->1	
mar,	 ->14	
mar.	B->1	H->1	J->2	
marb	e->88	
mare	 ->38	,->4	.->5	n->37	
marg	i->6	
mari	t->3	
mark	 ->23	,->3	.->4	a->3	e->9	n->187	o->1	s->2	
marl	e->1	
marn	a->26	
mars	 ->5	,->3	.->2	c->1	
mas 	a->2	b->1	f->1	o->1	p->3	r->1	s->2	u->1	ö->1	
mas,	 ->1	
mask	e->2	i->6	u->1	
maso	c->1	
mass	a->5	i->3	m->3	
mast	 ->1	,->1	e->12	o->1	
mat 	a->2	e->1	f->2	s->2	u->6	v->1	
mat.	D->1	
matc	h->2	
mate	m->1	r->28	t->7	
matf	ö->4	
mati	,->1	k->5	o->72	s->38	v->2	
matn	y->1	
matp	e->1	r->1	
mats	 ->2	
matt	a->3	n->1	
matu	m->1	
mavt	a->3	
maxb	e->1	
maxi	m->7	
mb h	a->1	
mb.A	n->1	
mbad	s->1	
mbal	a->1	
mban	d->47	
mbar	 ->1	a->1	d->1	g->1	
mbas	s->1	
mbat	t->2	
mbed	s->1	
mben	 ->1	i->3	
mber	 ->31	,->9	.->6	v->1	
mbes	ö->2	
mbet	e->5	s->3	t->2	
mbex	p->1	
mbin	a->1	
mbit	i->26	
mble	m->1	
mbli	c->5	
mbni	n->1	
mbol	 ->2	i->7	
mbor	d->1	
mbro	t->2	
mbry	o->1	
mbud	 ->2	s->10	
mbul	a->1	
mbur	g->8	
mbus	 ->1	
mbyg	d->1	
mbär	l->4	
md a	t->1	
md h	ö->1	
md i	n->1	
md o	m->1	
md t	i->2	
md v	i->1	
md, 	e->1	h->1	
mda 	a->1	m->1	o->1	r->1	v->1	å->3	
mda,	 ->1	
mde 	T->1	i->1	m->2	s->1	
mde.	D->1	
mdef	i->1	
mden	 ->1	
mdes	 ->1	
mdhe	t->1	
mdir	i->1	
mdri	v->6	
mdöm	e->2	
me e	g->1	
me f	å->1	ö->5	
me k	o->1	
me o	c->2	m->1	
me s	o->4	
me å	t->2	
me, 	d->1	
me-f	a->1	
me.K	o->1	
med 	"->3	-->1	1->6	2->8	3->2	5->1	8->1	A->3	B->2	D->2	E->19	F->4	G->1	H->4	I->3	J->1	K->2	L->3	M->4	O->2	P->1	R->1	S->5	T->3	U->4	V->2	a->195	b->23	d->250	e->136	f->89	g->19	h->52	i->40	j->3	k->58	l->14	m->68	n->38	o->48	p->50	r->38	s->122	t->75	u->30	v->52	y->5	Ö->2	ä->9	å->6	ö->15	
med,	 ->14	
med.	D->3	F->1	V->2	
meda	n->23	r->2	
medb	e->15	o->168	r->1	
medd	e->59	
mede	l->217	
medf	i->2	ö->20	
medg	e->18	i->2	ö->2	
medh	j->1	
medi	a->8	c->1	e->5	n->1	
medk	ä->5	
medl	a->3	e->347	i->4	
medv	e->61	
mega	p->1	
meka	.->1	n->10	
mell	 ->1	a->211	e->67	i->1	t->11	
mels	 ->1	e->145	
men 	(->1	-->3	A->1	C->1	E->1	F->1	I->1	K->2	L->1	a->23	b->11	d->97	e->13	f->75	g->2	h->6	i->39	j->40	k->6	l->1	m->24	n->11	o->49	p->4	r->5	s->33	t->13	u->4	v->46	ä->15	ö->2	
men,	 ->26	
men.	D->5	F->1	H->1	J->5	L->1	M->1	O->1	U->1	V->1	
men;	 ->2	
men?	V->1	
mena	d->2	n->2	r->27	s->2	
mend	a->33	e->12	
mene	r->3	t->2	
meni	n->53	s->2	
mens	 ->10	a->196	b->2	i->13	k->194	
ment	 ->153	,->21	.->19	a->56	e->557	f->6	k->1	o->1	p->2	r->1	s->40	t->1	v->2	ä->2	
mer 	-->4	2->2	6->1	B->2	E->4	G->1	I->3	J->2	N->1	S->1	T->1	a->433	b->9	d->61	e->23	f->51	g->8	h->11	i->48	j->15	k->28	l->10	m->30	n->15	o->84	p->23	r->7	s->46	t->17	u->11	v->49	ä->42	å->2	ö->6	
mer!	"->2	
mer,	 ->15	
mer.	 ->2	B->1	D->8	F->1	H->1	I->2	J->1	K->1	M->1	O->1	S->1	T->1	V->6	
mera	 ->39	d->7	n->1	r->4	s->5	y->1	
merf	o->22	
merg	e->1	
meri	k->17	n->18	t->1	
mern	a->22	
merp	a->1	
mers	 ->1	a->1	i->7	
merv	ä->5	
mes,	 ->1	
mesg	i->1	
mest	 ->39	a->5	e->4	
met 	"->2	(->1	-->4	A->2	K->2	L->1	S->1	a->4	b->5	e->4	f->29	g->4	h->4	i->10	k->2	l->2	m->25	n->1	o->5	p->4	s->14	t->3	u->1	v->3	ä->19	
met)	 ->2	.->1	
met,	 ->15	
met.	 ->1	1->1	B->1	D->4	E->1	H->2	I->3	J->6	M->4	N->1	O->1	P->1	V->2	
met:	 ->1	
met?	K->1	
meta	l->11	
mete	r->5	
meto	d->29	
metr	a->1	
mets	 ->3	
meur	o->4	
mexi	s->2	
mfar	t->1	
mfat	t->83	
mfin	a->1	
mfly	t->1	
mfor	m->3	s->1	
mfun	d->5	
mfäl	l->1	
mfån	g->2	
mför	 ->108	a->143	b->11	d->42	e->2	h->2	k->1	s->23	t->30	
mger	 ->1	
mgic	k->2	
mgiv	a->1	n->1	
mgri	p->4	
mgän	g->1	
mgå 	e->1	i->1	
mgå.	F->1	
mgåe	n->1	
mgån	g->43	
mgår	 ->15	.->1	
mgåt	t->3	
mhet	 ->58	,->6	.->7	?->1	e->21	s->7	
mhul	d->1	
mhäl	l->49	
mhär	d->1	
mhäv	a->3	e->1	
mhål	l->17	
mhög	e->14	
mhöl	l->2	
mi -	 ->1	
mi a	t->1	
mi m	e->5	
mi o	c->12	
mi ä	r->1	
mi, 	l->1	m->1	v->1	
mi.D	e->2	
mi.F	ö->1	
mi? 	O->1	
mibe	s->2	
midd	a->13	
midi	g->3	s->1	
mier	 ->1	,->1	.->1	n->5	
mifi	n->1	
mig 	a->39	b->9	d->8	e->6	f->13	g->4	h->5	i->15	k->3	l->2	m->10	n->5	o->25	p->11	r->1	s->12	t->8	u->5	v->12	y->1	ä->8	å->6	ö->2	
mig!	"->1	
mig,	 ->15	
mig.	D->1	E->1	J->3	
mig:	 ->1	
mig?	V->1	
miga	,->1	
migh	e->2	
migr	a->10	e->1	
migt	 ->1	
miin	n->1	
mik 	e->1	o->1	
mika	l->5	p->1	
miko	n->1	
mikr	a->2	o->4	
mild	a->1	r->3	
mili	a->1	s->1	t->8	
milj	 ->1	a->15	e->14	o->63	ö->189	
mill	e->7	
mils	t->1	
milä	n->1	
milö	n->1	
min 	-->1	a->2	b->5	d->6	e->5	f->14	g->23	i->3	k->27	m->19	o->13	p->5	r->8	s->7	t->5	u->15	v->2	å->9	ö->2	
min,	 ->3	
min.	C->1	D->1	L->1	M->1	V->1	
mina	 ->72	l->4	n->1	r->1	t->2	
mind	e->1	r->52	
mine	l->3	r->44	
ming	 ->4	"->1	)->3	
mini	m->27	r->1	s->95	v->1	
minn	a->23	e->21	s->6	
mino	r->24	
mins	 ->3	k->63	t->58	
minu	s->5	t->16	
minä	r->3	
mipa	r->1	
mira	k->1	
mire	f->2	g->3	
mis-	f->1	n->1	
mis.	F->1	
misk	 ->49	.->1	a->145	t->28	
mism	 ->3	e->2	
miss	 ->7	,->5	.->2	a->3	b->10	e->1	f->7	g->7	h->1	i->1151	k->6	l->19	n->3	r->2	t->24	u->2	
mist	e->4	i->11	l->1	y->4	
misä	r->2	
mit 	d->1	e->2	f->7	h->1	i->2	m->5	n->2	t->6	u->4	v->1	ö->6	
mit,	 ->3	
mit.	M->1	P->1	
mita	 ->1	
mite	t->7	
miti	s->3	v->1	
mitn	i->1	
mitr	a->5	
mits	 ->2	
mitt	 ->68	a->1	e->2	é->59	
mium	 ->2	,->1	
mix.	D->1	
mixe	n->1	
miär	m->10	
miål	d->1	
mja 	a->2	d->4	e->8	f->3	g->2	h->1	i->1	k->4	l->2	p->1	s->4	v->1	y->1	å->2	
mja.	K->1	
mjan	d->17	
mjar	 ->6	
mjas	,->1	
mjat	 ->1	
mjuk	a->1	n->2	
mka 	i->1	
mkar	 ->2	
mkas	t->1	
mkat	 ->1	,->1	
mkom	m->10	
mkri	n->15	
mla 	U->1	b->7	d->1	f->6	h->1	i->5	k->5	l->1	m->2	o->1	r->1	s->5	t->1	u->1	
mlad	e->2	
mlag	d->3	t->9	
mlan	d->3	
mlar	 ->2	f->1	
mlas	 ->1	t->1	
mlat	 ->3	s->2	
mlen	,->1	
mlev	n->1	
mlig	 ->5	.->1	a->18	e->48	g->1	h->19	t->21	
mlik	 ->1	h->12	
mlin	g->59	
mlok	a->2	
mläg	g->8	
mlän	d->1	
mläs	n->2	t->1	
mläx	o->1	
mlös	a->2	h->3	
mm a	v->1	
mma 	-->1	1->1	E->1	a->22	b->10	d->18	e->9	f->23	g->3	h->8	i->45	j->5	k->14	l->7	m->28	n->9	o->11	p->21	r->16	s->101	t->14	u->13	v->11	ä->3	å->4	ö->8	
mma,	 ->7	
mma.	H->1	J->3	O->1	
mma:	 ->2	
mmad	 ->1	e->4	
mmal	 ->4	
mman	 ->20	,->1	.->1	b->6	d->69	f->15	h->101	j->1	k->12	l->2	s->57	t->35	
mmap	l->1	
mmar	 ->18	!->1	,->8	.->1	e->64	l->1	n->3	
mmas	 ->6	,->1	
mmat	 ->4	e->1	s->1	
mme 	e->1	f->6	k->1	o->3	s->4	å->2	
mme,	 ->1	
mmel	s->143	
mmen	 ->25	,->6	.->10	;->1	d->45	t->37	
mmer	 ->761	,->6	.->6	f->22	s->9	
mmet	 ->56	)->2	,->6	.->12	:->1	s->2	
mmig	a->1	h->2	r->7	t->1	
mmip	a->1	
mmis	s->1150	
mmit	 ->37	,->3	.->2	s->2	t->59	
mmon	 ->1	
mmor	 ->8	,->1	.->1	
mmun	.->1	a->3	e->10	i->20	
mmöb	l->1	
mn K	o->1	
mn b	y->1	
mn i	 ->1	
mn k	a->1	
mn m	e->1	å->2	
mn o	c->1	
mn p	å->1	
mn s	o->1	p->1	v->1	
mn, 	f->1	m->1	u->1	
mn.D	e->2	
mn.M	e->1	
mn.V	i->1	
mna 	A->1	L->1	a->4	b->1	d->9	e->7	f->5	g->1	h->5	i->8	k->1	m->2	n->1	o->2	p->2	r->3	s->7	t->5	u->3	v->2	
mna,	 ->2	
mna.	T->1	
mnad	 ->1	e->9	
mnan	d->4	
mnar	 ->61	.->3	e->4	n->6	
mnas	 ->12	,->2	
mnat	 ->13	s->5	
mnav	g->2	
mnbe	s->1	
mnda	 ->7	s->1	
mnde	 ->11	,->4	.->2	s->1	
mne 	h->1	i->1	s->1	
mne.	D->2	
mne:	 ->1	
mnen	 ->12	,->2	.->6	a->1	
mner	 ->4	.->1	
mnet	 ->4	.->2	
mnin	g->84	s->1	
mnko	n->2	
mns 	a->1	e->1	f->1	h->1	i->1	m->1	o->1	u->1	
mns.	D->1	
mnt 	b->1	e->1	f->1	g->1	i->1	k->1	l->1	n->1	p->1	
mnt,	 ->2	
mnt.	D->2	
mnts	 ->2	,->2	.->2	
mnup	p->4	
mnvi	k->1	
mnvä	r->1	
mo, 	H->1	d->1	
mobi	l->7	
moco	,->1	
mod 	a->1	e->1	f->1	i->1	m->1	s->1	ä->1	
mode	l->12	r->40	t->6	
modi	f->3	g->4	
modl	i->12	
mofo	b->1	
moge	n->3	t->1	
mogr	a->3	
moko	 ->5	
mokr	a->137	
moln	 ->1	
mome	n->5	
momr	å->3	
moms	p->1	
mon 	l->1	
monb	e->1	
mone	t->7	
moni	 ->1	s->17	t->1	
monn	ä->1	
mono	k->3	p->17	
mons	t->7	
mont	e->12	
mor 	a->1	b->1	o->1	p->3	s->1	u->1	
mor,	 ->1	
mor.	V->1	
mora	l->7	
mord	 ->3	,->1	.->1	b->1	e->8	i->1	n->38	
morg	a->2	o->37	
mors	e->6	
moru	m->1	
mos 	O->1	
mose	x->1	
moso	r->1	
mot 	-->2	1->1	5->1	A->1	D->1	E->9	F->3	G->1	H->3	I->1	J->3	L->1	M->1	R->2	S->1	T->2	U->1	W->1	a->35	b->21	d->60	e->26	f->14	g->2	h->9	i->10	k->8	l->2	m->11	n->7	o->7	p->7	r->9	s->26	t->4	u->3	v->16	y->1	Ö->3	ä->2	å->1	ö->6	
mot!	 ->7	
mot,	 ->17	
mot.	 ->1	F->2	V->1	
mota	r->1	
mote	n->26	
motg	å->1	
moti	o->1	v->21	
moto	r->9	
motp	a->4	
mots	a->23	t->16	v->17	ä->17	
mott	a->17	
motv	e->4	i->2	
motå	t->3	
mout	i->1	
mp J	ö->1	
mp a	t->2	
mp f	ö->2	
mp i	 ->3	
mp m	e->1	o->4	
mp s	j->1	
mp.D	e->1	
mpa 	-->1	a->7	b->3	d->12	e->4	f->12	g->3	i->1	k->5	m->1	n->1	o->2	p->5	r->2	s->6	t->1	u->2	å->1	
mpad	 ->2	
mpag	n->1	
mpak	e->1	
mpan	d->4	j->6	
mpar	 ->12	.->1	
mpas	 ->34	,->1	.->8	:->1	s->1	
mpat	 ->3	i->8	s->5	
mpel	 ->72	,->5	.->3	:->3	v->28	
mpen	 ->14	,->1	.->1	s->10	
mper	a->6	i->3	
mpet	e->11	
mpic	 ->1	
mpis	k->1	
mpla	n->9	r->2	
mple	m->11	n->3	t->17	x->4	
mpli	c->12	g->60	m->4	n->1	
mpni	n->85	
mpon	e->7	
mpop	u->1	
mpor	,->1	t->6	ä->2	
mpro	c->10	g->15	j->1	m->22	
mprö	v->8	
mpso	n->1	
mpto	m->1	
mpul	s->6	
mpun	k->1	
mpål	e->1	
mra 	e->1	i->1	k->1	
mrad	 ->7	e->4	
mran	d->1	
mrap	p->2	
mrar	 ->3	
mras	 ->1	.->1	
mrat	 ->2	
mre 	b->1	f->2	h->1	l->1	s->1	
mres	t->1	
mrin	g->1	
mrum	 ->1	,->1	
mrun	d->1	
mrät	t->1	
mråd	 ->3	,->1	.->1	a->2	e->317	s->1	
mrös	t->57	
ms B	l->1	
ms a	n->2	
ms e	f->2	
ms f	ö->1	
ms i	 ->1	
ms s	ä->1	
ms t	u->1	
ms u	t->1	
ms v	a->1	
ms- 	o->3	
ms-,	 ->1	
msa 	d->2	u->1	
msan	 ->1	.->1	
msar	 ->1	
msav	t->2	
msbe	t->2	
msbr	o->1	
mses	i->5	
msfr	å->3	
msfu	l->1	
msgr	ä->1	
msha	v->1	
mshe	m->1	
msid	e->1	
msig	n->2	
msk 	k->1	
mska	 ->3	n->1	p->2	s->1	
mski	n->1	
mskj	u->1	
mskr	i->1	
msky	d->4	
msla	g->3	n->9	
mslu	t->3	
mslä	n->27	
msni	t->11	
msol	l->1	
msor	g->9	
mspa	r->1	
mspl	i->1	
mspä	n->1	
msre	g->1	
msrä	t->1	
msrå	d->2	
msst	a->284	
mst 	I->1	a->2	d->2	e->2	f->1	g->2	i->6	k->3	l->3	m->1	o->4	p->5	s->1	t->2	u->3	v->7	ö->1	
mst.	F->1	
msta	 ->13	d->1	
mste	g->32	n->2	r->45	
mstf	ö->1	
msth	ä->1	
mstk	ä->1	
msto	l->86	
mstr	a->1	i->4	u->10	
mstä	l->35	m->5	n->34	
mstå	 ->1	e->5	r->1	
mstö	t->1	
msve	p->1	
msvä	t->1	
msyn	 ->2	,->1	
msyr	a->3	
msät	t->8	
msåt	g->1	
mt A	u->1	
mt G	a->1	
mt H	e->1	
mt W	a->1	
mt a	l->1	n->2	r->1	s->1	t->14	v->3	
mt b	a->1	e->3	i->1	o->1	ö->1	
mt d	e->3	
mt e	k->3	n->2	r->1	t->3	u->2	
mt f	a->1	o->1	r->3	ö->9	
mt h	a->1	å->3	
mt i	 ->3	n->2	
mt j	ä->1	
mt k	o->3	u->1	v->1	
mt l	u->1	ä->2	
mt m	e->1	i->1	o->1	y->1	å->2	
mt n	e->1	
mt o	c->5	m->10	
mt p	a->2	o->1	å->1	
mt r	a->1	e->3	y->1	ä->2	
mt s	a->1	i->4	k->1	t->6	y->1	
mt t	a->6	i->4	
mt u	n->2	p->2	t->5	
mt v	a->2	i->1	ä->1	
mt y	t->1	
mt ä	n->1	v->2	
mt å	t->1	
mt ö	k->1	v->2	
mt, 	f->2	g->1	v->1	ä->2	
mt.D	e->1	
mt.P	å->1	
mt.U	n->1	
mt.Å	r->1	
mta 	s->2	u->1	
mtag	a->3	i->1	n->1	
mtal	 ->4	a->2	e->9	s->2	
mtan	d->1	k->1	
mtar	 ->1	
mtas	 ->1	
mtat	 ->1	
mte 	F->1	b->1	d->1	h->1	k->1	p->2	r->6	v->1	
mted	e->2	
mtid	 ->7	,->3	.->6	:->1	a->22	e->64	i->67	s->4	
mtie	l->1	
mtio	 ->1	e->1	n->2	
mtli	g->25	
mtni	n->1	
mton	 ->5	
mträ	d->2	
mts 	a->2	i->1	
mtsa	m->1	
mtvi	n->2	
mtyc	k->6	
mtän	k->1	
mtål	i->1	
mugg	l->1	
mula	 ->1	n->4	t->3	
mule	r->26	
mull	,->1	
mult	i->9	
mum 	-->1	a->1	m->1	p->1	
mun.	D->1	
muna	l->3	
mune	r->10	
muni	c->2	k->16	s->1	t->1	
munt	l->8	r->21	
mura	r->1	
mus 	e->1	
mus-	b->1	
musi	k->4	
muss	e->2	l->1	
mutf	o->1	
muto	r->1	
muts	a->2	i->1	
mvan	d->5	
mver	k->4	
mvet	e->1	s->1	
mvik	t->2	
mvil	l->3	
mvis	t->1	
mväg	 ->1	e->1	
mväl	v->4	
mvän	d->4	t->1	
mvär	d->1	
mväx	l->1	
myck	e->452	
mygg	o->1	
myll	r->1	
mynd	a->1	i->161	
mynn	a->2	
myti	s->1	
mán,	 ->1	
mäde	l->1	
mäkt	a->1	i->2	
mäla	 ->2	n->1	
mäld	a->1	
mäle	r->1	
mäln	i->12	
mäls	 ->2	
mält	 ->1	n->1	
män 	a->2	d->2	e->2	f->4	g->3	h->1	i->5	l->1	n->1	o->13	p->3	r->2	s->12	t->4	u->2	å->6	
män,	 ->1	
män.	I->1	J->1	T->1	
mänd	r->3	
mäng	d->22	i->1	
mänh	e->47	
mäni	e->1	
männ	a->39	e->29	i->93	y->2	
mäns	 ->4	k->42	
mänt	 ->16	,->1	
märk	a->4	b->3	e->19	l->4	n->13	s->54	t->32	
märr	e->1	
märt	a->1	s->1	
mäss	i->31	
mäst	a->2	
mäta	 ->2	r->1	s->1	
mäte	r->1	
mäti	g->1	
mätt	a->1	e->2	
må E	u->1	
må a	n->1	
må b	e->1	l->1	
må e	k->1	
må f	a->1	r->1	ö->2	
må h	a->1	e->1	
må l	ä->2	
må m	e->2	ä->1	ö->1	
må o	c->33	
må p	l->1	
må r	å->1	
må s	p->1	t->4	
må v	a->1	
må å	t->1	
må, 	m->1	s->1	
må.D	e->1	
måen	d->2	
måfö	r->6	
måga	 ->19	,->2	.->2	n->8	
mågr	ä->1	
måhä	n->5	
mål 	(->1	1->16	2->10	5->2	a->3	b->2	e->1	f->20	g->1	h->2	i->5	j->1	l->1	n->1	o->8	p->2	r->1	s->15	t->1	u->2	ä->4	
mål,	 ->16	
mål-	2->1	
mål.	B->1	D->3	E->1	F->1	H->2	I->2	J->1	K->1	M->2	N->2	Ä->1	
mål:	 ->1	
måla	r->1	
måle	n->15	t->28	
måli	g->1	n->4	
målm	e->1	
måls	d->1	e->2	s->1	ä->17	
mån 	b->1	d->5	f->11	h->1	l->1	o->1	s->2	
mån,	 ->1	
måna	 ->3	d->71	
månd	a->3	e->1	
måne	r->2	
mång	a->141	f->17	s->3	
måni	n->4	
måns	p->1	
mår.	H->1	L->1	
måri	g->1	
mårs	p->2	
måsk	a->1	
måst	e->696	
måt 	i->5	m->3	o->2	p->1	v->1	
måt,	 ->3	
måt.	D->3	F->1	H->1	J->1	V->1	
måtg	ä->1	
mått	 ->1	.->1	f->1	o->2	
mé o	c->2	
mé p	e->1	
méav	t->1	
méko	n->1	
mén 	o->1	
mén.	W->1	
més 	R->1	
möbl	e->2	
möda	 ->3	
mödo	s->1	
mödr	a->1	
möge	l->1	
mögn	a->1	
möjl	i->307	
möns	t->2	
mör 	s->1	v->1	
mörd	a->5	
mörk	 ->1	l->1	
möss	o->1	
möta	 ->10	
möte	 ->13	n->4	r->87	s->5	t->21	
möts	 ->2	
mött	e->1	
möve	r->2	
n "E	u->1	
n "L	o->1	
n "T	i->2	
n "d	e->1	ö->1	
n "e	n->1	u->2	
n "h	e->1	
n "n	o->1	
n "r	e->2	
n "s	p->1	
n "u	t->1	
n "å	t->1	
n (1	4->2	9->1	
n (A	5->5	
n (B	5->2	
n (C	E->2	
n (E	I->1	
n (F	U->1	
n (H	-->21	
n (I	M->1	
n (K	O->1	
n (e	l->1	
n (f	o->1	ö->2	
n (i	n->1	
n (m	a->1	
n (o	c->1	
n (s	å->1	
n , 	b->1	
n - 	"->1	'->1	2->1	6->1	A->1	R->1	a->4	b->2	d->9	e->6	f->3	h->5	i->3	j->2	l->2	m->3	n->1	o->8	s->6	t->2	u->2	v->3	Ö->1	ä->3	ö->1	
n 1 	j->6	m->2	o->2	p->2	s->1	
n 1,	 ->1	
n 10	 ->2	0->4	5->1	
n 11	 ->2	
n 12	/->3	4->2	6->1	
n 13	 ->3	,->1	
n 14	 ->7	
n 15	 ->2	0->1	
n 16	 ->2	
n 17	 ->3	,->1	
n 18	 ->5	
n 19	 ->1	1->1	4->1	6->5	7->1	8->3	9->30	
n 2 	d->1	o->1	
n 2,	 ->1	
n 20	 ->1	0->16	
n 21	 ->2	
n 23	 ->1	
n 24	 ->1	
n 26	 ->3	
n 28	 ->1	
n 29	,->1	
n 3 	f->1	j->1	m->1	o->1	
n 3,	 ->1	8->1	
n 30	 ->3	
n 31	 ->3	
n 34	.->1	
n 38	 ->1	
n 39	,->1	
n 4 	e->1	j->2	
n 4,	 ->2	
n 5 	0->2	o->1	
n 50	-->1	
n 52	0->1	
n 57	,->1	
n 6 	d->1	
n 7 	d->1	o->1	
n 79	/->1	
n 8 	o->2	
n 89	 ->1	
n 9 	d->1	f->1	
n 90	 ->1	
n 95	 ->1	
n AB	B->1	C->1	
n AD	R->1	
n Ac	t->1	
n Af	r->1	
n Al	b->1	t->2	
n Am	o->1	s->5	
n An	n->1	
n Ar	i->1	
n At	a->2	
n Au	t->1	
n BS	E->1	
n Ba	r->2	s->1	
n Be	l->1	r->3	
n Bo	e->1	n->1	
n Br	e->1	o->2	u->1	y->1	
n CE	N->4	
n Ca	n->1	s->1	
n Ce	n->1	
n Ch	a->1	
n Cr	e->2	
n Da	l->1	m->2	n->1	
n De	 ->6	
n Du	i->1	
n EG	-->3	
n EK	S->1	
n EM	U->1	
n EU	 ->1	,->1	-->1	:->2	?->1	
n Ei	e->1	
n En	 ->1	l->2	
n Er	i->6	
n Eu	r->50	
n FE	O->1	
n FM	I->1	
n FN	,->1	
n Fl	o->4	
n Fo	l->1	n->1	
n Fr	a->2	
n Fö	r->2	
n GU	E->1	
n Ga	l->1	r->1	z->1	
n Go	l->1	r->1	
n Gr	a->1	e->1	u->1	
n Gö	t->1	
n Ha	i->2	r->2	
n He	l->2	
n Hu	l->23	
n I 	-->1	o->1	
n IM	O->1	
n IR	A->1	
n IX	,->1	
n Im	b->2	
n In	d->1	t->2	
n Is	a->2	r->12	
n Ja	c->2	p->1	
n Jo	r->1	
n Ju	g->1	n->1	
n Ka	l->2	r->3	
n Ki	n->4	
n Ko	c->4	m->1	r->1	s->1	
n Ky	o->2	
n Kö	l->1	p->1	
n La	n->3	
n Le	a->1	
n Li	s->1	
n Lo	i->1	y->1	
n Ma	r->1	
n Mi	n->1	
n Na	t->5	
n Ni	e->1	
n No	i->1	
n OS	S->1	
n PP	E->2	
n PR	-->1	
n PS	E->1	
n Pa	l->2	r->1	
n Pl	a->1	
n Po	l->1	r->4	
n Pr	o->7	
n Ra	n->2	
n Re	d->2	
n Ro	t->1	v->2	
n SP	Ö->1	
n SS	 ->1	
n Sa	m->3	
n Sc	h->2	
n Se	b->1	
n Sh	a->2	
n So	l->1	
n Sy	d->1	r->4	
n Sã	o->1	
n Ta	m->4	
n Te	r->1	
n Th	e->1	
n To	t->1	
n Ty	s->4	
n UN	I->1	
n US	A->1	
n Un	i->2	
n VI	I->2	
n Va	l->3	
n Ve	l->1	n->1	
n Vi	v->1	
n Wa	l->1	
n Wi	e->4	
n Wo	g->18	
n Wu	r->1	
n XX	V->1	
n a 	p->1	
n ab	s->4	
n ac	c->15	
n ad	e->1	m->5	r->1	v->1	
n ag	e->3	r->1	
n ak	t->12	
n al	b->2	d->4	l->65	
n am	b->2	e->3	
n an	 ->1	a->11	b->1	d->73	g->11	i->3	l->24	m->5	n->40	o->2	p->1	s->47	t->13	v->17	
n ap	p->2	
n ar	a->2	b->22	k->1	t->5	
n as	p->7	y->1	
n at	t->429	
n au	k->2	t->1	
n av	 ->471	.->2	b->7	d->1	f->6	g->15	i->2	l->3	s->45	t->1	v->5	
n ax	e->1	
n ba	d->1	k->4	l->8	n->4	r->23	
n be	a->7	d->14	f->17	g->25	h->24	k->15	l->8	m->6	n->1	r->20	s->37	t->42	u->1	v->6	
n bi	b->1	d->13	l->23	n->1	o->2	t->2	
n bl	a->8	e->4	i->24	o->3	
n bo	e->1	k->3	m->1	n->2	r->17	s->2	t->4	
n br	a->14	e->7	i->14	o->7	u->1	ä->2	
n bu	d->13	
n by	g->3	r->6	t->2	
n bä	r->5	s->6	t->17	
n bå	d->3	
n bö	r->56	
n ce	n->10	r->1	
n ch	a->6	e->2	o->1	
n co	n->1	r->1	s->4	
n da	g->22	m->1	n->7	
n de	 ->86	a->1	b->30	c->8	f->6	g->1	l->75	m->21	n->103	p->1	r->11	s->19	t->195	
n di	a->7	k->2	r->8	s->17	t->1	v->1	
n dj	u->7	ä->1	
n do	c->3	g->1	k->2	m->9	
n dr	a->9	i->2	o->1	u->3	y->1	ö->2	
n du	b->1	m->1	n->1	
n dy	k->1	n->1	
n dä	r->57	
n då	 ->16	l->1	v->1	
n dö	d->2	l->2	m->2	p->3	r->3	
n ef	f->24	t->31	
n eg	e->22	n->4	
n ej	 ->2	
n ek	o->55	
n el	e->3	l->36	o->2	
n em	e->6	i->1	
n en	 ->122	a->14	b->5	d->31	e->4	g->8	h->17	k->4	l->10	o->9	s->12	t->1	v->1	
n ep	o->1	
n er	 ->2	,->1	a->1	b->3	f->2	h->2	i->1	k->6	s->3	t->2	
n et	n->3	t->52	
n eu	r->145	
n ev	e->4	
n ex	 ->1	a->3	e->1	i->5	k->1	p->10	t->7	
n fa	k->7	l->4	n->2	r->9	s->12	t->9	
n fe	d->2	l->3	m->7	
n fi	c->3	l->1	n->39	
n fj	o->1	ä->6	
n fl	a->3	e->8	i->1	o->1	y->1	
n fo	k->1	l->2	n->4	r->33	
n fr	a->47	e->9	i->13	o->2	u->4	y->1	ä->4	å->159	
n fu	l->12	n->13	s->1	
n fy	l->1	r->3	s->2	
n fä	l->1	r->1	s->4	
n få	 ->20	,->1	n->1	r->24	s->1	t->1	
n fö	d->2	l->8	n->1	r->787	
n ga	m->8	n->7	r->20	v->1	
n ge	 ->16	d->1	m->100	n->51	o->1	r->6	s->2	t->2	
n gi	c->2	g->2	l->2	v->3	
n gj	o->14	
n gl	a->1	e->1	o->3	ä->9	
n gn	u->2	
n go	d->35	
n gr	a->15	e->5	i->1	u->57	ä->3	ö->1	
n gu	m->1	
n gy	n->1	
n gä	l->26	r->1	
n gå	 ->8	n->56	r->10	t->1	
n gö	r->51	
n ha	 ->11	d->17	f->7	l->8	m->4	n->26	r->321	v->1	
n he	b->1	j->2	l->43	m->4	r->1	
n hi	n->2	s->3	t->8	
n hj	ä->10	
n ho	n->1	p->10	r->1	s->10	t->6	
n hu	n->2	r->8	v->7	
n hy	p->1	s->1	
n hä	l->1	m->2	n->22	r->80	v->6	
n hå	l->17	r->4	
n hö	g->26	j->4	r->5	
n i 	A->5	B->9	C->2	D->2	E->34	F->5	G->4	H->3	I->5	K->13	L->9	M->8	N->2	O->1	P->1	R->2	S->12	T->9	V->2	W->2	a->21	b->12	c->2	d->106	e->28	f->58	g->8	h->9	i->4	j->2	k->9	l->8	m->30	n->1	o->7	p->16	r->14	s->56	t->5	u->19	v->26	z->1	Ö->14	ä->2	å->3	ö->1	
n i,	 ->1	
n ib	l->1	
n ic	k->4	
n id	e->6	é->4	
n if	r->3	
n ig	n->1	
n ih	ä->1	å->1	
n il	l->3	
n im	p->1	
n in	 ->1	b->4	c->1	d->7	e->2	f->33	g->7	h->3	i->1	k->2	l->9	n->29	o->50	r->70	s->29	t->250	v->5	
n ir	a->1	l->2	
n is	r->11	t->1	
n it	a->5	
n ja	g->130	k->2	n->1	
n ju	 ->4	b->1	l->2	n->1	r->7	s->15	
n jä	m->8	
n ka	b->1	l->5	m->6	n->143	p->1	r->2	s->2	t->17	
n ke	d->1	l->1	
n ki	n->1	
n kl	.->12	a->19	i->1	
n kn	a->3	
n ko	a->4	l->30	m->258	n->85	p->3	r->5	s->13	
n kr	a->11	i->12	ä->20	ö->1	
n ku	l->11	n->18	r->1	
n kv	a->4	i->4	o->6	
n ky	l->1	
n kä	l->3	n->16	r->2	
n kö	n->3	r->1	
n la	d->3	g->19	n->1	r->1	w->1	
n le	d->20	g->2	v->2	
n li	b->4	d->1	g->9	k->11	n->5	t->11	v->4	
n lo	g->2	k->8	v->3	
n lu	c->1	
n ly	c->8	d->1	s->4	
n lä	g->21	m->7	n->11	r->2	s->5	t->4	
n lå	g->3	n->20	t->3	
n lö	j->1	k->1	n->1	p->1	s->20	
n m.	m->1	
n ma	g->2	j->6	k->5	l->1	n->47	r->17	s->6	x->2	
n me	d->216	l->41	n->31	r->24	s->2	t->5	
n mi	l->18	n->43	s->13	t->1	
n mo	d->14	n->3	r->2	t->48	
n mu	l->1	n->3	
n my	c->69	n->12	
n mä	n->15	r->3	t->2	
n må	 ->2	h->1	l->3	n->14	s->139	
n mö	j->21	r->2	t->4	
n na	t->36	
n ne	d->7	g->5	u->1	
n ni	 ->13	o->1	v->3	
n no	g->1	l->1	m->2	r->5	t->5	
n nu	 ->28	,->1	m->1	v->16	
n ny	 ->25	a->38	c->2	e->1	h->1	l->5	n->1	s->4	t->8	
n nä	m->15	r->42	s->2	
n nå	 ->3	b->2	g->36	
n nö	d->15	j->1	t->1	
n oa	c->2	n->2	v->2	
n ob	a->1	e->21	l->5	
n oc	h->585	k->97	
n oe	g->1	n->1	r->2	
n of	a->1	f->26	t->2	ö->5	
n oh	ä->1	
n ok	l->2	o->1	ä->2	
n ol	i->8	j->2	y->7	
n om	 ->376	"->1	,->4	.->2	I->1	b->1	d->1	e->5	f->14	i->1	m->1	o->1	p->5	r->7	s->5	v->6	ö->4	
n on	d->1	e->1	ö->2	
n op	e->2	p->2	t->2	
n or	d->19	g->7	i->1	k->1	m->1	o->25	s->3	t->1	ä->1	
n os	s->6	
n ot	a->1	i->2	j->1	
n ou	m->2	n->1	
n ov	a->2	i->3	
n oä	n->1	
n oö	n->1	v->2	
n p.	g->1	
n pa	l->4	r->34	s->2	
n pe	d->1	k->2	l->2	n->1	r->27	t->1	
n pl	a->22	i->1	u->1	ö->2	
n po	e->1	l->57	o->1	r->5	s->15	t->1	ä->2	
n pr	a->2	e->14	i->12	o->30	
n pu	n->28	r->1	
n py	r->1	
n på	 ->239	:->1	?->1	b->1	f->1	g->5	m->3	p->6	s->6	t->2	v->5	
n ra	d->23	m->4	p->11	s->3	t->1	
n re	a->4	d->28	e->3	f->18	g->66	k->5	l->5	m->1	n->8	p->1	s->39	v->9	
n ri	g->1	k->20	m->3	s->17	
n ro	l->11	s->1	
n ru	n->2	s->1	
n ry	s->1	
n rä	c->2	d->4	k->7	t->48	
n rå	d->26	g->1	
n ré	f->1	
n rö	d->2	r->5	s->17	
n sa	d->17	g->9	k->22	m->47	n->5	t->8	
n sc	e->1	o->1	
n se	 ->12	d->10	g->2	k->2	n->12	p->1	r->19	t->2	x->1	
n si	f->1	g->12	n->11	s->20	t->23	
n sj	u->5	ä->29	
n sk	a->191	e->5	i->9	j->3	o->2	r->11	u->72	y->9	ä->3	ö->4	
n sl	a->4	o->1	u->22	å->1	
n sm	i->1	u->1	ä->2	å->1	
n sn	a->21	e->2	
n so	 ->1	c->41	l->6	m->353	r->6	
n sp	a->4	e->19	l->2	o->1	r->3	ä->1	
n sr	i->1	
n st	a->56	i->5	o->57	r->43	u->7	y->4	ä->26	å->24	ö->44	
n su	b->2	c->2	m->1	n->2	p->1	v->1	
n sv	a->6	e->2	å->3	
n sy	f->3	m->3	n->9	r->4	s->6	
n sä	g->25	k->9	l->2	r->17	t->5	
n så	 ->43	,->1	:->1	d->47	g->1	h->1	l->2	n->1	s->4	v->1	
n sö	d->2	k->1	
n t.	e->1	
n ta	 ->16	c->10	g->7	l->29	n->2	p->1	r->10	s->5	
n te	c->2	k->9	n->1	r->4	x->2	
n ti	b->4	d->43	l->316	m->1	o->1	t->6	
n tj	ä->8	
n to	g->4	l->2	m->1	n->2	p->2	t->11	
n tr	a->7	e->36	o->12	ä->4	ö->1	
n tu	f->1	n->5	r->9	
n tv	e->19	i->22	ä->5	å->7	
n ty	c->5	d->15	g->1	n->3	p->5	s->12	v->6	
n tä	n->9	v->1	
n un	d->79	g->1	i->15	
n up	p->106	
n ur	 ->5	m->1	s->6	v->1	
n ut	,->1	a->18	b->6	e->3	f->12	g->13	i->1	j->1	k->1	l->3	m->7	n->6	p->1	r->2	s->30	t->16	v->34	ö->5	
n va	d->16	l->10	n->6	r->87	t->1	
n ve	c->3	d->2	k->1	m->2	r->41	t->20	
n vi	 ->133	,->1	.->1	c->1	d->60	f->1	k->59	l->56	n->2	s->52	t->5	
n vo	l->1	r->3	
n vr	i->1	
n vu	n->1	
n vä	c->2	d->2	g->7	l->14	n->17	r->8	s->6	v->1	x->7	
n vå	g->1	l->4	r->13	
n wa	l->1	
n we	b->1	
n yt	t->8	
n zi	g->2	
n Ös	t->3	
n äg	a->3	e->1	n->4	t->1	
n äl	s->1	
n än	 ->11	d->31	n->10	t->1	
n är	 ->302	,->3	.->4	:->2	a->1	l->1	
n äv	e->32	
n å 	a->1	d->3	e->4	
n åb	e->1	
n åk	l->8	
n ål	a->1	d->2	ä->1	
n år	 ->9	l->1	
n ås	i->22	t->5	y->1	
n åt	 ->7	a->1	e->23	f->3	g->11	m->3	s->1	t->1	
n öd	e->1	
n ök	a->23	n->9	
n öm	 ->1	
n ön	s->9	
n öp	p->8	
n ör	e->1	
n ös	t->18	
n öv	e->74	n->2	r->4	
n! A	l->2	t->1	v->2	
n! B	e->2	
n! D	a->1	e->30	ä->1	í->1	
n! E	U->1	n->1	r->1	u->3	
n! F	r->3	å->1	ö->8	
n! G	r->2	
n! H	e->1	
n! I	 ->9	n->1	
n! J	a->75	
n! K	o->5	
n! L	i->1	å->5	
n! M	a->1	i->5	
n! N	i->1	u->1	ä->4	
n! O	l->1	m->1	
n! P	a->1	r->1	å->2	
n! R	e->1	o->1	å->2	
n! S	c->1	e->3	k->1	o->3	t->1	
n! T	a->1	h->1	i->4	o->1	r->1	
n! U	n->2	t->2	
n! V	a->3	i->12	å->2	
n! Ä	n->1	v->6	
n! Å	 ->3	
n! Ö	s->1	
n!Am	s->1	
n!De	n->1	t->2	
n!Ef	t->1	
n!En	 ->1	
n!He	r->1	
n!Ja	g->6	
n!Mi	n->1	
n!Nä	r->2	
n!Rö	s->1	
n!Sa	n->1	
n!Ta	c->1	
n!Ti	l->1	
n!Un	d->1	
n!Vi	 ->2	
n" a	l->1	t->1	
n" e	t->1	
n" g	e->1	
n" i	 ->1	
n" o	c->1	
n" p	å->1	
n" s	o->1	
n", 	"->1	d->1	o->1	s->2	
n".D	e->3	
n".O	r->1	
n".R	å->1	
n) (	K->2	S->1	
n) f	ö->1	
n) h	a->1	
n) z	o->1	
n)(P	a->2	
n), 	o->1	
n).D	e->2	
n).H	e->1	
n)Ja	g->1	
n)Nä	s->1	
n, "	o->1	
n, 1	 ->1	0->1	5->1	9->1	
n, 5	0->1	
n, 8	,->1	
n, A	m->2	
n, B	N->1	e->3	r->1	
n, C	u->1	
n, D	u->1	
n, E	u->2	
n, I	V->1	r->1	
n, J	o->1	
n, K	a->2	o->2	
n, L	o->2	
n, N	e->1	
n, O	l->1	
n, P	a->3	e->1	
n, R	a->1	o->1	
n, S	h->1	l->1	v->1	
n, T	o->1	y->1	
n, U	z->1	
n, V	 ->1	l->1	
n, W	i->1	
n, a	l->4	n->7	r->1	t->20	v->3	
n, b	a->3	e->1	l->6	o->1	r->1	ä->2	å->3	ö->5	
n, d	e->44	u->1	v->6	ä->14	å->3	ö->1	
n, e	f->19	k->1	l->5	n->16	t->11	x->1	
n, f	a->2	i->3	l->1	r->35	å->4	ö->55	
n, g	a->1	e->5	j->2	r->1	
n, h	a->14	e->57	o->1	ä->1	ö->1	
n, i	 ->21	g->1	n->29	
n, j	a->8	u->4	
n, k	a->6	o->19	r->2	u->1	v->1	ä->27	
n, l	i->5	ä->2	å->1	
n, m	a->2	e->55	i->19	u->1	ä->1	å->7	
n, n	a->1	u->1	ä->23	å->5	
n, o	c->118	f->1	m->15	s->1	
n, p	a->4	r->2	u->1	å->11	
n, r	a->1	ä->1	å->4	
n, s	a->11	e->1	k->13	l->2	n->2	o->79	t->3	ä->6	å->24	
n, t	.->3	a->4	i->13	r->5	v->3	y->4	
n, u	n->2	p->2	t->31	
n, v	a->10	e->1	i->45	o->1	ä->2	
n, y	t->1	
n, Î	l->1	
n, ä	g->1	n->2	r->27	v->14	
n, å	t->1	
n, ö	p->1	
n- o	c->4	
n-Cl	a->1	
n-Ha	r->1	
n-Ke	e->1	
n-SS	:->1	
n-gr	u->1	
n-rå	d->3	
n. D	e->7	ä->1	
n. F	o->1	
n. H	a->1	ä->1	
n. I	 ->1	n->1	
n. J	a->3	
n. L	å->1	
n. M	e->3	
n. N	ä->1	
n. O	c->3	
n. R	å->1	
n. V	i->2	
n." 	Ä->1	
n.(E	L->1	
n.(I	T->1	
n.(L	i->1	
n.(P	a->2	
n.) 	H->1	T->1	
n.).	H->1	
n.)A	n->1	
n.)B	e->4	
n.)F	r->3	
n.)G	e->1	
n.)H	e->1	
n.. 	(->9	D->1	
n..(	E->2	N->1	
n..H	e->1	
n.14	 ->1	
n.15	 ->1	
n.Al	l->11	
n.An	d->1	n->1	
n.Ar	b->1	t->1	
n.At	t->4	
n.Av	 ->6	s->2	
n.Be	d->1	t->2	
n.Bi	l->1	
n.Br	i->1	y->1	
n.Ce	n->1	
n.Cu	n->1	
n.DE	B->1	
n.De	 ->21	n->48	s->10	t->176	
n.Dä	r->28	
n.Då	 ->3	
n.EU	 ->2	
n.Ef	f->1	t->3	
n.Em	e->1	
n.En	 ->9	d->2	l->6	
n.Er	 ->1	i->1	
n.Et	t->10	
n.Eu	r->5	
n.Ev	e->1	
n.FE	O->1	
n.Fa	k->1	r->1	
n.Fi	n->1	
n.Fl	e->1	
n.Fo	r->1	
n.Fr	u->5	å->4	
n.Fy	r->1	
n.Fö	l->2	r->43	
n.Ge	n->1	
n.Go	l->1	
n.Gä	l->1	
n.Gå	 ->1	
n.Ha	d->1	n->5	r->2	
n.He	l->1	r->56	
n.Hi	t->2	
n.Ho	n->2	
n.Hu	r->5	
n.Hä	r->7	
n.I 	E->1	T->1	a->2	d->14	e->5	f->1	m->3	r->2	s->7	v->1	
n.Il	l->1	
n.In	g->2	o->1	r->1	s->1	t->2	
n.Ja	,->1	c->1	g->133	
n.Jo	r->1	
n.Ju	s->2	
n.Ka	n->5	
n.Ko	c->1	m->20	n->3	r->1	
n.Kr	a->1	
n.Ku	l->1	
n.Kv	a->1	
n.Le	d->1	
n.Li	k->1	v->1	
n.Lå	n->1	t->10	
n.Ma	n->6	r->1	x->1	
n.Me	d->5	n->35	
n.Mi	n->6	t->1	
n.Mo	t->4	
n.My	n->1	
n.Mä	n->1	r->1	
n.Må	n->1	
n.Mö	j->1	
n.Na	t->2	
n.Ni	 ->8	e->1	
n.Nu	 ->4	
n.Ny	l->1	
n.Nä	r->9	
n.Oc	h->10	k->1	
n.Om	 ->18	
n.Or	d->4	s->1	
n.Oz	 ->1	
n.Pa	r->4	
n.Pe	r->1	
n.Pl	a->1	
n.Pr	e->1	o->2	
n.På	 ->9	
n.Re	f->1	n->1	
n.Ri	k->1	
n.Ro	t->1	
n.Rä	t->1	
n.Rå	d->4	
n.Sa	m->5	n->2	
n.Sc	h->1	
n.Se	d->3	t->1	
n.Si	s->2	t->1	
n.Sk	a->1	u->1	
n.Sl	u->11	
n.Sn	a->1	
n.So	c->1	m->10	
n.St	a->1	å->1	ö->2	
n.Su	b->1	
n.Sy	f->2	
n.Sä	k->1	r->2	
n.Så	 ->7	l->1	
n.Ta	c->5	
n.Th	e->1	y->1	
n.Ti	d->1	l->5	
n.To	r->2	
n.Tr	o->3	
n.Tv	ä->1	
n.Ty	 ->2	v->3	
n.Un	d->8	i->2	
n.Up	p->1	
n.Ut	a->1	i->1	s->1	v->1	
n.Va	d->13	l->1	n->1	r->2	
n.Ve	t->1	
n.Vi	 ->85	d->4	l->5	s->2	t->2	
n.Vå	r->5	
n.Wo	r->1	
n.Än	 ->1	d->2	
n.Är	a->2	
n.Äv	e->4	
n.Å 	E->1	a->1	e->1	
n.Ög	o->2	
n.Öv	e->1	
n/No	r->2	
n/år	)->1	,->1	
n: "	d->1	
n: A	t->1	
n: D	e->2	
n: E	r->1	
n: H	a->1	
n: J	a->2	
n: K	o->3	
n: R	e->1	
n: T	å->1	
n: V	a->1	i->1	
n: a	t->1	
n: d	e->2	ä->1	
n: e	n->1	
n: f	o->1	ö->2	
n: i	 ->1	n->1	
n: j	a->1	
n: m	e->2	
n: n	ä->2	
n: v	a->3	i->2	
n:Fö	r->1	
n; J	a->1	
n; a	v->1	
n; d	e->9	ä->1	
n; e	n->1	
n; f	i->1	ö->1	
n; i	n->1	
n; m	e->1	
n; o	c->1	
n; p	u->1	
n; s	a->1	k->1	
n; v	i->1	
n; ä	n->1	
n? 2	1->1	
n? D	e->1	
n? I	n->1	
n?. 	(->1	
n?An	s->1	
n?De	n->3	s->1	t->4	
n?Ef	t->1	
n?Fo	l->1	
n?Fr	u->2	
n?Fö	r->2	
n?He	r->3	
n?Hu	r->1	
n?I 	d->1	
n?Ja	,->1	g->3	
n?Ka	n->3	
n?Ko	m->2	
n?Nä	r->1	
n?Om	 ->1	
n?Pa	r->1	
n?Se	d->1	
n?Va	d->1	
n?Ve	m->1	t->1	
n?Vi	 ->4	l->4	
n?Är	 ->4	
n?Äv	e->1	
nFrå	g->3	
nHer	r->2	
nI d	e->1	
nJag	 ->2	
nNäs	t->7	
na (	K->1	
na -	 ->23	
na 1	 ->2	2->1	3->1	6->1	
na 3	3->1	
na 6	 ->1	
na 8	1->4	5->3	7->1	
na A	l->1	z->1	
na B	 ->1	
na E	l->1	u->1	
na I	X->1	
na L	i->1	
na M	o->1	
na P	r->1	
na T	e->2	u->2	
na a	b->1	d->1	f->1	k->2	l->2	m->2	n->30	r->7	s->1	t->67	v->58	
na b	a->8	e->37	i->13	l->12	o->6	r->4	u->5	y->5	ä->1	ö->7	
na c	a->1	e->2	
na d	a->42	e->72	i->11	o->3	r->8	y->1	ä->12	å->3	ö->2	
na e	f->6	g->15	k->5	l->18	m->4	n->23	r->5	t->10	u->4	x->3	
na f	a->15	e->1	i->7	o->12	r->111	u->4	å->20	ö->210	
na g	a->9	e->38	i->2	j->3	l->1	o->1	r->19	ä->5	å->8	ö->16	
na h	a->56	e->6	i->1	j->2	o->6	u->4	y->1	ä->12	å->6	ö->5	
na i	 ->196	b->1	d->2	f->1	g->2	k->1	n->77	
na j	o->2	u->2	ä->1	
na k	a->40	l->3	n->1	o->81	r->5	u->7	v->7	ä->11	
na l	a->5	e->6	i->7	j->1	o->2	u->1	y->1	ä->8	å->2	ö->11	
na m	a->9	e->80	i->9	o->6	u->2	y->10	ä->3	å->24	ö->6	
na n	a->6	e->2	o->2	r->2	y->4	ä->9	å->7	
na o	b->1	c->170	f->1	j->1	l->4	m->75	p->2	r->15	s->9	
na p	a->10	e->6	l->3	o->8	r->35	u->10	å->41	
na r	a->8	e->78	i->8	o->2	ä->11	å->5	ö->7	
na s	a->8	e->20	i->42	j->10	k->59	l->10	m->2	n->3	o->64	p->11	t->46	u->2	v->3	y->8	ä->12	å->7	ö->2	
na t	.->1	a->20	e->8	i->61	j->2	o->6	r->7	v->6	y->14	ä->3	
na u	l->1	n->17	p->36	r->2	t->40	
na v	a->23	e->11	i->47	o->1	ä->12	å->6	
na y	r->2	t->2	
na ä	m->1	n->17	r->51	v->2	
na å	k->1	r->4	s->3	t->20	
na ö	d->2	g->2	k->3	n->2	p->1	s->1	v->11	
na!D	e->1	
na!H	e->1	
na!O	m->1	
na".	D->1	K->1	
na"i	n->1	
na, 	B->1	S->1	a->12	b->4	d->21	e->13	f->10	g->1	h->9	i->18	j->3	k->3	l->5	m->25	n->8	o->36	p->1	r->3	s->42	t->12	u->9	v->18	ä->2	ö->1	
na-I	s->1	
na. 	D->3	H->1	J->1	K->2	S->1	V->1	Å->1	
na.(	T->1	
na.)	B->1	
na.-	 ->2	
na..	(->1	
na.A	l->6	m->1	v->2	
na.B	e->2	
na.D	e->61	o->1	ä->6	
na.E	f->3	m->1	n->1	t->5	u->3	
na.F	a->2	r->1	ö->13	
na.G	e->1	i->1	
na.H	a->1	e->5	u->3	ä->2	
na.I	 ->12	b->1	n->3	
na.J	a->29	u->2	
na.K	a->2	o->8	
na.L	i->2	å->2	
na.M	a->1	e->13	i->5	
na.N	a->1	i->2	u->1	ä->3	
na.O	c->1	m->5	r->1	
na.P	r->1	å->4	
na.R	e->1	
na.S	e->1	k->1	l->3	o->3	t->1	y->1	å->2	
na.T	a->2	i->1	r->2	
na.U	n->2	p->1	r->1	t->4	
na.V	a->4	e->1	i->32	ä->2	å->1	
na.Ä	n->2	r->1	v->2	
na.Å	 ->1	
na/E	u->1	
na/s	a->1	
na: 	F->1	m->1	v->1	
na; 	j->2	l->1	o->1	p->1	
na?E	t->1	
na?H	a->1	u->1	
na?I	 ->1	
na?J	a->1	o->1	
na?M	a->1	
na?P	å->1	
na?S	v->1	
na?V	a->2	i->2	
na?Ä	r->1	
naHe	r->1	
nabb	 ->4	a->24	t->43	v->1	
nabi	s->1	
nack	a->2	d->8	
nad 	-->1	a->7	b->2	d->1	e->2	f->8	h->1	i->8	j->1	k->4	m->6	n->1	o->4	r->2	s->7	t->1	u->3	ö->1	
nad,	 ->11	
nad.	D->2	E->1	H->2	J->2	P->1	
nad:	 ->1	
nad;	 ->1	
nad?	H->1	V->1	
nada	,->2	
nade	 ->64	,->1	.->3	n->164	r->165	s->9	
nads	-->4	/->1	a->5	b->4	d->1	e->18	f->5	i->3	k->1	l->2	m->2	n->1	o->1	p->5	s->3	t->1	u->1	v->3	
nafl	y->1	
nafr	å->1	
naga	v->3	
nage	 ->1	l->1	r->1	t->1	
nagi	v->3	
naiv	a->1	i->1	
naki	s->2	
nakn	a->1	
nakr	y->1	
nal 	C->1	d->1	f->4	i->3	m->1	o->5	p->1	r->1	s->3	t->2	u->2	v->2	
nal,	 ->3	
nal-	s->2	
nal.	 ->1	D->1	F->1	P->1	S->1	V->1	
nala	 ->46	g->1	
nale	k->4	n->2	r->11	
nalf	a->1	ö->3	
nali	s->30	t->8	
nall	i->1	
nalp	a->1	o->40	r->1	
nalr	e->3	ä->1	
nals	o->1	t->5	y->1	
nalt	 ->1	
nalu	t->1	
nalv	e->1	
naly	s->58	
namb	a->1	
nami	k->1	s->4	
namm	a->4	
namn	 ->7	,->2	.->2	e->2	u->4	
nan 	E->3	a->3	b->3	c->1	d->11	e->2	f->3	g->1	h->1	i->6	j->3	k->1	m->8	n->1	o->3	p->1	r->3	s->9	t->1	v->16	å->2	
nan,	 ->4	
nan.	L->1	
nand	e->67	
nane	r->1	
nans	 ->2	d->1	e->2	i->79	l->1	m->1	t->2	v->1	
nant	 ->1	
napp	 ->1	a->11	n->1	t->5	
napr	o->2	
nar 	C->1	E->1	R->1	a->17	b->4	d->39	e->9	f->6	h->4	i->19	j->18	k->16	l->1	m->21	n->4	o->22	p->2	r->4	s->17	t->7	u->5	v->17	Ö->1	ä->2	å->2	ö->1	
nar,	 ->7	
nar.	.->1	D->4	H->2	M->1	O->1	S->2	U->1	V->1	
nar:	 ->1	
nara	r->24	s->13	
narb	e->1	
nard	 ->1	
nare	 ->35	,->5	.->5	l->1	n->5	p->1	
nari	e->1	o->4	u->1	
nark	o->7	
narl	i->1	
narn	a->17	
nars	 ->18	,->1	a->4	
nart	 ->26	.->1	
narå	d->1	
nas 	E->7	S->2	a->37	b->5	c->1	d->9	e->19	f->30	g->5	h->5	i->24	j->2	k->19	l->9	m->15	n->13	o->30	p->15	r->15	s->34	t->16	u->6	v->9	y->1	ä->2	å->4	ö->2	
nas!	E->1	
nas,	 ->10	
nas.	 ->1	D->3	E->1	J->1	K->1	M->1	V->1	Å->1	
nast	 ->13	?->1	e->63	å->2	
nat 	-->1	3->1	E->1	I->1	K->1	a->3	b->8	d->7	e->3	f->16	g->5	h->2	i->14	j->1	k->9	l->4	m->5	o->8	p->6	r->3	s->15	t->13	u->7	v->6	ä->13	å->3	ö->1	
nat,	 ->4	
nat.	 ->1	D->1	G->1	J->1	K->1	Ä->1	
nate	n->1	
nati	o->271	v->12	
nats	 ->11	,->2	.->2	
natt	 ->1	e->2	
natu	r->121	
naue	r->1	
navg	i->2	
navi	s->1	
navt	a->3	
nazi	s->16	
nban	a->1	
nbar	 ->1	.->2	a->1	l->12	n->1	t->51	
nbeg	r->12	
nbeh	a->1	
nber	 ->2	g->3	
nbes	t->1	
nbet	ä->5	
nbil	a->8	
nbin	d->1	
nbju	d->6	
nbjö	d->1	
nbla	n->16	
nbli	c->16	
nboe	n->1	
nbok	 ->1	e->1	
nbro	t->1	
nbry	t->1	
nbud	s->4	
nbul	 ->1	
nbun	d->1	
nbur	g->3	
nbyg	g->1	
nc d	å->1	
nc, 	d->1	
nca,	 ->1	
ncas	 ->1	
nce,	 ->1	
nce.	.->1	
ncen	t->31	
ncep	t->7	
ncer	!->1	,->1	a->1	b->1	n->2	
nche	n->1	z->1	
ncht	i->1	
ncid	e->1	
ncil	 ->1	
ncip	 ->28	,->3	.->4	e->151	i->8	s->1	
ncis	 ->2	t->1	
ncit	a->8	
nckh	e->14	
nd (	e->1	k->1	r->1	
nd -	 ->4	
nd 8	0->1	
nd E	U->1	
nd L	T->1	a->3	
nd S	v->1	
nd T	i->1	
nd a	c->1	l->4	n->22	t->11	v->80	
nd b	e->7	i->1	y->1	å->1	
nd c	i->1	
nd d	e->17	ä->5	
nd e	f->1	l->3	n->9	r->2	
nd f	i->1	o->1	r->6	y->1	ö->26	
nd g	e->3	o->1	r->1	
nd h	a->13	
nd i	 ->20	n->5	v->1	
nd j	u->1	
nd k	a->1	o->4	v->3	ä->1	
nd l	a->1	ä->2	
nd m	e->55	i->3	y->1	å->3	
nd n	y->1	ä->5	ö->1	
nd o	c->26	m->15	s->6	
nd p	a->1	å->5	
nd r	e->2	
nd s	e->6	i->1	j->1	k->4	m->1	o->25	t->5	y->1	ä->4	å->2	
nd t	.->1	a->1	i->11	v->1	
nd u	n->4	p->1	t->3	
nd v	a->4	e->2	i->4	ä->1	å->1	
nd ä	n->1	r->17	
nd å	t->1	
nd ö	v->1	
nd! 	L->1	N->1	
nd),	 ->1	
nd, 	5->1	D->1	E->1	F->1	I->2	N->1	S->2	b->1	d->4	f->3	h->2	k->2	l->1	m->5	n->1	o->7	p->1	r->2	s->6	t->1	u->2	v->2	
nd- 	(->1	
nd. 	V->1	
nd.A	n->1	t->1	
nd.D	e->8	i->2	
nd.E	m->1	
nd.F	r->1	
nd.G	e->1	
nd.H	e->1	
nd.I	 ->2	n->3	r->1	
nd.J	a->7	
nd.K	o->2	
nd.L	å->1	
nd.M	e->1	i->1	
nd.N	i->1	u->1	ä->1	
nd.O	m->2	
nd.P	å->1	
nd.S	o->1	
nd.U	p->1	
nd.V	a->1	i->2	
nd.Å	 ->1	
nd? 	H->1	
nd?.	 ->1	
nd?F	ö->1	
nd?J	a->1	
nda 	-->1	1->1	2->1	E->2	a->18	b->3	c->1	d->21	e->10	f->18	g->2	h->3	i->13	j->4	k->1	l->4	m->9	n->3	o->7	p->12	r->6	s->36	t->5	u->3	v->4	ä->4	ö->2	
nda,	 ->7	
nda.	B->1	D->3	F->2	H->1	I->1	K->1	M->1	N->2	R->1	V->2	
nda?	D->1	
ndab	o->2	
ndad	 ->6	e->11	
ndag	 ->1	e->2	s->2	
ndah	å->43	
ndai	r->1	
ndal	!->1	,->1	a->1	e->5	ö->1	
ndam	a->1	e->1	å->13	
ndan	 ->14	,->2	.->1	b->2	d->18	f->1	h->1	m->1	o->1	r->6	t->39	
ndar	 ->9	d->24	e->10	n->4	s->1	
ndas	 ->20	,->1	.->6	t->82	
ndat	 ->12	,->4	e->5	i->33	p->9	
ndba	r->9	
ndbe	t->1	
ndbu	l->1	
nde 	"->3	(->30	-->15	1->1	A->3	B->1	D->1	E->4	G->5	I->1	J->1	K->4	L->2	M->4	N->1	O->1	P->14	R->3	S->4	a->213	b->67	d->70	e->54	f->180	g->19	h->39	i->106	j->4	k->58	l->21	m->74	n->14	o->149	p->103	r->95	s->137	t->65	u->42	v->41	ä->33	å->40	ö->16	
nde!	 ->6	A->1	J->1	N->1	
nde"	,->1	
nde(	A->1	
nde,	 ->117	
nde.	 ->3	-->1	.->1	A->2	D->28	E->6	F->4	G->1	H->11	I->4	J->26	K->4	L->3	M->13	N->3	O->4	P->2	S->7	T->5	U->2	V->10	Å->1	
nde:	 ->37	
nde;	 ->4	
nde?	F->1	H->2	V->1	
ndeb	e->1	u->9	ä->1	
ndef	r->1	ö->12	
ndeh	ö->1	
ndek	o->9	r->1	
ndel	 ->12	,->4	.->3	a->9	e->1	n->3	s->60	
ndem	e->5	i->1	
nden	 ->231	"->1	,->43	.->38	:->3	;->1	?->1	N->1	a->40	b->2	s->24	
nder	 ->516	"->1	,->27	.->37	?->2	a->36	b->3	d->4	e->3	g->4	h->5	k->5	l->36	m->3	n->132	o->4	r->3	s->96	t->17	u->3	v->1	ä->3	ö->1	
ndes	 ->12	,->1	k->115	t->1	
ndet	 ->383	)->1	,->22	.->34	;->1	?->1	a->1	s->15	
ndev	a->6	i->2	
ndfu	l->1	
ndfä	l->4	
ndfö	r->4	
ndgä	n->2	
ndgå	r->2	t->1	
ndi 	r->1	s->1	
ndi:	 ->1	
ndic	a->1	
ndid	a->14	
ndie	,->1	n->5	r->1	
ndig	 ->25	,->2	.->3	a->39	h->210	t->120	
ndik	a->10	
ndin	a->1	
ndir	e->7	
ndis	 ->1	k->1	
ndit	 ->3	i->1	
ndiv	i->14	
ndku	r->1	
ndla	 ->21	.->2	d->10	r->118	s->14	t->7	
ndli	g->22	n->186	
ndlä	g->75	
ndlö	s->1	
ndme	d->3	
ndmä	n->1	
ndna	 ->4	
ndni	n->74	
ndo.	F->1	
ndom	 ->2	l->2	r->14	s->1	
ndon	 ->1	,->2	.->1	
ndor	s->1	
ndpe	l->1	
ndpr	i->1	
ndpu	n->103	
ndra	 ->357	,->22	.->7	:->4	;->2	b->5	d->21	g->3	h->1	k->1	n->4	r->33	s->23	t->24	
ndre	 ->52	.->1	?->1	n->3	s->2	
ndri	n->314	
ndro	m->1	
ndrä	n->2	
nds 	a->1	b->3	d->2	e->1	f->5	g->1	i->4	l->1	m->3	n->1	o->2	p->7	r->1	v->1	å->1	
nds,	 ->1	
ndsa	m->4	n->1	t->1	v->3	
ndsb	e->1	y->43	
ndsd	e->12	
ndsj	u->1	
ndsk	 ->5	-->1	a->30	o->5	t->1	
ndsl	ä->2	
ndsm	e->6	ä->3	
ndsp	l->3	o->2	r->3	
ndsr	e->5	ö->1	
ndss	y->1	
ndst	a->2	e->1	
ndsv	ä->1	
ndsä	n->1	
ndt 	f->1	h->1	o->1	s->1	t->1	u->1	
ndt,	 ->1	
ndte	s->1	
ndup	p->3	
ndus	t->114	
ndut	y->1	
ndva	g->1	l->24	t->1	
ndvi	k->39	n->2	
ndzi	o->4	
ndär	r->1	
ndå 	A->1	a->8	b->5	d->1	e->5	f->5	g->2	h->3	i->4	k->4	l->1	o->2	s->4	t->4	u->4	v->1	ä->2	
ndå,	 ->1	
ndå.	.->1	
ndée	,->1	
ndöv	t->1	
ne F	o->1	
ne a	n->2	t->3	v->1	
ne b	l->1	
ne d	e->1	i->1	
ne e	k->1	
ne f	o->1	r->2	å->1	ö->4	
ne g	ä->1	
ne h	a->5	j->1	ö->1	
ne i	 ->4	n->3	
ne j	a->1	e->1	
ne k	a->1	o->1	
ne l	o->1	
ne n	ä->4	å->1	ö->1	
ne o	c->6	m->2	
ne p	å->2	
ne q	u->2	
ne r	y->1	
ne s	o->5	å->1	
ne t	i->2	o->1	
ne v	a->1	i->1	
ne ä	r->2	
ne å	k->1	
ne! 	N->1	
ne, 	E->1	R->1	d->2	g->1	k->1	n->1	t->1	ä->1	
ne- 	o->1	
ne-A	l->1	r->1	
ne-M	a->1	
ne-s	t->1	
ne.D	e->3	
ne.J	a->1	
ne: 	N->1	
near	b->1	v->1	
neba	r->1	
nebo	e->1	
nebä	r->108	
nebö	r->7	
ned 	a->2	d->1	e->3	f->1	i->5	m->3	n->1	o->1	p->2	t->1	v->1	
ned.	E->1	J->1	
nede	r->9	
nedg	å->2	
nedl	a->1	ä->4	
nedm	o->3	
nedo	m->1	
nedr	a->2	u->1	
neds	k->4	t->3	
nedv	r->12	ä->1	
neex	e->1	
nefa	t->6	
neff	e->3	
nefi	t->5	
nega	t->26	
neha	r->2	v->1	
nehå	l->78	
nehö	l->4	
nej 	l->1	t->1	
nej,	 ->2	
nej.	(->1	
neka	 ->4	,->1	.->1	d->1	n->2	r->2	s->2	
nela	g->1	
nele	r->1	
neli	g->2	
nell	 ->50	,->3	.->2	a->198	t->28	
neln	,->1	.->1	
nels	e->1	
nelt	r->1	
nelu	x->1	
nema	n->4	
nen 	"->1	(->6	-->7	C->1	E->2	I->1	J->1	P->1	a->113	b->36	d->9	e->17	f->89	g->22	h->64	i->88	j->1	k->68	l->9	m->36	n->14	o->119	p->28	r->18	s->99	t->24	u->21	v->24	ä->43	å->3	ö->4	
nen!	N->1	
nen"	.->1	
nen)	N->1	
nen,	 ->113	
nen.	 ->4	(->1	)->6	.->7	1->1	A->2	B->2	D->37	E->7	F->6	G->1	H->11	I->4	J->16	K->2	L->2	M->6	N->6	O->4	P->7	R->2	S->3	T->1	U->2	V->16	Ä->2	
nen:	 ->1	
nen;	 ->3	
nen?	H->1	K->1	V->1	Ä->1	
nenJ	a->2	
nena	 ->2	
nene	r->8	
nens	 ->389	,->1	
nent	 ->7	,->1	.->1	a->4	e->4	i->1	
neon	a->1	l->1	
nepo	t->5	
ner 	(->3	-->6	E->1	I->4	J->1	K->2	[->1	a->19	b->12	d->24	e->28	f->30	g->8	h->10	i->46	j->5	k->10	l->2	m->46	n->5	o->67	p->7	r->2	s->80	t->34	u->5	v->13	ä->7	å->1	ö->1	
ner"	)->1	
ner,	 ->52	
ner-	p->10	
ner.	 ->2	(->1	-->1	.->1	A->1	B->1	D->13	F->1	G->1	H->2	I->6	J->11	K->2	L->1	M->2	N->1	R->1	S->1	T->1	U->1	V->5	Ä->2	
ner;	 ->1	
ner?	-->1	H->1	J->1	K->1	V->1	
nerN	ä->2	
nera	 ->16	d->25	l->20	n->7	r->10	s->10	t->11	
nere	 ->2	.->1	l->16	r->3	
nerg	i->111	
nerh	e->46	
neri	e->1	n->63	
nerl	i->14	
nern	a->208	
ners	 ->12	h->1	k->17	t->2	
nerö	s->4	
nes 	a->3	b->3	e->2	f->3	i->1	k->5	m->2	o->2	s->2	t->2	u->1	v->1	
nes,	 ->1	
nese	r->2	
nesi	s->8	
nesm	a->1	ä->1	
nesr	ö->1	
ness	 ->1	
nest	a->1	
net 	"->1	a->1	f->4	i->1	m->1	n->1	o->2	p->2	s->1	t->1	u->1	v->1	ä->1	
net,	 ->6	
net.	 ->1	D->4	F->1	I->1	J->1	M->1	N->1	O->1	V->1	
neta	r->1	
nete	c->6	
neti	s->1	
nett	 ->1	.->1	e->1	
netä	r->6	
neut	r->2	
nevå	n->2	
nez 	a->1	
nezu	e->1	
nfal	l->2	
nfat	t->12	
nfed	e->1	
nfek	t->2	
nfer	e->170	
nfes	s->1	
nfid	e->2	
nfil	t->1	
nfin	i->1	n->1	
nfis	k->2	
nfli	k->16	
nfly	k->1	t->12	
nfor	d->2	m->90	
nfra	s->15	
nfre	d->1	
nfri	a->1	
nfro	n->1	
nfrå	g->4	
nfär	d->1	
nför	 ->109	,->1	.->2	:->1	a->68	d->4	e->5	l->19	s->8	t->9	
ng (	1->1	E->1	a->2	r->1	å->1	
ng -	 ->11	,->1	
ng 1	7->1	9->1	
ng 2	0->2	
ng 3	7->1	
ng 6	0->1	8->1	
ng 8	0->2	
ng D	e->1	
ng E	c->1	u->1	
ng F	ä->1	
ng I	V->2	
ng T	a->1	
ng V	I->1	
ng a	j->1	l->4	n->8	r->1	t->27	v->329	
ng b	a->2	e->7	i->1	l->3	o->1	r->1	y->1	ö->5	
ng d	e->9	i->1	y->1	ä->7	
ng e	.->1	f->2	l->9	n->8	t->7	x->2	
ng f	i->5	o->1	r->29	u->1	å->2	ö->89	
ng g	a->1	e->8	j->1	l->1	r->1	å->1	
ng h	a->25	e->1	o->3	ä->1	å->1	
ng i	 ->90	a->1	n->32	r->1	
ng j	a->1	
ng k	a->7	n->1	o->19	r->2	u->1	
ng l	e->1	i->5	ä->2	å->1	
ng m	a->5	e->46	i->2	o->10	å->12	
ng n	e->1	i->4	r->2	u->1	ä->3	ö->1	
ng o	c->150	f->2	l->1	m->34	
ng p	e->2	l->1	o->1	r->4	å->53	
ng r	a->2	e->2	i->1	ä->3	ö->2	
ng s	a->3	e->2	i->11	k->21	o->108	t->6	y->1	ä->4	å->4	
ng t	a->7	i->74	r->3	y->2	
ng u	n->6	p->2	r->1	t->11	
ng v	a->9	e->3	i->16	o->1	ä->2	
ng ä	g->1	n->6	r->39	v->2	
ng å	t->5	
ng ö	k->1	v->2	
ng!J	a->1	
ng" 	a->1	o->1	
ng",	 ->2	
ng".	J->1	N->1	
ng) 	i->2	o->2	
ng).	V->1	
ng)N	ä->1	
ng, 	O->1	a->6	b->4	d->13	e->15	f->25	g->2	h->4	i->14	k->5	l->4	m->19	n->8	o->22	p->6	r->2	s->29	t->5	u->9	v->14	ä->4	å->3	ö->1	
ng-P	M->1	
ng. 	D->2	E->1	M->1	S->1	
ng.(	A->1	
ng..	 ->2	(->1	
ng.A	l->3	n->1	v->4	
ng.D	a->1	e->66	o->2	ä->6	
ng.E	f->1	n->5	t->1	u->1	
ng.F	l->1	r->5	ö->10	
ng.G	e->2	
ng.H	a->1	e->12	u->1	ä->1	ö->1	
ng.I	 ->13	n->2	
ng.J	a->32	
ng.K	a->1	o->8	
ng.L	i->1	å->2	
ng.M	a->6	e->4	y->1	å->2	
ng.N	a->1	i->3	u->2	ä->2	å->1	
ng.O	c->7	f->1	m->9	
ng.P	P->1	a->1	r->1	å->2	
ng.R	e->1	
ng.S	a->1	e->1	l->4	å->1	
ng.T	a->1	i->2	r->1	
ng.V	a->1	i->17	å->1	
ng.Ä	r->3	
ng: 	e->1	f->1	i->1	
ng:D	e->1	
ng; 	d->1	e->1	f->2	
ng?D	e->2	
ng?H	ä->1	
ng?J	a->1	
ng?O	l->1	
ng?T	y->1	
ng?Ä	r->1	
nga 	-->1	a->37	b->12	c->1	d->11	e->4	f->16	g->8	h->2	i->5	k->9	l->3	m->21	n->6	o->13	p->3	r->8	s->21	t->9	u->4	v->7	ä->7	å->10	ö->1	
nga,	 ->5	
nga.	J->2	V->1	
ngad	e->6	
ngag	e->18	
ngal	u->3	
ngan	d->13	
ngar	 ->330	!->1	"->1	)->1	,->52	-->1	.->83	:->7	;->1	?->1	e->9	i->15	n->159	s->3	
ngas	 ->12	.->2	t->2	
ngat	 ->3	s->1	
ngav	 ->1	
ngbr	o->1	
ngd 	a->1	b->2	f->5	i->1	n->1	o->4	s->2	y->1	ä->1	å->1	
ngda	 ->1	
ngde	 ->2	n->5	r->5	
ngdo	m->15	
ngdp	u->4	
ngdr	a->1	
ngdy	r->1	
nge 	E->1	a->4	b->1	d->4	e->1	h->2	i->2	k->2	m->1	n->2	o->5	p->4	s->12	t->1	u->1	v->5	ä->1	å->1	
nge,	 ->1	
ngef	ä->10	
ngel	 ->1	i->1	n->2	s->11	ä->23	
ngem	a->4	
ngen	 ->746	"->1	,->80	.->95	:->4	;->2	?->7	I->1	a->3	b->1	j->2	k->1	o->1	r->1	s->25	t->22	ä->1	
nger	 ->47	,->5	.->3	a->56	
nges	 ->6	,->2	.->1	f->1	
nget	 ->49	,->1	d->1	t->1	
ngfa	l->15	
ngfl	ö->1	
ngfo	n->1	r->20	
ngfr	i->1	u->1	
ngfu	n->1	
ngfä	r->2	
nggå	 ->1	s->1	
ngig	g->1	t->1	
ngil	t->1	
ngiv	a->5	e->1	i->6	n->1	
ngkö	r->1	
ngle	w->2	
ngli	g->37	
ngme	t->6	
ngmå	l->1	
ngna	 ->8	
ngni	n->44	
ngom	 ->3	.->1	
ngpo	l->2	
ngra	 ->2	n->2	
ngre	 ->56	,->1	.->6	d->2	m->1	p->11	s->2	
ngri	n->1	p->16	
ngro	d->1	
ngrä	n->1	
ngs 	b->1	d->1	e->1	h->1	k->1	p->1	s->3	v->1	
ngs-	 ->12	
ngsa	k->3	l->1	m->6	n->7	r->7	v->6	
ngsb	a->2	e->11	i->11	o->3	
ngsc	e->5	h->8	
ngsd	i->2	o->1	r->1	
ngse	n->1	r->1	t->1	
ngsf	a->7	e->2	i->31	l->1	o->22	r->15	u->11	ö->232	
ngsg	r->6	
ngsh	a->1	o->1	
ngsi	d->4	k->7	n->10	
ngsk	a->1	l->3	o->170	r->14	u->1	v->1	
ngsl	a->2	i->59	o->1	ä->6	ö->5	
ngsm	a->4	e->7	i->1	o->5	ä->2	å->4	ö->4	
ngsn	i->5	o->1	y->1	
ngso	m->10	r->2	
ngsp	a->4	e->3	l->23	o->21	r->46	u->11	å->1	
ngsr	e->18	i->15	u->1	ä->2	å->1	
ngss	a->2	e->4	i->2	k->14	p->1	t->19	y->24	ä->15	
ngst	 ->3	.->1	a->9	e->3	j->5	m->2	r->1	ä->1	
ngsu	m->1	t->6	
ngsv	e->4	i->33	ä->7	å->1	
ngsy	s->2	
ngsä	r->1	t->1	
ngså	r->1	t->5	
ngsö	v->1	
ngt 	a->1	b->3	d->5	f->3	h->2	i->7	k->2	m->5	n->2	s->7	u->2	v->1	ö->1	
ngt,	 ->1	
ngt.	D->1	M->1	V->1	
ngta	r->1	
ngte	r->8	
ngtg	å->11	
ngti	d->4	
ngto	n->5	
ngtv	ä->4	
ngue	r->2	
ngva	r->6	
ngäl	d->1	
ngå 	e->1	i->5	s->2	
ngå.	A->1	
ngåe	n->53	
ngån	g->1	
ngår	 ->14	.->2	
ngåt	t->6	
ngör	 ->1	i->2	
nham	n->1	
nhan	d->1	g->47	
nhas	 ->1	
nhed	r->2	
nhem	s->2	
nhet	 ->47	"->2	,->12	.->24	e->111	l->36	s->10	
nhil	l->1	
nho 	f->1	p->1	s->1	v->1	
nho.	 ->1	
nhos	 ->1	
nhun	d->1	
nhäl	l->32	
nhäm	t->6	
nhän	g->5	
nhål	l->55	
nhår	d->1	
nhöj	d->4	
ni 1	9->6	
ni 2	0->2	
ni a	l->4	n->1	r->1	t->18	v->1	
ni b	e->7	l->1	r->1	ä->1	
ni d	e->2	i->1	ä->1	å->3	
ni e	f->1	n->1	r->2	
ni f	i->1	r->3	å->1	ö->10	
ni g	e->2	ö->3	
ni h	a->19	e->1	ä->2	å->2	
ni i	 ->3	n->12	
ni j	u->3	
ni k	a->3	o->8	u->1	ä->5	
ni l	e->1	ä->1	ö->1	
ni m	e->2	å->1	
ni n	u->2	ä->6	
ni o	c->5	m->2	s->1	
ni p	a->1	e->1	å->1	
ni r	a->2	e->2	ä->1	
ni s	a->11	e->4	j->2	k->6	l->1	o->2	t->2	ä->5	
ni t	a->5	i->1	o->1	
ni u	n->1	p->3	t->1	
ni v	a->4	e->8	i->9	ä->2	å->1	
ni ä	r->6	v->1	
ni ö	n->1	
ni, 	b->1	d->1	f->4	h->4	i->1	m->1	o->3	t->1	
ni.(	P->1	
ni.A	l->1	
ni.D	ä->1	
nial	i->1	
nice	r->2	
nied	 ->1	.->1	
nief	u->1	
nien	 ->14	,->4	.->3	?->1	s->2	
nier	 ->15	,->2	.->1	a->12	i->1	n->5	s->2	
nies	k->2	
niet	 ->1	.->2	
nife	s->1	
nifr	å->2	
nig 	h->1	i->1	o->1	
niga	 ->2	,->1	.->2	
nigh	e->12	
nigt	 ->1	
nik 	D->1	s->5	u->1	
nik-	 ->1	
nika	 ->1	t->16	
nike	n->4	r->3	
nikt	 ->1	
nila	t->2	
nima	l->1	
nimb	u->1	
nime	r->1	
nimi	b->2	f->1	i->1	k->4	l->2	n->3	r->5	s->1	
nimo	r->1	
nimu	m->4	s->1	
nind	e->1	u->1	
nine	r->1	
ning	 ->841	"->2	)->2	,->125	.->157	:->4	;->2	?->4	a->308	d->1	e->580	f->1	o->4	p->2	r->1	s->410	t->4	
nins	p->1	
ninv	å->1	
nio 	V->1	b->2	f->1	l->1	m->7	p->1	t->1	
nio;	 ->1	
nion	 ->15	,->5	.->6	d->1	e->415	s->8	
nipa	.->1	
nipe	n->1	
nipp	a->3	
nire	f->1	
nisa	t->43	
nisc	h->1	
nise	r->57	
nisk	 ->25	a->38	o->91	t->8	
nism	 ->3	,->2	.->2	e->9	
nist	a->2	e->56	i->7	r->41	
nit 	d->1	e->2	f->2	v->1	
nit,	 ->1	
nit.	N->1	
nite	t->14	
niti	a->80	e->2	o->14	s->1	v->9	
nito	r->1	
nits	 ->7	,->1	
nitt	 ->7	,->1	e->5	l->1	s->1	
nitu	d->1	m->1	
nitz	 ->1	
nitä	r->1	
nium	 ->2	!->1	.->2	
nive	r->4	
nivå	 ->46	,->13	.->21	;->1	?->1	e->14	g->3	n->11	
nié 	u->1	
nj f	ö->2	
nj m	o->1	
nj.D	e->1	
nje 	(->1	m->5	o->1	s->4	
nje.	G->1	J->1	
njen	 ->3	.->1	
njer	 ->36	"->1	,->6	.->3	:->1	n->31	
njor	 ->1	
njun	k->1	
njut	e->1	n->1	
njuv	e->1	
njäm	k->1	
njär	e->1	
njör	 ->2	
nk b	a->1	
nk e	n->1	
nk h	o->1	
nk p	å->1	
nk r	a->1	
nk t	i->1	
nk u	t->1	
nk v	ä->1	
nk" 	f->1	
nk- 	e->1	
nk.D	e->1	
nka 	a->4	b->1	d->2	e->2	h->2	m->2	n->1	o->2	p->16	s->7	v->1	ö->2	
nka,	 ->1	
nka.	E->1	Å->1	
nkal	l->9	
nkan	d->288	
nkar	 ->10	,->1	.->4	a->1	n->2	
nkas	 ->2	,->1	
nkat	a->1	
nkba	r->4	
nke 	a->1	l->1	o->1	p->40	r->1	t->2	ä->2	
nke,	 ->2	
nkeb	a->1	
nkef	r->1	
nkeg	å->1	
nkel	 ->9	.->3	:->2	m->1	n->2	r->1	t->28	v->2	
nken	 ->20	,->2	.->1	:->1	s->1	
nkep	o->1	
nker	 ->45	,->2	n->3	s->1	ä->1	
nkes	i->1	
nkfa	r->7	
nkfo	r->1	
nkfö	r->1	
nkir	e->1	
nkit	 ->2	
nkla	 ->10	d->1	g->4	r->5	s->3	t->1	
nkli	g->5	n->1	
nklu	d->4	s->17	
nkna	 ->1	d->1	r->1	t->1	
nkni	n->15	
nkny	t->1	
nko.	T->1	
nkol	e->1	
nkom	l->3	m->1	p->3	s->12	
nkon	s->1	t->2	v->3	
nkop	p->1	
nkra	 ->1	d->3	f->22	r->5	
nkre	n->2	t->58	
nkri	k->39	s->1	
nkrä	k->1	
nks 	o->2	t->1	
nksa	m->2	
nksc	h->1	
nkse	k->1	
nkt 	(->2	-->2	1->3	2->3	4->2	5->1	6->1	7->1	D->1	a->6	b->1	d->4	e->2	f->6	g->4	h->5	i->16	k->2	m->4	n->2	o->6	p->29	r->1	s->21	t->2	u->1	v->3	ä->8	
nkt,	 ->14	
nkt.	 ->1	A->1	D->5	I->1	M->3	N->2	P->1	T->2	V->4	
nkt:	 ->2	
nkt?	E->1	
nkta	 ->6	,->1	.->1	
nkte	 ->3	n->88	r->86	
nkti	o->41	v->1	
nkts	 ->4	p->1	
nktu	r->1	
nkur	r->285	
nkän	n->1	
nköp	 ->1	s->1	
nkör	s->1	
nlag	t->1	
nlam	p->1	
nlan	d->7	
nlar	 ->1	n->1	
nled	a->31	d->10	e->8	n->57	s->5	
nlet	t->13	
nlig	 ->14	,->1	.->1	a->36	e->17	g->1	h->37	t->139	
nlit	a->1	
nlys	n->1	
nläg	g->32	
nläm	n->5	
nlän	d->6	k->1	t->1	
nlås	t->1	
nlåt	a->1	
nlöp	a->2	e->3	
nlös	 ->1	
nman	ö->1	
nmar	k->26	
nmäl	a->3	d->1	e->1	n->12	s->2	t->1	
nmär	k->12	
nmäs	s->2	
nmöt	e->2	
nn d	e->1	
nn e	u->1	
nn o	c->1	
nn t	i->1	
nn ä	r->1	
nn, 	d->1	e->1	
nn-g	r->1	
nna 	-->2	E->1	T->2	a->34	b->45	c->2	d->49	e->21	f->131	g->49	h->16	i->26	j->1	k->66	l->23	m->37	n->6	o->37	p->53	r->74	s->98	t->42	u->36	v->44	y->2	ä->6	å->15	ö->8	
nna,	 ->4	
nna.	 ->2	-->1	D->1	J->3	O->1	U->1	V->2	Ä->1	
nna?	S->1	
nnab	i->1	
nnad	e->6	
nnag	a->3	e->3	i->3	
nnak	i->2	
nnal	a->1	
nnam	b->1	
nnan	 ->76	,->4	.->1	d->28	s->2	
nnar	 ->11	e->1	s->19	
nnas	 ->52	!->1	,->2	.->3	
nnat	 ->111	,->1	.->4	
nndr	a->1	
nne 	F->1	a->4	f->4	h->4	n->1	o->1	p->2	s->1	t->1	ä->2	å->1	
nne!	 ->1	
nne,	 ->5	
nne.	D->1	J->1	
nneb	a->1	o->1	ä->108	ö->7	
nned	o->1	
nnef	a->6	
nneh	a->3	å->78	ö->4	
nnel	a->1	i->1	n->2	t->1	
nnen	 ->39	,->2	.->5	a->1	s->11	
nner	 ->129	,->5	.->5	h->46	l->12	s->2	
nnes	 ->24	,->1	m->2	r->1	
nnet	 ->1	.->2	e->6	
nnev	å->2	
nnhe	t->1	
nnie	f->1	n->14	r->5	s->2	t->3	
nnig	 ->2	a->1	h->3	t->1	
nnin	g->79	
nnis	k->98	
nnit	 ->6	,->1	.->1	s->8	
nniu	m->3	
nniv	å->1	
nnla	n->1	r->2	
nnli	g->2	
nnly	s->1	
nnlä	n->1	
nnoc	k->24	
nnol	i->9	
nnop	r->2	
nnor	 ->37	,->3	.->4	?->1	l->2	n->5	s->12	
nnov	a->6	
nns 	2->1	G->1	S->1	a->17	b->5	c->1	d->59	e->53	f->25	g->4	h->5	i->43	j->2	k->3	l->1	m->23	n->20	o->12	p->8	r->10	s->15	t->15	u->1	v->5	y->2	ä->3	å->1	ö->2	
nns,	 ->3	
nns.	D->3	E->1	J->1	M->1	V->1	
nnsa	k->1	m->3	
nnsk	a->1	
nnu 	a->1	e->12	f->1	h->6	i->32	m->8	n->1	p->1	s->10	v->2	ä->1	
nnu.	D->1	K->2	V->1	
nnu;	 ->1	
nnyt	t->2	
nnäe	r->1	
nnäm	n->2	
no L	e->1	
no P	r->2	
no i	 ->1	
no k	o->1	
no o	c->1	m->1	
no u	n->1	
no, 	T->1	m->1	
no.J	a->1	
no.O	r->1	
nock	 ->12	,->6	.->3	s->3	
nodl	a->2	i->1	
nog 	a->3	b->1	d->2	h->2	i->1	k->1	n->1	o->1	p->1	ö->1	
nog,	 ->1	
nog.	M->2	
noga	 ->9	,->1	.->2	
nogg	r->12	
nogr	a->2	
nois	e->1	
noku	l->3	
noli	k->9	
noll	,->1	n->1	r->1	
nolo	g->3	
nom 	-->1	2->1	5->1	A->1	D->1	E->39	F->1	G->1	I->1	L->1	S->2	V->1	W->1	a->115	b->8	d->70	e->38	f->14	g->9	h->7	i->10	j->4	k->26	l->5	m->14	n->5	o->14	p->8	r->59	s->21	t->13	u->22	v->17	y->1	ä->2	å->4	ö->7	
nom,	 ->3	
nom.	 ->1	H->2	J->1	M->1	V->1	
noma	r->2	
nomb	l->5	r->2	
nomd	r->6	
nome	n->6	r->1	u->1	
nomf	ö->161	
nomg	i->1	r->4	å->11	
nomi	 ->20	,->2	.->3	?->1	e->8	n->33	s->219	
noml	ä->2	
nomr	å->1	
noms	k->1	l->3	n->11	y->3	
nomt	ä->1	
non 	e->1	f->2	o->1	
non,	 ->1	
non.	E->1	
non?	K->1	
none	r->1	
nony	m->5	
nopo	l->17	
nopr	o->2	
nor 	a->1	e->1	f->1	i->10	o->14	s->9	t->1	
nor,	 ->3	
nor.	D->2	F->3	J->2	V->1	
nor?	H->1	
nord	a->4	e->1	i->3	k->1	l->4	n->9	t->1	v->1	
nore	r->4	
nori	t->22	
norl	u->2	
norm	 ->7	a->31	e->32	t->7	
norn	a->6	
norr	?->1	a->4	
nors	 ->10	t->2	
nos 	h->1	i->1	o->1	t->1	
nos!	 ->1	
nos,	 ->2	
nota	n->1	
note	r->28	
noti	s->1	
nott	i->1	
nova	t->6	
nove	m->11	r->3	
now-	h->1	
npas	s->14	
npor	n->2	
npri	n->2	
npro	b->1	
nprä	n->1	
npun	k->31	
npå 	d->1	
nr 1	 ->1	2->2	7->2	
nr 2	8->1	9->1	
nr 3	0->1	1->1	2->1	3->2	5->1	6->1	7->1	8->1	9->1	
nr 4	0->1	1->1	2->1	3->1	4->1	5->1	6->1	
nr 5	 ->1	
nr 6	 ->1	
nr 7	.->1	
nr 8	 ->1	
nr 9	 ->1	
nra 	k->1	o->10	
nrad	 ->1	
nrar	 ->1	
nras	 ->1	
nre 	a->2	e->2	g->1	m->69	v->9	
nreg	e->1	
nren	i->1	
nres	a->5	u->1	
nrik	e->13	t->44	
nry 	F->1	
nrym	s->1	
nrät	t->56	
nråd	e->1	
nröj	a->5	t->1	
nröt	t->1	
ns -	 ->1	
ns 2	4->1	8->1	
ns B	N->3	
ns E	U->1	u->2	
ns G	e->1	
ns H	e->1	
ns I	s->1	
ns S	O->1	
ns V	D->1	
ns X	X->1	
ns a	b->2	d->1	g->2	k->1	l->11	m->1	n->25	r->17	t->11	u->1	v->12	
ns b	a->2	e->47	i->2	l->3	r->1	u->7	y->1	ä->1	å->2	
ns c	e->1	i->1	
ns d	a->12	e->66	i->5	o->6	ä->7	ö->1	
ns e	f->6	g->6	k->18	l->1	m->2	n->38	t->18	u->1	x->4	
ns f	a->9	e->2	i->4	l->5	o->11	r->21	u->3	y->1	å->1	ö->78	
ns g	a->2	e->13	o->3	r->10	ä->1	å->1	
ns h	a->7	e->1	i->5	o->2	u->2	ä->8	å->1	
ns i	 ->29	d->1	k->1	m->1	n->71	
ns j	o->2	u->5	
ns k	a->2	o->31	r->4	u->5	v->6	ä->2	
ns l	a->13	e->2	i->4	j->1	o->2	u->1	ä->9	ö->1	
ns m	a->6	e->67	i->6	o->5	y->4	ä->1	å->17	ö->5	
ns n	a->6	e->1	i->3	u->8	y->1	ä->2	å->16	ö->1	
ns o	b->3	c->36	d->1	i->2	l->2	m->34	r->15	s->1	t->3	
ns p	a->11	e->2	l->2	o->13	r->13	å->10	
ns r	a->16	e->41	i->8	o->8	u->1	ä->18	å->1	ö->1	
ns s	a->16	c->1	e->5	i->20	j->1	k->14	l->7	m->1	n->3	o->17	p->4	t->38	v->3	y->3	ä->9	å->4	
ns t	a->4	e->9	i->15	j->7	o->1	r->6	u->1	v->6	
ns u	n->1	p->8	r->5	t->46	
ns v	a->5	e->10	i->23	o->1	ä->13	
ns y	t->9	
ns ä	g->4	n->4	r->7	v->1	
ns å	l->2	r->3	s->3	t->5	
ns ö	d->3	k->2	r->1	v->9	
ns!V	i->1	
ns, 	b->2	d->6	e->1	f->4	j->1	m->5	n->3	o->11	p->1	s->4	t->1	v->2	ä->2	
ns- 	o->6	
ns.D	e->10	ä->2	
ns.E	n->1	u->1	
ns.F	ö->1	
ns.I	 ->1	
ns.J	a->3	
ns.L	å->1	
ns.M	a->1	e->1	y->1	
ns.O	a->1	
ns.S	o->1	
ns.V	a->1	
ns/d	e->1	
ns: 	h->1	
ns; 	v->1	
ns?.	H->1	
ns?E	t->1	
ns?J	a->1	
nsa 	a->2	d->2	m->1	p->1	s->3	t->2	u->3	
nsa,	 ->1	
nsad	 ->13	,->1	.->3	e->10	
nsaf	f->2	
nsak	a->1	
nsam	 ->50	,->1	l->8	m->135	r->1	t->28	
nsan	a->1	d->3	
nsar	 ->6	b->8	
nsas	 ->5	
nsat	 ->7	.->3	i->3	s->49	t->4	
nsav	g->1	t->1	
nsbe	g->3	r->1	s->6	v->2	
nsbo	l->1	
nsbr	i->1	
nsbu	t->1	
nsch	 ->3	.->1	?->1	e->4	
nsda	g->5	
nsde	b->2	p->1	
nsdi	r->1	
nsdo	k->1	m->1	
nsdu	g->2	
nsdö	m->1	
nse 	a->8	d->2	h->1	m->4	o->1	v->4	
nse,	 ->1	
nse.	E->1	
nse;	 ->1	
nsee	n->11	
nsek	v->61	
nsem	e->3	
nsen	 ->124	,->13	.->39	?->1	N->1	l->1	s->18	
nser	 ->263	,->6	.->10	?->3	a->15	i->1	n->36	v->7	
nses	 ->5	
nset	t->2	
nseu	r->1	
nsfo	r->1	
nsfr	i->3	ä->1	å->5	
nsfu	n->1	
nsfö	r->22	
nsgr	u->1	
nsha	u->1	
nshi	n->10	
nshä	m->2	
nsib	i->1	
nsid	i->4	
nsie	l->28	r->50	
nsif	i->3	
nsik	t->5	
nsin	 ->11	.->1	d->1	i->1	n->2	r->1	s->1	
nsio	n->27	
nsis	k->2	t->6	
nsit	e->1	i->2	l->3	r->1	t->1	
nsiv	 ->3	a->3	t->6	
nsiä	r->1	
nsjo	v->17	
nsk 	T->1	b->1	d->1	k->1	l->2	n->1	p->2	r->1	s->1	
nska	 ->178	,->3	.->6	d->13	f->1	m->1	n->16	p->317	r->32	s->6	t->15	
nske	 ->66	,->1	m->3	
nski	l->28	
nskl	i->43	
nskn	i->41	
nsko	m->19	n->18	s->2	
nskr	a->36	i->5	ä->12	
nskt	 ->6	.->1	a->1	
nsku	l->6	r->6	
nskv	ä->10	
nsla	 ->13	"->1	,->1	g->30	
nsle	d->11	n->2	r->1	s->5	
nsli	e->1	g->21	
nslo	g->1	l->1	m->1	r->5	
nslu	t->29	
nslä	g->1	
nslå	 ->1	d->1	r->1	s->2	
nsme	d->5	
nsmi	n->2	
nsmo	m->1	
nsmy	n->8	
nsmä	l->1	n->5	s->1	
nsmå	l->1	
nsmö	t->1	
nsna	c->2	
nsni	n->19	v->2	
nsol	i->3	
nsom	r->3	
nsor	d->2	
nspa	k->1	r->1	
nspe	k->12	l->1	
nspi	r->3	
nspl	a->2	
nspo	l->79	r->108	
nspr	i->6	o->6	å->7	
nsra	d->1	m->1	
nsre	g->12	l->1	
nsro	l->1	
nsrä	t->43	
nssa	m->7	
nssc	h->1	
nsse	k->1	
nssi	t->1	
nssk	a->2	y->2	
nsst	r->2	ä->20	ö->1	
nssv	å->1	
nssy	s->6	
nst 	-->1	1->2	3->2	4->1	a->1	b->1	d->2	f->1	i->3	l->1	m->2	n->1	o->4	p->2	r->1	s->5	u->2	v->2	å->1	
nst,	 ->3	
nst.	J->2	
nsta	 ->5	b->1	g->2	k->5	l->2	n->37	t->46	
nste	e->5	f->6	k->2	l->1	m->39	n->5	p->1	r->77	s->2	
nstf	u->1	
nstg	ö->3	
nsti	g->3	l->3	n->3	t->158	
nstj	ä->1	
nstm	a->1	
nsto	n->27	r->2	
nstr	a->4	e->14	u->89	ä->46	å->1	
nsts	v->1	
nstä	l->58	m->23	n->5	
nstå	e->1	
nsul	t->5	
nsum	e->61	t->2	
nsun	d->3	
nsup	p->1	
nsut	b->3	s->2	
nsva	r->311	
nsve	r->1	
nsvi	l->10	
nsvä	n->1	r->12	
nsyn	 ->74	,->1	.->3	;->1	e->4	s->2	
nsäg	a->1	
nsäk	e->3	
nsäm	n->1	
nsär	e->2	
nsät	t->9	
nsåg	 ->12	
nsåt	e->1	g->1	
nsök	a->8	n->1	t->1	
nsöv	e->12	n->1	
nt (	t->1	
nt -	 ->7	
nt 1	9->2	
nt A	s->1	
nt C	l->1	
nt E	u->2	
nt a	l->5	n->5	r->1	t->16	v->54	
nt b	a->2	e->2	i->1	o->1	r->1	u->1	ö->2	
nt c	e->1	
nt d	e->6	i->1	
nt e	k->1	l->3	n->3	t->1	x->3	
nt f	a->5	i->1	r->5	u->1	y->1	ö->44	
nt g	a->1	e->4	r->1	ä->2	
nt h	a->9	e->1	o->1	u->2	å->1	
nt i	 ->17	d->1	f->1	g->1	n->13	
nt k	a->5	o->8	r->2	u->1	v->1	ä->1	
nt l	e->1	i->1	j->1	ö->1	
nt m	a->1	e->8	i->1	o->2	å->3	ö->1	
nt n	u->1	y->1	ä->1	å->2	
nt o	c->27	m->11	
nt p	l->1	r->4	u->1	å->5	
nt r	e->2	
nt s	a->2	e->6	i->2	j->2	k->4	l->1	n->1	o->37	t->5	v->1	y->2	ä->12	å->2	
nt t	a->2	e->3	i->16	v->1	
nt u	n->6	p->2	r->1	t->5	
nt v	a->2	e->1	ä->1	å->1	
nt ä	m->1	n->1	r->5	
nt å	t->1	
nt ö	n->1	v->3	
nt!"	J->1	
nt, 	L->1	S->1	a->2	b->1	d->5	e->2	f->3	g->1	h->2	i->6	k->1	l->1	m->3	o->5	r->2	s->2	u->2	v->1	
nt-E	x->1	
nt. 	V->1	
nt.D	e->13	
nt.E	n->1	u->1	
nt.F	r->1	ö->3	
nt.H	e->3	
nt.I	 ->4	
nt.J	a->6	
nt.L	å->1	
nt.M	a->1	e->2	
nt.N	ä->1	
nt.O	K->1	
nt.P	l->1	
nt.S	a->2	å->2	
nt.V	i->3	
nt: 	U->1	v->1	
nta 	-->1	1->1	M->1	N->1	S->2	a->4	b->6	d->5	e->12	f->25	h->1	i->4	k->4	l->1	m->6	n->11	o->2	p->5	r->2	s->20	t->4	u->1	ä->2	å->1	
nta,	 ->1	
nta.	 ->1	D->1	
ntab	l->1	r->3	
ntad	e->1	
ntag	 ->12	,->4	.->2	?->1	a->17	e->6	i->22	l->1	n->4	s->10	
ntai	n->1	
ntak	t->17	
ntal	 ->41	,->1	a->4	e->19	i->1	s->11	
ntam	i->2	
ntan	 ->4	.->1	?->1	a->1	d->2	s->6	t->13	
ntar	 ->55	,->1	.->1	e->21	i->31	
ntas	 ->13	,->2	.->1	i->2	t->9	
ntat	 ->8	.->1	e->1	i->18	
ntav	 ->1	
nte 	-->3	1->1	B->1	E->3	a->138	b->141	c->1	d->56	e->59	f->123	g->74	h->166	i->47	j->1	k->102	l->65	m->62	n->49	o->32	p->46	r->35	s->104	t->72	u->50	v->50	ä->85	å->6	ö->12	
nte!	D->1	M->1	
nte,	 ->15	
nte.	A->1	B->1	D->3	H->2	J->2	S->1	V->2	Å->2	
nte:	 ->1	
nte?	F->1	H->1	
nteg	r->42	
ntek	n->3	
ntel	l->9	s->5	
ntem	o->27	
nten	 ->30	"->1	)->1	,->6	.->6	?->1	s->16	t->1	
nter	 ->23	,->2	-->1	.->7	a->128	i->48	n->138	p->1	v->10	
ntes	.->1	
ntet	 ->308	,->37	-->1	.->29	:->1	?->1	s->103	
ntex	t->1	
ntfr	å->6	
nti 	-->1	f->5	h->2	i->4	k->1	o->3	p->1	s->1	v->1	
nti!	 ->3	
nti,	 ->3	
nti-	g->1	i->1	r->1	
nti.	H->1	J->1	V->1	
ntia	l->3	
ntib	e->1	
ntid	e->1	
ntie	l->8	r->20	u->1	
ntif	a->3	i->15	o->3	
ntik	a->1	o->1	r->2	
ntil	 ->1	e->1	i->1	
ntim	e->1	t->1	ö->1	
ntin	 ->3	e->5	g->72	s->1	u->2	
ntio	n->41	
ntiq	u->1	
ntis	e->5	k->6	y->1	
ntit	a->4	e->8	r->1	
ntka	t->1	
ntku	s->1	
ntli	g->249	
ntni	n->8	
ntog	 ->16	s->10	
ntol	e->4	
ntom	 ->1	
nton	s->1	
ntor	 ->5	,->2	e->2	g->1	
ntpo	l->2	
ntpr	a->1	
ntra	 ->12	,->1	d->1	k->4	l->76	n->3	p->1	r->8	s->5	t->17	
ntre	a->2	l->1	p->5	r->15	s->120	t->1	
ntro	d->6	l->180	v->4	
ntru	m->9	
ntry	c->15	
nträ	d->36	f->26	t->1	
ntrå	n->1	
nts 	a->6	b->1	e->1	f->1	h->1	i->3	m->3	o->1	p->1	t->1	v->1	ä->1	
nts,	 ->2	
nts.	D->1	J->1	
ntsa	t->1	
ntsb	e->1	
ntsf	o->1	
ntsi	f->1	
ntsk	a->1	o->1	y->5	
ntsl	e->28	
ntsu	t->2	
ntti	l->1	
ntue	l->21	
ntun	n->1	
ntur	e->1	
ntus	i->3	
ntva	r->1	
ntve	r->2	
ntvä	n->1	
ntyd	d->2	i->4	
ntyg	 ->1	a->3	
ntyr	a->9	
ntäk	t->5	
ntär	a->2	
ntón	i->1	
ntör	e->2	s->1	
nu -	 ->1	
nu 3	4->1	
nu E	r->1	
nu a	l->1	n->1	t->5	v->1	
nu b	e->4	l->4	
nu d	e->4	i->2	ö->1	
nu e	f->1	g->1	n->12	t->8	u->1	
nu f	a->2	i->3	l->1	r->2	å->3	ö->10	
nu g	e->5	ä->3	å->3	ö->3	
nu h	a->13	å->3	ö->5	
nu i	 ->3	g->1	n->38	
nu k	a->5	o->6	
nu l	i->1	y->1	ä->3	
nu m	e->8	i->1	ä->1	å->8	
nu n	u->1	ä->8	å->1	
nu o	c->4	f->2	m->1	
nu p	l->1	r->2	å->4	
nu r	u->1	å->2	ö->1	
nu s	e->2	i->1	k->7	l->1	m->1	o->1	p->1	t->11	v->1	ä->2	å->2	
nu t	a->5	i->3	y->3	
nu u	n->1	p->3	
nu v	a->1	e->2	i->6	
nu ä	l->1	n->6	r->10	
nu å	t->1	
nu, 	e->1	i->1	m->2	u->1	ö->1	
nu..	T->1	
nu.D	e->1	
nu.J	a->1	
nu.K	o->2	
nu.L	å->1	
nu.V	i->2	
nu: 	g->1	
nu; 	i->1	
nu?J	a->1	
nuar	i->16	
nuc 	s->1	
nuer	l->2	
nuft	 ->1	.->1	e->1	i->11	
null	i->1	
nulä	g->1	
num 	f->1	h->1	i->1	ä->1	
num.	D->1	
nume	r->5	
numm	e->2	
nunn	o->1	
nupp	r->4	
nus 	2->1	f->1	t->1	
nusd	i->1	
nusg	r->2	
nuss	l->1	
nut 	f->2	n->1	
nut.	(->1	)->1	J->1	
nute	n->3	r->10	t->1	
nutn	a->2	
nutp	u->1	
nuts	-->1	
nutt	a->2	
nutv	e->1	
nuva	r->45	
nval	d->1	
nvan	d->18	
nvap	e->12	
nvar	a->4	o->4	
nvec	k->2	
nven	t->25	
nver	g->5	k->7	s->1	
nves	t->15	
nvet	e->1	
nvik	t->5	
nvin	k->12	
nvis	a->27	h->3	n->10	t->1	
nvit	 ->1	
nvol	v->9	
nväg	 ->8	,->1	.->2	a->9	s->3	
nvän	d->187	t->12	
nvär	d->1	
nvån	a->9	
ny b	i->1	
ny e	u->1	
ny f	a->1	o->1	ö->2	
ny g	r->1	
ny h	ä->1	
ny i	n->2	
ny k	e->1	o->3	u->3	v->1	
ny l	a->1	e->1	i->1	
ny m	y->1	
ny o	c->1	l->1	
ny p	e->2	
ny r	ö->2	
ny s	e->1	i->1	p->1	t->1	y->2	
ny t	y->1	
ny u	p->1	
ny v	e->1	i->2	
nya 	"->1	8->1	E->3	a->12	b->14	d->5	e->2	f->10	g->3	i->4	j->1	k->17	l->7	m->17	n->2	o->6	p->13	r->16	s->7	t->8	u->3	v->4	ä->2	å->6	
nya,	 ->1	
nya;	 ->1	
nyan	d->1	s->3	
nyar	 ->1	
nyas	 ->1	t->1	
nyba	r->39	
nybi	l->2	
nyck	e->8	
nyda	n->1	
nye 	o->1	
nyel	s->6	
nyet	a->1	
nyfa	s->1	
nyfö	r->1	
nyhe	t->13	
nykt	e->2	r->1	
nyli	b->1	g->29	
nym 	m->1	s->1	
nym.	D->1	
nyma	 ->1	
nymi	t->1	
nyna	z->6	
nyo 	s->1	
nyon	 ->2	,->1	
nypl	a->1	
nysk	a->1	
nyss	 ->10	,->2	.->1	
nyta	 ->5	
nyte	r->2	
nytn	i->1	
nyts	 ->1	
nytt	 ->40	,->3	.->3	a->20	i->13	j->41	o->2	
nyva	l->1	
nyår	s->1	
nz F	i->3	l->2	
nz b	e->1	
nz e	t->1	
nz f	r->1	ö->1	
nz o	c->6	m->1	
nz t	o->1	
nz)(	T->1	
nz).	H->1	
nz, 	L->3	
nzFr	u->1	
nzbe	t->1	
nzes	-->1	
nzál	e->1	
nÄra	d->1	
näck	a->2	
näer	;->1	
nägn	a->1	
näll	a->1	e->1	
näml	i->43	
nämn	a->30	d->26	e->5	i->3	s->9	t->19	v->1	
nämt	 ->1	
när 	-->2	A->1	B->9	C->1	E->1	K->5	M->14	N->1	P->18	R->2	S->2	V->4	W->1	a->9	b->3	c->1	d->199	e->8	f->7	g->2	h->13	i->1	j->14	k->7	l->1	m->23	n->10	o->1	p->1	r->3	s->3	t->1	v->43	ä->2	ö->2	
när!	 ->29	.->1	E->1	J->1	
när,	 ->75	
när.	 ->1	D->2	G->1	J->6	V->1	
nära	 ->27	,->1	
näre	n->46	r->20	
närf	r->1	
närh	e->5	
näri	n->12	
närm	a->36	e->1	n->5	
närp	e->1	
närs	 ->1	y->1	
närv	a->46	
näsd	u->1	
näst	a->47	
nät 	k->1	o->2	s->2	
nät.	 ->1	
näte	n->2	t->2	
näts	t->1	
nätt	e->1	
nätv	e->11	
näva	r->1	
nå a	n->1	
nå d	a->1	e->12	
nå e	k->2	n->20	t->6	
nå f	a->1	r->5	
nå g	e->1	
nå h	ö->1	
nå m	e->2	å->1	
nå n	å->1	
nå p	å->2	
nå r	e->1	
nå s	i->1	
nå v	å->5	
nå y	t->1	
nå ä	n->1	
nå å	t->1	
nå ö	n->1	
nå, 	n->1	
nå. 	D->1	
nå.F	r->1	
nå.J	a->1	
nå.S	l->1	
nåba	r->2	
nåd 	a->1	
nåda	 ->1	
nådd	a->3	e->3	
någo	n->165	r->1	t->192	
någr	a->147	
nåla	 ->2	,->1	r->2	
når 	d->5	e->5	m->3	s->1	v->1	
nåri	g->1	n->1	
nås 	b->1	e->1	g->1	i->2	
nås.	F->1	L->1	
nått	 ->13	,->1	.->1	s->5	
nçoi	s->1	
nève	 ->1	,->1	k->1	
nödb	e->1	
nöde	n->1	
nödi	g->12	n->1	
nöds	i->1	
nödv	ä->124	
nöja	 ->8	k->2	
nöjd	 ->2	a->9	
nöje	 ->4	r->1	t->2	
nöjt	 ->1	
nör 	t->1	
nör,	 ->1	
nörs	k->2	
nöst	e->19	
nöt.	D->1	
nötk	ö->3	
nöts	k->1	
nött	e->1	
növa	d->1	
növi	t->1	
növr	a->1	
o (K	O->2	
o - 	d->1	e->1	t->1	
o 19	9->1	
o Ca	d->5	
o Eu	r->1	
o Le	o->1	
o Pr	o->2	
o Ro	j->1	
o Sá	n->1	
o To	m->2	
o Tr	a->1	
o Va	l->3	
o Vi	t->1	
o ac	c->1	
o an	g->1	
o at	t->8	
o be	a->1	s->2	
o bl	a->1	
o bä	r->1	
o de	t->1	
o di	s->1	
o då	,->1	
o et	t->1	
o fa	r->1	t->1	
o fr	a->1	å->1	
o fu	l->1	
o fö	r->19	
o go	d->1	
o gr	a->2	
o gå	n->3	
o ha	r->4	
o hå	r->1	
o i 	a->1	d->1	e->2	f->3	h->1	l->1	m->1	n->1	
o in	t->1	
o ka	n->2	
o ko	m->1	
o kv	a->1	
o kä	m->1	
o le	d->1	
o lä	n->1	
o me	d->1	l->1	
o mi	l->6	n->1	
o må	l->1	n->2	s->1	
o nä	r->2	
o nå	g->3	
o oc	h->16	k->2	
o om	 ->3	
o pe	r->2	
o pu	n->1	
o på	 ->4	p->1	
o re	s->1	
o sa	d->1	f->1	
o si	n->1	
o sk	i->1	u->1	
o so	m->15	
o så	 ->2	
o ti	l->5	m->1	
o tr	e->1	
o un	d->2	
o ut	a->1	t->1	
o va	r->2	
o vi	k->1	l->1	
o vä	l->1	
o än	d->1	
o är	 ->7	
o äv	e->2	
o år	 ->4	,->1	e->2	s->1	
o åt	e->1	
o öp	p->1	
o öv	e->1	
o!Al	l->1	
o, A	s->1	
o, H	e->1	
o, T	a->1	
o, W	y->1	
o, a	n->1	t->1	
o, d	e->4	ä->1	
o, e	l->1	t->2	
o, f	ö->2	
o, h	e->1	u->1	
o, i	 ->2	
o, k	o->1	
o, m	e->2	o->1	
o, o	c->5	r->1	
o, s	a->1	e->1	o->6	t->1	y->1	
o, t	i->2	
o, v	i->2	
o, ä	n->1	
o- o	c->1	
o-Pl	a->4	
o-af	f->1	
o-an	a->1	
o-pr	o->1	
o-rå	d->1	
o. D	e->1	
o.- 	(->1	
o.At	t->1	
o.Av	s->1	
o.Be	t->1	
o.De	s->1	t->4	
o.Dä	r->1	
o.Eu	r->1	
o.Fl	e->1	
o.Fö	r->3	
o.He	r->2	
o.Hu	r->1	
o.Ja	g->5	
o.Kn	a->1	
o.Ko	m->1	
o.Lå	t->1	
o.Me	n->1	
o.Nä	r->2	
o.Oc	h->1	
o.Om	 ->2	
o.Or	d->1	
o.Se	d->1	
o.Tr	o->1	
o.Ty	 ->1	
o.Vi	 ->5	
o.m.	 ->6	,->1	
o/Oi	l->1	
o: v	i->1	
o; d	e->1	
o? D	e->1	
o?Hu	r->1	
oNäs	t->1	
oU, 	n->1	
oU-r	a->1	
oa f	ö->1	
oa o	s->1	
oa s	i->1	
oacc	e->31	
oad 	ö->3	
oade	 ->2	
oakl	u->1	
oakt	a->1	i->13	
oali	t->14	
oana	l->1	
oand	e->9	
oans	t->1	v->5	
oanv	ä->1	
oar 	e->1	k->1	o->1	s->2	
oard	,->1	
oare	s->1	
oate	r->1	
oavb	r->2	
oavs	e->8	i->2	
ob S	ö->2	
obak	,->1	s->1	
obal	 ->1	a->10	i->5	t->2	
obas	e->1	
obb 	e->1	o->1	
obb,	 ->2	
obby	,->1	a->1	b->1	g->2	i->2	m->1	n->3	v->1	
obeb	o->1	
obef	o->1	
obeg	r->5	
obeh	a->2	
ober	 ->8	o->50	t->1	ä->1	
obes	t->2	v->3	
obet	ä->1	
obil	i->7	
obin	,->1	
obje	k->1	
oble	m->183	s->1	
obli	g->14	
obod	a->3	
obse	r->2	
oc-d	i->1	
oc-t	r->1	
oca 	C->1	
oced	u->1	
ocen	t->94	
oces	s->109	
och 	"->3	(->1	-->6	0->1	1->21	2->13	3->7	4->10	5->3	6->2	7->6	8->11	9->4	A->4	B->6	C->4	D->4	E->35	F->15	G->7	H->3	I->14	J->2	K->9	L->8	M->5	N->2	O->2	P->15	R->3	S->25	T->8	U->1	V->2	W->1	X->1	a->290	b->119	c->10	d->588	e->210	f->320	g->91	h->161	i->231	j->152	k->197	l->93	m->278	n->79	o->95	p->115	r->188	s->440	t->152	u->106	v->229	y->7	Ö->7	ä->54	å->37	ö->43	
och)	D->1	
och,	 ->14	
och.	J->1	
och/	e->1	
ochI	 ->1	I->1	
ochi	s->1	
ochs	 ->1	
ocia	l->206	
ocie	r->1	t->1	
ocil	o->1	
ocio	e->3	
ock 	a->12	d->3	e->3	f->6	g->2	h->3	i->8	k->6	l->2	m->3	n->3	o->3	p->1	s->7	t->3	u->1	v->6	ä->1	å->2	
ock"	 ->1	
ock,	 ->8	
ock.	 ->1	J->1	K->1	
ocka	 ->3	d->3	n->2	r->1	
ockb	i->1	
ocke	r->4	t->1	
ockh	o->3	
ocks	 ->3	k->1	å->585	
ocku	p->5	
oco,	 ->1	
od a	d->1	n->1	t->3	v->4	
od b	i->1	ö->1	
od d	e->3	ä->1	
od e	f->2	n->1	
od f	a->1	i->2	r->1	å->1	ö->14	
od h	a->1	
od i	 ->5	d->2	n->2	
od j	a->1	o->1	
od k	o->2	
od l	e->1	
od m	e->3	i->1	y->1	
od n	y->1	
od o	m->2	
od p	r->1	å->3	
od r	e->1	ö->1	
od s	k->1	o->8	
od t	a->1	i->5	r->1	ä->1	
od u	p->1	
od v	i->2	
od ä	r->4	
od å	t->1	
od, 	e->1	f->1	m->1	n->1	v->1	
od.D	e->1	
od.F	a->1	
od.V	i->1	
od?-	 ->1	
oda 	a->4	c->1	e->1	f->8	g->1	h->2	i->1	k->1	l->2	n->1	o->3	p->2	r->4	s->1	t->3	v->3	
oda.	V->1	
odac	 ->3	"->1	-->1	
odaf	o->1	
odas	 ->2	.->3	
odda	.->1	
odde	 ->8	
odds	 ->1	
odel	b->1	l->12	
oden	 ->37	,->3	.->7	s->2	
oder	 ->13	,->4	.->6	a->1	m->1	n->39	s->4	t->1	
odet	 ->6	
odfi	l->1	
odi 	a->3	b->1	h->2	i->1	l->2	o->5	s->1	t->2	
odi,	 ->1	
odi.	S->1	V->1	
odi;	 ->1	
odif	i->5	
odig	a->3	t->1	
odin	s->1	
odis	 ->7	k->15	
odju	r->2	
odkä	n->89	
odla	r->3	
odli	g->12	n->2	
odo.	D->1	H->1	O->1	
odon	t->1	
odos	e->1	
ods 	a->1	b->1	i->1	l->1	o->1	p->18	s->4	t->1	v->1	ö->1	
ods,	 ->1	
ods.	 ->1	B->1	D->1	U->1	
ods;	 ->1	
odsN	ä->1	
odse	t->2	
odta	 ->10	.->1	g->17	r->3	s->7	
odto	g->2	
odty	c->6	
oduc	e->31	
odug	l->1	
oduk	t->53	
odwi	l->1	
oebb	e->1	
oedt	e->14	
oeff	e->2	i->1	
oeft	e->1	
oege	n->5	
oek 	s->1	
oeko	n->9	
oeli	g->1	
oelv	a->1	
oend	e->130	
oeni	g->4	
oens	e->4	
oerh	ö->12	
oers	ä->1	
oet 	a->1	
oeti	s->1	
oett	e->5	i->1	
of -	 ->1	
of a	v->1	
of e	l->1	x->1	
of f	ö->5	
of h	a->2	
of i	 ->1	n->2	
of k	u->1	
of l	i->1	
of o	c->2	
of s	o->4	
of t	h->1	
of u	t->1	
of ä	g->1	
of, 	h->1	m->1	o->1	s->1	
of.D	e->1	ä->1	
of.E	n->1	
of.J	a->1	
ofal	a->1	
ofan	t->2	
ofdr	a->1	
ofed	e->1	
ofel	b->1	
ofem	 ->2	
ofen	 ->13	,->5	.->2	
ofer	 ->17	"->1	,->5	.->5	n->4	
ofes	s->7	
offe	n->80	r->13	
offi	c->5	
offr	a->2	e->14	
ofhj	ä->1	
ofi 	o->1	s->1	
ofi,	 ->1	
ofil	 ->1	.->2	s->1	
ofin	 ->1	-->2	a->1	
ofis	k->1	
ofob	i->1	
ofre	d->1	
ofrå	n->3	
ofsi	t->1	
ofst	r->1	ö->2	
oft 	l->1	
ofta	 ->49	.->1	r->3	s->1	
oful	l->2	
oför	a->1	d->2	e->6	f->1	k->1	l->2	m->5	s->3	t->2	ä->2	
og 1	9->1	
og a	k->1	t->4	v->1	
og b	a->1	e->3	
og d	e->4	i->1	
og e	n->3	r->1	t->3	v->1	
og f	a->1	r->1	ö->3	
og h	a->2	e->1	ä->1	
og i	 ->8	n->1	
og k	a->1	o->3	
og l	a->4	ä->1	
og m	a->1	e->9	å->2	
og n	i->1	o->1	
og o	c->2	m->2	
og p	a->1	å->1	
og r	e->3	å->1	
og s	i->1	o->4	t->2	
og t	i->3	
og u	p->9	
og v	i->1	
og ä	r->1	
og å	t->1	
og ö	k->1	
og, 	i->1	o->1	v->1	
og.D	a->1	e->1	
og.F	r->1	ö->1	
og.H	a->1	
og.J	a->2	
og.M	e->1	ö->1	
og.N	ä->1	
og.S	a->1	
oga 	a->5	f->5	m->2	p->1	s->1	ö->1	
oga,	 ->1	
oga.	J->1	V->1	
ogad	.->1	e->2	
ogam	 ->1	,->1	
ogan	d->11	s->1	t->1	
ogar	 ->8	,->1	.->1	n->7	
ogat	 ->3	i->1	
ogau	 ->7	,->5	.->1	M->1	b->1	s->3	
ogbe	r->1	
oge 	f->1	
oge,	 ->1	
ogen	 ->10	,->2	.->3	a->2	h->27	o->2	t->2	
oger	 ->2	
oget	 ->2	
oggr	a->12	
ogi 	-->2	o->2	
ogi.	.->1	V->1	
ogik	 ->1	,->2	.->3	e->2	
ogin	,->1	
ogis	k->34	
ogjo	r->1	
ogku	l->1	
ogm 	e->1	
ogma	t->1	
ogra	f->14	m->238	
ogre	s->1	
ogri	k->1	
ogru	n->3	
ogs 	-->1	a->5	b->1	d->1	e->1	i->3	k->2	m->3	n->1	o->2	p->1	s->1	t->1	u->3	
ogs,	 ->2	
ogsa	r->1	v->1	
ogsb	r->6	
ogse	r->1	
ogsf	a->1	
ogsk	o->1	
ogso	m->1	
ogsp	o->1	
ogss	e->4	
ogsu	t->1	
ogsv	å->1	
ogsä	g->2	
ogue	i->1	
ogyn	n->1	
ogår	d->1	
ogör	 ->1	a->4	e->3	s->1	
ohan	d->3	
oher	e->1	
ohja	m->1	
ohjä	l->1	
ohol	,->1	
ohäm	m->1	
ohöv	l->1	
oige	n->1	
oij-	v->1	
oins	k->2	
oint	r->4	
oire	 ->1	,->1	-->1	
oirm	o->1	
ois 	M->1	
oise	 ->1	
oisk	 ->1	
oiss	y->1	
oist	i->2	
ojal	a->2	i->5	
ojek	t->64	
ojka	n->1	
ojko	t->1	
ojos	 ->1	
ojus	t->6	
ojäm	l->5	n->2	
ok a	v->1	
ok d	e->1	
ok f	ö->2	
ok g	j->1	
ok h	e->1	
ok i	 ->1	
ok m	e->1	
ok o	c->2	m->7	
ok s	a->1	k->1	o->2	
ok t	i->1	
ok ä	r->2	
ok, 	d->1	f->1	k->1	m->1	s->1	
ok.D	e->1	
ok.H	u->1	
ok.J	a->1	
ok.T	a->1	
ok.V	i->1	
oka 	h->1	s->1	
okal	 ->7	a->31	i->3	p->1	t->2	
okas	t->1	
okat	 ->2	.->1	e->2	
oken	 ->31	,->1	.->4	:->1	s->1	
oker	i->1	
okig	 ->1	t->1	
okla	d->1	m->1	n->2	r->12	
oko 	C->5	
okol	l->26	
okon	f->1	t->2	
okor	 ->1	
okra	t->138	
okre	d->2	
okri	g->1	t->1	
okrä	n->1	
oksl	u->1	
okst	a->1	
okt 	d->2	s->2	v->1	
okto	b->8	
okul	t->3	
okum	e->46	
okun	n->2	s->1	
okus	 ->1	.->1	e->3	
okän	d->1	s->1	
ol a	t->1	v->1	
ol b	e->1	
ol d	ä->1	
ol f	ö->2	
ol i	 ->2	n->1	
ol m	e->1	å->1	
ol o	c->9	
ol s	o->4	
ol t	i->1	
ol v	i->1	
ol, 	d->1	e->1	i->1	o->2	p->1	t->1	
ol- 	o->1	
ol-f	ö->1	
ol.D	e->1	
ol.E	t->1	u->1	
ol.H	e->1	
ol.K	ä->1	
ol.M	e->1	
ol; 	f->1	
ola 	d->2	f->1	s->1	v->1	ä->1	
ola,	 ->1	
olad	d->1	
olag	 ->3	,->1	e->8	l->4	
olan	 ->5	,->1	.->2	?->1	a->4	h->4	
olar	 ->12	,->1	.->2	n->8	s->2	
olav	t->1	
olbe	s->2	
olda	t->2	
oldi	o->5	
ole 	p->1	
olem	i->1	
olen	 ->28	,->5	.->7	s->8	
oler	a->17	e->7	i->1	
oleu	m->1	
olf 	H->2	
olfe	n->4	
olfr	å->1	
olfs	t->3	
olfö	r->2	
olib	a->1	
olic	y->4	
olid	a->30	e->3	
olig	 ->4	,->1	a->2	e->6	t->5	
olik	 ->1	.->1	:->1	a->116	e->2	h->7	t->5	
olin	t->1	
olis	,->1	.->1	;->1	a->1	e->8	i->1	k->6	m->3	s->2	v->1	
olit	a->1	i->533	
oliv	 ->2	.->1	
olja	 ->4	,->2	.->1	n->3	
olje	b->13	f->1	i->3	k->2	s->1	t->10	u->2	
olk 	a->1	b->2	h->1	i->2	o->2	r->1	s->3	t->1	u->1	
olk,	 ->1	
olk.	A->1	D->1	M->1	O->1	V->4	
olka	 ->4	d->1	r->5	s->6	t->1	
olke	n->6	s->1	t->14	
olkf	r->1	
olkg	r->2	
olkh	ä->9	
olkl	i->1	
olkn	i->57	
olko	m->6	n->1	
olkp	a->10	
olkr	e->4	ä->1	
olks	 ->3	t->1	w->1	ä->1	
olkv	a->2	
oll 	-->1	E->1	a->21	d->2	f->8	g->2	i->19	k->2	m->1	n->3	o->7	p->1	s->12	u->1	v->4	ä->3	ö->5	
oll!	J->1	
oll,	 ->20	
oll-	 ->1	
oll.	D->5	E->1	F->2	H->1	I->2	J->3	K->2	M->1	P->2	S->2	T->2	U->1	V->4	
oll:	 ->1	
olla	n->1	r->9	
olle	g->196	k->10	n->27	r->60	t->16	
ollf	u->1	
olli	s->3	
ollm	a->1	y->1	ä->1	ö->2	
olln	i->2	
ollo	m->1	r->1	
ollr	i->1	
olls	b->1	y->3	
ollu	t->15	
ollv	e->1	
olly	w->1	
olm 	d->1	
olm,	 ->1	
olm.	H->1	
oln 	o->1	
olog	,->1	i->30	
olon	i->1	
olor	 ->2	,->1	
olos	s->1	
olpe	 ->1	
ols 	a->1	m->1	u->1	
olsa	v->1	
olsb	u->1	
olsf	a->1	ö->1	
olsi	t->1	
olsk	a->4	e->1	
olsp	r->1	
olss	y->1	
olst	v->1	
olsu	t->1	
olsv	ä->1	
olt 	ö->6	
olta	 ->3	
olth	e->2	
olun	t->4	
olut	 ->38	a->3	i->100	
olv 	å->1	
olve	r->9	t->1	
olyc	k->48	
olym	 ->2	e->2	p->1	
olzm	a->2	
oläm	p->5	
olös	t->2	
om "	E->2	K->1	n->1	o->1	v->1	ö->1	
om -	 ->10	
om 1	 ->1	5->1	6->1	9->2	
om 2	0->2	8->1	
om 3	-->2	1->1	5->3	
om 4	0->3	5->1	
om 5	b->1	
om 6	,->1	
om A	g->1	h->1	l->2	m->3	p->1	t->1	
om B	S->1	a->1	e->6	l->1	o->1	r->2	
om C	E->1	e->1	o->2	
om D	a->4	e->1	i->1	u->1	
om E	G->3	M->1	U->19	h->1	l->1	r->1	t->1	u->72	
om F	B->1	P->1	l->1	r->2	ö->4	
om G	U->1	a->1	e->2	o->2	r->2	
om H	a->5	e->1	i->1	
om I	N->1	n->1	r->1	s->1	t->2	
om J	o->2	ö->2	
om K	a->1	o->5	
om L	a->6	i->1	l->1	
om M	a->2	c->2	
om N	e->1	
om O	f->1	
om P	P->1	a->3	o->4	r->1	
om R	a->1	i->1	o->1	
om S	E->1	c->2	e->2	j->1	k->1	p->1	
om T	a->1	h->3	i->2	o->2	u->4	
om V	ä->1	
om W	a->2	i->1	
om a	 ->1	b->2	d->2	g->4	l->53	m->2	n->66	p->1	r->21	s->3	t->334	v->39	
om b	)->1	a->7	e->127	i->12	l->9	o->15	r->13	u->3	y->2	ä->7	å->5	ö->16	
om c	)->1	a->1	e->1	h->2	o->1	
om d	a->6	e->617	i->17	j->1	o->5	r->16	u->1	y->1	ä->8	å->5	ö->3	
om e	f->8	g->5	j->1	k->5	l->2	m->1	n->182	r->14	t->98	u->8	x->15	
om f	a->31	e->2	i->43	j->1	l->11	o->21	r->60	u->5	y->2	ä->2	å->9	ö->208	
om g	a->7	e->48	i->3	j->10	l->1	o->8	r->16	ä->22	å->11	ö->34	
om h	a->195	e->55	i->14	j->6	o->14	u->34	y->1	ä->35	å->8	ö->7	
om i	 ->94	c->4	d->1	f->2	g->1	h->1	n->185	s->1	
om j	a->133	o->6	u->13	ä->3	
om k	a->63	e->1	l->2	o->186	r->26	u->9	v->1	ä->12	ö->2	
om l	a->18	e->38	i->40	j->1	o->1	y->6	ä->24	å->3	ö->2	
om m	a->95	e->48	i->30	o->14	u->1	y->15	ä->14	å->32	ö->51	
om n	a->13	e->4	i->62	o->1	u->25	y->7	ä->12	å->26	ö->2	
om o	a->1	b->2	c->36	f->7	g->1	l->6	m->41	n->1	r->17	s->4	t->1	
om p	a->23	e->7	l->4	o->7	r->22	u->2	å->38	
om r	a->56	e->88	i->14	o->1	u->3	y->2	ä->15	å->35	ö->17	
om s	.->1	a->47	c->1	e->16	i->11	j->4	k->127	l->6	m->3	n->3	o->6	p->11	t->81	u->4	v->3	y->18	ä->20	å->26	ö->3	
om t	.->3	a->20	i->73	j->3	o->10	r->26	u->1	v->5	y->11	ä->4	
om u	n->39	p->35	r->8	t->75	
om v	a->59	e->25	i->337	o->5	r->1	u->1	ä->13	å->17	
om y	r->1	t->3	
om Ö	s->4	
om ä	g->4	n->26	r->176	t->1	v->14	
om å	k->1	l->2	r->4	s->5	t->22	
om ö	a->1	k->3	m->1	n->1	p->7	r->1	s->2	v->17	
om!T	r->1	
om".	D->1	
om) 	o->1	
om);	 ->1	
om, 	a->5	d->7	e->4	f->1	g->1	h->3	i->4	j->2	k->1	l->1	m->2	n->2	o->5	p->1	s->4	t->1	u->4	v->4	ä->6	
om- 	o->1	
om. 	D->1	H->1	
om.A	v->1	
om.D	e->9	ä->1	
om.E	K->1	x->1	
om.H	e->1	u->1	
om.I	n->1	
om.J	a->7	
om.M	e->4	
om.N	ä->1	
om.O	c->1	
om.S	t->1	å->1	
om.V	i->3	
om/r	i->1	
omI.	 ->1	
omad	e->1	
omag	n->1	
oman	e->1	o->2	
omar	 ->9	,->3	.->2	b->2	e->5	k->1	n->8	
omat	e->1	i->18	
omb 	h->1	
omb.	A->1	
omba	d->1	r->1	t->2	
ombe	d->1	n->1	r->2	s->2	t->2	x->1	
ombi	n->1	
ombl	i->5	
ombn	i->1	
ombo	r->1	
ombr	o->2	
ombu	d->12	
omde	f->1	
omdi	r->1	
omdr	i->6	
omdö	m->2	
omed	e->18	g->2	v->1	
omen	 ->10	,->3	.->1	e->5	t->5	
omer	 ->2	,->3	a->4	n->1	
omes	,->1	
omet	 ->1	e->1	
omeu	r->4	
omfa	t->83	
omfl	y->1	
omfo	r->4	
omfå	n->2	
omfö	r->162	
omge	r->1	
omgi	c->1	v->2	
omgr	i->4	
omgå	 ->1	.->1	e->1	n->5	r->4	t->2	
omhu	l->1	
omi 	-->1	a->1	m->5	o->12	ä->1	
omi,	 ->2	
omi.	D->2	F->1	
omi?	 ->1	
omie	r->8	
omin	 ->20	,->2	.->5	a->1	e->10	s->3	
omis	k->215	s->22	t->5	
omkr	i->15	
omla	s->1	
omli	g->18	
omlo	k->2	
omlä	s->2	
omma	 ->102	,->1	.->3	n->55	r->3	s->1	
omme	l->15	n->84	r->730	t->5	
ommi	s->1150	t->103	
ommo	n->1	r->2	
ommu	n->33	
ommö	b->1	
omna	 ->13	,->1	.->1	n->1	r->28	s->1	
omof	o->1	
omog	e->2	
omor	a->1	d->7	g->2	
omos	e->1	
ompa	s->1	
ompe	n->10	t->11	
ompl	a->1	e->28	i->16	
ompo	n->4	
ompr	o->22	ö->8	
omri	n->1	
omru	m->2	
områ	d->316	
omrö	s->42	
oms 	f->1	s->1	
oms-	 ->2	,->1	
omsa	 ->3	r->1	
omsb	r->1	
omsf	r->3	u->1	
omsg	r->1	
omsh	e->1	
omsk	i->1	
omsl	a->3	u->3	
omsn	i->11	
omso	r->9	
omsp	l->1	ä->1	
omsr	ä->1	
omst	 ->7	e->8	f->1	h->1	k->1	o->86	r->15	ä->35	å->2	
omsv	e->1	ä->1	
omsy	r->3	
omsä	t->8	
omta	l->1	
omtä	n->1	
omul	l->1	
omva	n->5	
omvä	g->2	l->4	n->5	x->1	
omán	,->1	
omäs	s->1	
omål	 ->2	e->1	
omé 	o->1	p->1	
oméa	v->1	
omék	o->1	
omés	 ->1	
omöj	l->16	
on (	A->5	f->2	
on -	 ->5	
on 1	2->5	9->1	
on 3	4->1	
on 5	2->1	7->1	
on A	c->1	
on B	o->1	
on E	i->1	
on H	a->1	
on I	 ->1	
on P	r->2	
on V	I->2	a->3	
on W	o->17	
on a	l->2	n->13	p->1	r->1	t->6	v->27	
on b	e->8	i->1	l->1	o->1	ä->2	ö->1	
on c	h->1	
on d	e->3	ä->8	å->1	
on e	f->6	l->2	n->5	t->1	u->1	
on f	a->1	o->1	r->5	u->1	å->1	ö->33	
on g	e->3	r->1	å->8	ö->1	
on h	a->13	o->1	ä->3	ö->1	
on i	 ->29	d->1	n->17	
on j	a->1	u->3	
on k	a->13	l->12	o->15	
on l	a->3	i->2	y->1	ö->1	
on m	.->1	e->19	i->2	o->4	y->1	å->2	ö->2	
on n	e->1	i->1	y->4	ä->2	
on o	c->41	f->1	l->3	m->20	r->2	v->1	
on p	e->2	l->2	r->1	å->16	
on r	e->3	i->2	o->1	ä->3	
on s	a->4	e->1	k->13	o->72	p->1	t->7	y->1	ä->2	å->7	
on t	a->4	i->22	j->1	r->1	y->1	ä->1	
on u	n->2	p->5	r->1	t->3	
on v	a->1	e->4	i->6	å->1	
on ä	n->1	r->11	
on å	r->2	t->3	
on ö	v->1	
on" 	p->1	
on) 	(->2	
on, 	5->1	D->1	L->1	O->1	P->1	S->1	a->2	b->3	d->5	e->7	f->3	h->2	i->4	k->3	m->4	n->2	o->12	p->1	s->9	t->1	u->1	v->4	ä->3	
on- 	o->1	
on-H	a->1	
on. 	D->1	I->1	O->1	R->1	
on.1	4->1	
on.A	v->1	
on.B	r->1	
on.D	E->1	e->18	ä->2	å->1	
on.E	n->2	v->1	
on.F	l->1	r->1	ö->3	
on.G	ä->1	
on.H	a->1	e->6	
on.I	 ->7	
on.J	a->14	
on.K	o->2	
on.L	å->1	
on.M	e->1	i->2	ö->1	
on.N	i->2	
on.O	m->3	
on.S	a->1	e->1	o->2	å->1	
on.T	i->1	r->1	
on.U	n->1	
on.V	a->5	i->11	
on.Å	 ->1	
on/å	r->2	
on: 	D->1	a->1	i->1	
on; 	v->1	
on? 	D->1	I->1	
on?D	e->1	
on?J	a->1	
on?K	a->2	o->1	
on?V	i->1	
on?Ä	v->1	
onNä	s->1	
ona 	a->8	d->5	e->2	h->1	i->1	n->1	o->1	s->1	t->4	v->2	
onad	e->7	
onak	r->1	
onal	 ->16	,->2	-->2	.->4	a->44	e->5	f->3	i->28	l->1	p->40	r->4	s->7	t->1	u->1	
onan	d->1	s->1	
onap	r->2	
onar	 ->7	,->1	
onas	 ->3	
onat	 ->2	,->2	.->1	i->1	
onaz	i->2	
onbe	h->1	
onbl	i->15	
once	n->31	p->7	r->2	
onci	s->2	
onck	h->14	
ond 	c->1	f->4	k->1	s->2	
onda	 ->3	g->2	
onde	 ->5	.->1	n->45	r->69	
ondg	å->2	
ondi	t->1	
ondm	e->3	
ondo	.->1	n->4	
onds	k->1	p->3	
ondu	p->1	
one 	a->2	b->1	d->1	e->1	f->1	g->1	h->1	i->5	j->1	k->2	l->1	n->4	o->1	r->1	s->1	t->1	v->2	
one-	M->1	s->1	
onel	l->277	
onem	a->3	
onen	 ->883	!->1	"->1	)->1	,->103	.->137	:->1	;->3	?->4	J->2	s->375	t->5	
oner	 ->284	,->42	.->45	;->1	?->4	N->1	a->15	i->11	l->2	n->181	s->5	
onet	.->1	a->1	ä->6	
onfe	d->1	r->170	s->1	
onfi	d->2	s->2	
onfl	i->16	
onfr	o->1	
onge	n->1	
ongi	v->2	
ongr	e->1	
ongs	b->1	
onhu	n->1	
oni 	o->2	s->1	
oni.	(->1	
onia	l->1	
onik	-->1	
onin	d->1	g->5	
onis	e->15	k->13	m->3	t->2	
onit	o->1	
onju	n->1	v->1	
onjä	r->1	
onkr	e->58	
onku	r->285	
onla	m->1	
onli	g->34	
onmä	r->2	s->1	
onmö	t->2	
onna	m->1	
onnä	e->1	
onod	l->3	
onok	u->3	
onom	 ->22	,->2	.->4	e->4	i->283	
onop	o->17	
onra	d->1	
ons 	b->1	f->1	i->1	p->1	r->1	s->2	t->2	v->2	
ons-	 ->4	
onsa	f->2	n->1	r->8	v->1	
onsb	o->1	r->1	
onsd	a->5	i->1	o->1	ö->1	
onse	k->61	r->7	
onsf	o->1	r->2	u->1	ö->19	
onsh	a->1	i->8	
onsi	n->13	
onsk	a->2	o->5	r->1	u->6	
onsl	e->11	ä->1	
onsm	e->4	o->1	ä->1	ö->1	
onsn	i->2	
onso	l->3	r->1	
onsp	a->1	l->2	o->3	r->6	
onsr	a->1	e->3	o->1	ä->12	
onss	a->7	c->1	e->1	k->1	t->2	y->5	
onst	 ->1	,->1	a->45	e->3	i->29	j->1	r->42	
onsu	l->5	m->63	n->3	p->1	t->3	
onsv	i->1	
onsä	g->1	m->1	
onså	t->1	
ont 	a->1	o->1	
ont.	S->1	
onta	i->1	k->17	l->3	m->2	n->5	t->1	
onte	l->1	n->3	r->12	x->1	
onti	 ->10	!->3	,->2	.->2	n->46	
onto	r->7	
ontr	a->7	e->2	o->184	
onve	n->24	r->5	
onvi	k->4	
onym	 ->2	.->1	a->1	i->1	
onzá	l->1	
onär	 ->65	!->32	,->74	.->11	e->65	s->1	
onår	i->1	
onöd	i->11	
oo f	r->1	
ood 	o->1	
oodf	i->1	
oods	 ->1	
oodw	i->1	
ooij	-->1	
ool,	 ->1	
oomr	å->1	
oope	r->1	
oos 	a->1	
op a	l->1	
op b	e->1	
op d	e->1	
op f	ö->1	
op o	c->1	m->1	
op p	e->1	
op s	i->1	k->1	
op t	i->1	
op u	t->1	
op ä	n->1	
op, 	A->3	e->1	o->1	p->1	
op-s	h->1	
op.D	e->1	
op.I	n->1	
op.J	a->1	
op.S	o->1	
opa 	-->2	a->8	b->1	d->1	e->4	f->6	h->11	i->9	k->10	m->13	n->1	o->19	p->3	r->2	s->26	t->4	u->4	v->7	ä->11	
opa!	A->1	F->1	
opa"	.->1	
opa,	 ->36	
opa.	.->2	1->1	D->15	E->2	F->3	H->6	I->2	J->8	M->3	N->1	O->1	P->1	R->1	T->2	U->1	V->10	Ä->1	
opa;	 ->1	
opa?	H->1	V->2	
opaN	ä->1	
opad	e->2	
opag	a->3	e->1	r->1	
opak	o->1	
opam	i->1	
opan	i->1	
opap	a->166	
opar	 ->3	t->2	å->1	
opas	 ->48	
opat	j->1	
opav	a->3	
opei	s->712	
oper	a->12	e->1	
opet	 ->2	
opia	 ->1	
opie	n->3	r->1	
opil	o->1	
opin	i->4	
opla	s->1	
opol	 ->15	,->3	.->2	;->1	a->1	f->3	i->3	k->1	s->4	
opor	t->9	
opou	l->5	
opp 	-->1	a->2	f->8	h->2	i->1	p->1	s->1	
opp,	 ->1	
opp.	.->1	
oppa	 ->5	d->2	r->1	s->99	
oppe	 ->1	n->8	t->10	
oppl	a->4	i->2	ö->1	
oppm	ö->12	
oppn	i->12	
oppo	n->3	r->2	s->2	
opra	k->1	
opro	g->2	j->1	p->2	t->2	
opti	m->7	o->1	
opul	a->1	i->4	ä->2	
opyr	i->1	
opå 	b->1	
opé 	o->1	
opée	r->9	
or -	 ->3	
or F	r->1	
or M	o->2	
or T	e->1	s->2	
or a	l->1	n->3	r->1	t->85	v->10	
or b	e->14	i->2	l->1	o->1	r->2	ö->3	
or c	h->1	
or d	e->21	j->1	ä->7	ö->2	
or e	f->2	g->1	l->4	n->3	r->1	u->1	
or f	a->4	i->1	o->2	r->7	ö->27	
or g	a->1	e->3	r->1	ä->1	ö->1	
or h	a->12	i->1	j->3	ä->2	ö->1	
or i	 ->30	n->29	
or j	a->23	o->2	u->1	
or k	a->5	o->2	
or l	e->1	i->2	ö->1	
or m	a->7	e->12	i->1	y->1	ä->2	å->4	
or n	i->4	o->1	ä->1	
or o	c->70	m->16	r->2	
or p	e->1	o->2	r->1	å->20	
or r	e->5	o->1	
or s	a->2	e->3	j->1	k->4	o->94	t->2	y->1	å->3	
or t	i->24	j->1	r->1	
or u	n->1	p->8	r->1	t->14	
or v	a->5	e->2	i->12	ä->2	
or ä	n->3	r->11	v->1	
or ö	v->2	
or) 	o->1	
or, 	a->1	b->2	e->3	f->3	g->2	h->1	i->6	k->3	m->13	n->2	o->11	p->1	r->2	s->20	t->2	u->5	v->2	ä->4	
or. 	D->1	
or..	(->1	
or.A	l->1	
or.B	r->1	
or.D	e->23	ä->1	
or.E	t->1	
or.F	e->1	r->3	ö->6	
or.G	e->1	
or.H	e->2	u->1	
or.J	a->12	
or.K	a->1	o->2	
or.L	i->1	
or.M	a->1	e->2	y->1	
or.N	a->1	y->1	ä->1	
or.O	c->2	
or.R	e->1	
or.S	a->2	
or.T	i->1	y->1	
or.V	e->1	i->6	å->1	
or.Ä	v->1	
or.Ö	V->1	
or: 	d->1	f->1	o->1	t->1	
or; 	j->1	
or?,	 ->1	
or?H	a->1	u->1	
or?Ä	r->1	
ora 	1->1	a->9	b->6	d->5	e->5	f->47	g->7	h->2	i->8	k->3	m->4	n->1	o->11	p->13	r->3	s->18	t->5	u->3	v->4	å->3	
ora,	 ->2	
ora.	E->1	M->1	V->1	
ora?	A->1	
orad	 ->2	e->3	
oral	 ->1	,->1	e->1	i->5	
oran	d->1	
orar	 ->4	
orat	 ->7	,->3	.->2	e->13	i->4	o->3	s->1	
orbe	r->1	t->1	
orbi	h->1	
orbr	i->14	o->1	
orce	 ->1	
orcy	k->4	
ord 	-->1	I->2	a->4	b->1	e->1	f->6	i->6	j->1	k->3	m->1	n->1	o->11	s->6	t->4	v->3	
ord,	 ->4	
ord-	f->1	
ord.	B->1	E->1	U->1	V->2	
ord:	 ->2	
orda	 ->5	,->1	d->1	l->6	m->4	n->3	r->2	
ordb	r->57	ä->10	
orde	 ->100	,->1	.->2	a->1	n->31	r->6	s->5	t->22	u->1	
ordf	ö->216	
ordi	n->1	r->2	s->4	t->1	
ordk	u->1	
ordl	a->1	i->5	
ordm	å->1	
ordn	a->28	i->155	
ordo	n->65	
ordr	a->18	e->1	i->5	
ords	k->1	u->1	
ordt	i->1	y->1	
ordv	r->1	ä->2	
ore 	b->2	d->5	e->6	f->3	h->1	i->3	l->1	m->2	o->3	p->1	t->1	v->1	ö->1	
orea	 ->3	l->2	
oreb	o->1	
ored	l->1	
oreg	l->1	
orel	a->1	
oren	 ->17	,->1	.->4	a->19	i->9	z->19	
orer	 ->30	,->2	.->4	a->4	n->10	
ores	t->1	
oret	 ->1	i->2	
orfö	r->2	
org 	a->1	o->7	s->1	t->1	
orga	n->93	r->168	
orge	 ->1	,->1	r->3	
orgl	i->3	
orgm	ä->2	
orgo	n->37	
orgs	f->1	
orha	v->1	
orhe	t->1	
ori 	8->2	o->2	s->1	v->1	
oria	 ->6	,->2	.->2	
orie	l->5	n->13	r->10	t->3	
orig	i->2	
orik	 ->1	,->1	.->1	e->1	t->3	
orim	l->5	
orin	d->2	g->1	o->7	
oris	 ->1	e->2	k->35	m->2	o->3	t->8	
orit	a->1	e->104	l->1	
oriu	m->10	
ork 	v->1	
orka	,->1	n->3	p->1	
orkn	i->1	
orld	 ->1	
orli	g->2	
orlu	n->3	
orlä	r->1	
orm 	a->26	b->1	d->2	e->1	f->3	i->3	j->1	k->4	l->1	o->3	p->1	s->7	v->3	ä->1	ö->1	
orm,	 ->9	
orm.	D->1	E->1	M->1	N->1	S->1	V->1	Ä->1	
orm:	 ->1	
orma	 ->24	.->1	d->1	l->11	n->5	r->23	s->3	t->77	
orme	l->16	n->23	r->131	
ormf	ä->1	ö->2	
ormi	s->1	
ormn	i->26	
ormo	n->1	
ormp	a->1	r->14	
orms	t->1	
ormt	 ->7	
ormu	l->18	
ormå	t->1	
orn 	-->2	b->1	e->2	f->3	i->2	k->1	o->5	s->3	u->1	ä->2	
orn)	.->1	
orn,	 ->12	
orn.	D->4	F->3	H->1	K->1	M->1	
orn?	A->1	
orna	 ->69	,->10	.->12	?->1	s->7	
orne	t->1	
orno	g->2	
orns	 ->4	
oro 	-->1	E->1	b->1	d->1	f->5	i->3	l->1	n->2	o->4	p->1	s->12	ä->3	ö->1	
oro,	 ->4	
oro.	A->1	B->1	F->2	J->2	O->1	T->1	V->1	
oroa	 ->3	d->5	n->9	r->4	
orol	i->6	
oron	 ->5	
oros	m->4	
orov	ä->2	
orpe	t->2	
orpo	l->1	
orpu	s->5	
orr?	V->1	
orra	 ->4	i->2	
orre	c->1	k->27	n->1	s->1	y->3	
orri	d->2	
orru	m->2	p->7	
ors 	a->1	b->3	d->6	e->1	f->5	g->1	h->7	i->7	k->2	l->2	o->4	p->1	r->2	s->6	t->3	u->1	y->1	ö->1	
ors,	 ->7	
ors.	D->5	J->1	M->1	T->1	U->1	V->2	
orsa	k->36	n->1	
orsb	e->1	
orsd	a->8	
orse	 ->3	,->1	.->2	l->1	
orsi	n->1	
orsk	a->8	n->35	r->1	
orsl	a->2	i->1	
orst	 ->1	ä->2	
orsö	v->1	
ort 	-->1	E->1	a->42	b->6	d->14	e->15	f->21	g->5	h->7	i->13	k->7	l->2	m->7	n->8	o->35	p->9	r->4	s->37	t->10	u->6	v->7	ä->2	å->1	ö->2	
ort)	 ->1	
ort,	 ->26	
ort-	 ->1	s->2	
ort.	D->8	E->1	I->1	J->3	L->1	N->1	R->1	S->1	U->1	V->3	
ort:	 ->1	
ort?	J->1	
ortN	ä->1	
orta	 ->5	b->1	d->1	m->1	s->1	
ortb	e->2	i->1	
ortd	i->1	
orte	n->48	r->64	t->19	
ortf	a->97	e->1	r->1	ö->1	
ortg	r->1	å->5	
orti	o->9	
ortk	o->2	
ortl	e->1	
ortm	a->1	o->1	
ortn	i->1	ä->1	
orto	m->6	n->9	
ortp	r->2	
orts	 ->25	,->3	.->2	a->12	e->6	i->5	k->1	ä->89	
ortu	g->97	n->2	t->1	
ortv	i->1	
orty	r->1	
orum	 ->4	,->1	e->1	
orv 	f->1	
orve	n->5	
orwe	l->1	
oräk	n->1	
orär	 ->1	t->1	
orät	t->10	
orêt	s->1	
orös	 ->1	a->2	t->1	
os D	a->1	
os E	G->1	u->1	
os F	P->1	
os O	z->1	
os R	E->1	
os a	l->3	n->1	t->1	v->1	
os b	e->11	l->1	
os d	e->13	
os e	n->3	x->1	
os f	a->1	ö->5	
os h	a->1	
os i	n->3	
os k	l->1	o->6	
os l	e->1	
os m	e->3	i->1	ä->1	å->1	
os n	ä->1	
os o	c->8	r->3	s->3	
os p	r->2	
os r	å->1	
os s	e->1	i->2	t->1	
os t	a->1	i->1	
os v	u->1	ä->1	å->1	
os y	t->1	
os å	s->1	
os! 	J->1	
os, 	a->1	h->1	k->1	
osam	t->2	
osan	n->1	
osat	s->1	t->3	
osed	d->1	
osen	r->1	
osex	u->1	
osfä	r->1	
osio	n->1	
osit	i->87	
osiv	 ->1	
osju	 ->1	
oske	p->3	
osko	p->3	
oskr	i->1	
oskv	a->1	
osky	d->1	
osla	v->1	
oslä	k->1	
osmo	l->1	m->3	
osni	e->2	
osof	i->5	
osor	,->1	
osov	o->60	
ospi	c->1	n->1	
oss 	-->1	a->39	b->1	d->19	e->16	f->16	g->4	h->6	i->29	k->3	l->3	m->12	n->6	o->29	p->13	r->2	s->29	t->16	u->8	v->13	y->1	ä->10	å->10	ö->3	
oss,	 ->15	
oss.	D->3	E->2	F->2	H->1	J->4	N->1	V->3	Ä->2	
oss:	 ->1	
oss?	.->1	V->1	
ossa	l->1	r->1	
osse	t->2	
ossi	l->3	
ossn	i->1	
osst	ê->1	
ost 	a->1	f->2	o->1	t->1	u->1	v->1	
ost-	b->5	
ost.	N->1	
osta	 ->9	,->2	d->4	r->4	s->1	t->3	
ostb	i->1	
oste	n->1	r->6	u->1	
osth	å->1	
osti	t->1	
ostn	a->108	
ostr	a->2	o->3	
osts	a->2	
ostv	e->1	
ostä	d->4	
osv.	 ->3	,->1	?->1	S->1	
osyn	l->1	
osys	t->4	
osäk	e->12	
osät	t->5	
osår	b->1	
ot -	 ->2	e->1	
ot 1	3->1	
ot 5	 ->1	
ot A	i->1	
ot D	a->1	
ot E	G->1	U->2	u->7	
ot F	r->1	ö->2	
ot G	r->1	
ot H	a->3	
ot I	s->1	
ot J	o->3	
ot K	a->1	
ot L	a->1	
ot M	o->1	
ot R	a->2	
ot S	o->1	
ot T	i->1	o->1	
ot U	N->1	
ot W	a->1	u->1	
ot a	b->1	i->1	l->7	n->10	r->2	t->16	v->20	
ot b	a->18	e->6	r->2	ä->1	å->1	
ot d	e->60	i->4	o->3	
ot e	k->1	l->1	n->13	r->3	t->7	x->4	
ot f	e->1	o->2	r->10	ö->17	
ot g	e->1	l->1	
ot h	a->4	e->1	i->1	u->2	ä->2	
ot i	 ->7	d->1	n->8	
ot j	a->4	
ot k	a->1	l->1	o->7	ö->1	
ot l	a->1	e->1	i->1	o->1	y->1	ä->3	
ot m	a->4	e->8	i->2	o->6	y->4	ä->2	å->1	
ot n	a->3	ä->3	å->1	
ot o	c->1	e->1	k->1	l->3	m->9	s->3	
ot p	a->2	e->1	o->3	r->5	u->1	å->4	
ot r	a->2	e->5	å->4	
ot s	a->1	e->1	i->3	j->1	k->6	l->5	n->1	o->55	p->3	t->8	u->2	v->3	y->1	ä->12	å->3	
ot t	a->3	e->1	i->3	v->1	
ot u	n->2	p->2	t->1	
ot v	a->6	e->5	i->11	ä->1	å->4	
ot y	t->1	
ot Ö	s->3	
ot ä	n->1	r->2	
ot å	r->1	t->1	
ot ö	k->2	v->4	
ot! 	D->2	J->2	N->1	S->1	V->1	
ot!D	e->1	
ot, 	Z->1	a->5	d->1	e->2	h->2	o->1	s->2	t->1	u->1	v->1	ä->3	
ot. 	7->1	
ot.A	l->1	
ot.D	e->2	
ot.F	r->2	
ot.J	a->2	
ot.S	l->1	
ot.V	i->1	
ot.Ä	n->1	
ot?N	e->1	
ota 	d->1	f->1	h->1	k->1	
otac	k->1	
otad	.->2	e->6	
otal	 ->4	,->1	-->3	F->1	a->14	b->2	e->1	f->5	i->2	s->6	t->6	v->1	
otan	;->1	d->1	
otar	 ->10	b->1	
otas	 ->8	.->1	
otat	 ->1	i->1	
otbi	l->1	
otbo	l->1	
ote 	Q->1	
otek	e->2	t->4	
otel	s->1	
oten	 ->25	.->3	s->2	t->6	
oter	 ->1	.->1	a->27	i->5	n->4	
otes	e->1	t->9	
otet	 ->7	i->1	
otfu	l->1	
otfä	r->1	s->1	
otgå	n->1	
oth-	B->7	
otha	r->3	
othe	r->1	
otik	a->7	
otil	l->17	
otio	n->1	
otis	 ->1	k->1	m->5	
otiv	 ->2	a->1	e->18	
otjä	n->1	
otni	n->17	
oto 	k->1	o->1	
oto-	p->1	
oto.	V->1	
otok	o->26	
otop	r->2	
otor	 ->1	.->2	c->4	i->2	
otos	 ->1	
otpa	r->4	
otpr	o->2	
otro	l->2	
otry	g->1	
ots 	a->34	d->20	e->1	i->1	k->1	m->1	p->1	r->1	s->2	t->1	v->1	
otsa	t->23	
otsp	å->2	
otst	r->1	y->3	å->12	
otsv	a->17	
otsy	s->1	
otsä	g->8	t->9	
ott 	a->5	b->3	d->2	e->3	f->5	h->2	i->4	m->4	n->3	o->5	p->3	r->2	s->11	u->1	ä->1	
ott,	 ->11	
ott.	D->2	F->1	I->1	J->1	L->1	M->1	O->3	Ä->1	
otta	 ->2	,->1	d->3	g->16	n->1	r->1	s->1	t->2	
otte	n->8	r->3	t->136	
ottg	ö->1	
otti	 ->1	
ottl	a->5	
ottm	å->1	
ottn	a->3	e->1	
otto	r->1	
otts	 ->3	b->5	d->1	f->1	l->17	m->2	o->2	p->1	r->1	
otul	l->1	
otum	 ->1	
otur	i->1	
otus	e->1	
otve	r->4	t->2	
otvi	k->1	l->1	v->1	
otyd	l->4	
otän	k->1	
otål	i->1	
otåt	g->3	
ou f	r->1	
ou o	c->1	
ouch	n->12	
ouk 	a->1	
oula	d->1	
oulo	s->5	
oumb	ä->4	
ounc	i->1	
ound	g->2	v->4	
oup 	,->1	d->1	
oura	 ->6	,->2	
ourg	 ->2	.->3	
ouri	.->1	
ourl	a->6	
ourn	a->2	e->1	
ours	 ->1	
ouse	w->1	
ousk	o->1	
outh	ä->2	
outi	e->1	
outn	y->1	
oux-	a->1	
ov a	t->1	v->15	
ov f	ö->4	
ov i	 ->1	n->1	
ov k	o->1	
ov n	y->1	
ov o	c->7	
ov p	å->9	
ov s	o->1	y->1	å->1	
ov t	i->8	
ov",	 ->1	
ov, 	a->1	n->1	ä->1	
ov. 	D->1	
ov.A	v->1	
ov.D	e->1	
ov.H	e->1	
ov.U	p->1	
ova 	a->2	
ovad	e->4	
ovak	i->1	
ovan	,->1	.->1	a->1	i->1	l->1	n->2	p->1	s->2	
ovar	 ->2	
ovat	 ->5	.->1	i->6	s->1	
ovem	b->11	
oven	 ->5	.->1	s->1	
over	 ->1	,->1	a->1	h->1	i->3	s->4	
ovet	 ->36	,->2	
ovic	 ->1	
ovil	j->2	l->2	
ovin	s->3	
ovis	 ->1	)->1	a->3	b->9	e->1	f->3	k->2	n->1	o->2	s->1	
ovje	t->1	
ovka	r->1	
ovko	n->1	
ovo 	(->2	T->1	a->1	b->1	f->3	h->1	i->1	k->2	m->1	o->7	t->1	u->1	v->1	ä->3	
ovo,	 ->11	
ovo.	-->1	A->1	D->2	E->1	F->1	H->1	K->1	L->1	M->1	O->1	V->1	
ovo?	 ->1	H->1	
ovoN	ä->1	
ovok	o->1	r->1	
ovor	d->2	
ovos	 ->7	
ovsi	d->1	
ovsk	o->2	
ovsm	a->2	ä->3	
ovst	e->1	
ovvä	r->2	
ovyt	t->1	
oväc	k->3	
oväd	e->1	r->1	
oväl	k->1	
ovän	l->1	
ovär	d->15	
oväs	e->1	
ovåd	l->1	
ovår	d->2	
ow t	i->1	
ow-h	o->1	
owe.	E->1	V->1	
ower	 ->1	,->2	
owis	 ->2	
owit	t->1	
own 	a->1	ä->1	
own,	 ->1	
ox o	c->1	
ox s	a->1	
ox!J	a->1	
ox, 	j->1	s->1	
oxal	 ->2	a->1	t->2	
oxid	 ->4	u->1	
oxin	 ->1	k->1	
oxis	k->1	
oxni	n->1	
oyal	 ->1	
oyds	 ->1	
oyol	a->2	
oämn	e->1	
oänd	l->4	
oäng	 ->1	.->1	s->2	t->8	
oår 	f->1	
oöns	k->1	
oöve	r->6	
p (k	r->2	
p , 	m->1	
p - 	o->2	s->1	
p Ca	d->1	
p Eu	r->1	
p Jö	r->1	
p Ti	b->1	
p al	l->7	
p an	s->3	t->1	v->1	
p at	t->11	
p av	 ->76	s->1	
p be	g->1	t->2	
p bi	d->1	
p bå	d->1	
p bö	r->2	
p de	 ->11	b->2	m->2	n->14	s->3	t->12	
p do	m->1	
p dä	r->3	
p ef	t->3	
p el	l->3	
p en	 ->11	l->1	
p et	t->6	
p ex	p->1	
p fo	r->1	
p fr	a->2	å->13	
p fu	l->1	
p få	t->1	
p fö	r->21	
p ge	n->2	
p gr	u->1	ä->1	
p ha	d->1	r->6	
p he	l->1	
p hu	v->1	
p hä	n->2	r->1	
p hö	g->1	
p i 	E->1	S->1	b->2	d->6	e->2	f->2	h->1	k->1	m->3	p->2	r->3	s->2	t->2	u->1	v->2	ä->1	
p id	é->1	
p ig	e->4	
p in	l->2	o->2	t->6	
p ka	n->1	
p ko	m->6	n->1	
p la	g->1	
p li	v->1	
p lä	g->1	m->1	n->1	
p ma	n->1	
p me	d->8	l->3	
p mo	t->4	
p må	s->2	
p na	t->1	
p ni	 ->1	
p ny	a->1	
p nä	r->1	
p nå	g->3	
p oc	h->23	
p ol	j->1	
p om	 ->8	
p or	d->2	
p pe	r->1	
p po	s->1	
p pr	i->1	o->2	
p på	 ->11	.->2	
p re	f->1	g->1	
p rä	c->1	t->2	
p rå	d->1	
p rö	s->1	
p sa	d->1	
p si	g->1	n->1	t->1	
p sj	ö->1	
p sk	a->5	u->1	y->1	
p so	m->21	
p st	ä->2	
p sä	r->1	t->1	
p så	v->2	
p ti	l->18	
p to	g->1	
p tr	e->1	
p tv	å->1	
p ty	d->1	v->1	
p un	d->3	
p up	p->1	
p ut	a->2	g->1	t->3	v->2	
p va	d->4	
p vi	d->2	l->2	
p vä	l->2	
p än	 ->1	d->1	n->1	
p är	 ->8	,->1	e->2	
p äv	e->1	
p ön	s->1	
p öv	e->1	
p" f	r->1	
p"!I	 ->1	
p", 	a->1	v->1	
p, A	r->3	
p, E	D->1	
p, a	n->1	v->1	
p, b	l->1	
p, d	e->3	ä->1	å->1	
p, e	f->3	n->5	
p, f	o->1	å->1	ö->1	
p, g	e->1	
p, h	a->1	e->2	
p, i	 ->1	n->1	
p, j	u->1	
p, l	i->1	
p, m	e->3	i->1	
p, n	u->1	
p, o	c->6	m->1	
p, p	å->1	
p, r	i->1	
p, s	o->2	ä->1	
p, u	t->1	
p, v	a->1	i->2	
p, ä	v->1	
p-sh	o->1	
p. S	k->1	
p. s	ä->1	
p. t	r->1	
p..(	F->1	
p.Ah	e->1	
p.Da	g->1	
p.De	 ->1	n->2	t->12	
p.Ef	t->1	
p.Eu	r->1	
p.Fa	k->1	
p.Hä	r->1	
p.I 	a->1	d->1	o->1	
p.In	r->1	
p.Ja	g->12	
p.Me	n->1	
p.På	 ->1	
p.Sj	ä->1	
p.Sl	u->1	
p.So	m->1	
p.Ti	l->1	
p.Vi	 ->6	l->1	s->1	
p.g.	a->1	
p.Än	d->1	
p.Äv	e->1	
p: K	o->1	
p?Hu	r->1	
pa -	 ->3	
pa O	L->1	
pa W	a->1	
pa a	l->3	n->4	r->7	t->7	v->1	
pa b	e->7	ä->1	
pa d	a->1	e->27	i->2	r->1	ä->2	
pa e	f->2	k->1	l->1	n->29	r->1	t->14	u->2	x->2	
pa f	i->1	l->2	o->2	r->3	å->1	ö->20	
pa g	e->4	l->1	
pa h	a->11	e->1	o->1	å->1	ö->2	
pa i	 ->10	h->1	m->1	n->11	
pa j	ä->1	
pa k	a->5	l->1	o->10	r->3	u->2	v->2	
pa l	a->1	u->1	
pa m	a->1	e->10	i->6	o->1	ä->5	å->4	ö->2	
pa n	a->1	y->5	ä->1	å->5	
pa o	c->22	f->2	l->1	m->1	r->1	s->2	
pa p	a->1	e->2	l->1	o->1	r->2	å->4	
pa r	e->5	ä->3	
pa s	i->2	k->6	n->2	o->20	p->2	t->3	u->1	y->6	å->3	
pa t	a->3	e->2	i->12	r->4	v->2	y->2	
pa u	n->4	r->2	t->2	
pa v	a->1	e->1	i->4	ä->2	å->2	
pa y	t->1	
pa ä	n->1	r->11	
pa å	t->1	
pa ö	v->1	
pa!A	v->1	
pa!F	r->1	
pa".	J->1	
pa, 	K->1	S->1	b->1	d->5	e->3	f->1	h->1	i->1	n->1	o->12	p->1	s->4	t->2	v->3	ä->2	
pa..	 ->1	(->1	
pa.1	8->1	
pa.D	e->15	
pa.E	f->1	n->1	t->1	
pa.F	r->2	ö->1	
pa.H	e->6	
pa.I	 ->2	
pa.J	a->8	
pa.K	o->1	
pa.M	a->1	e->1	å->1	
pa.N	ä->1	
pa.O	c->1	
pa.P	r->1	
pa.R	e->1	
pa.T	r->1	y->1	
pa.U	n->1	
pa.V	a->1	i->9	
pa.Ä	v->1	
pa; 	e->1	
pa?H	e->1	
pa?V	a->1	i->1	
paNä	s->1	
paci	t->5	
pack	n->5	
pad 	a->1	b->1	k->1	
pade	 ->13	m->2	s->9	
paga	n->3	
page	r->1	
pagn	e->1	
pagr	u->1	
pake	t->7	
pako	n->1	
pakt	 ->1	e->4	
pale	s->12	
pami	n->1	
pan 	e->1	o->1	
pan,	 ->1	
pand	e->64	
pane	l->1	
pani	e->7	v->1	
panj	 ->3	.->1	e->2	o->1	
pans	i->1	k->11	
pant	e->1	
papa	r->166	
papp	e->5	
par 	-->1	a->6	b->2	d->10	e->8	f->4	g->1	h->1	i->3	j->1	k->1	m->8	n->1	o->5	p->5	r->1	s->6	u->1	v->5	å->2	ö->2	
par.	A->1	D->1	I->1	
para	 ->4	b->1	d->6	g->2	l->5	m->2	r->3	t->3	
parc	o->1	
pare	 ->5	,->1	.->1	r->4	
pari	c->1	n->3	
park	 ->4	a->3	e->7	
parl	a->558	
parn	a->1	
pars	a->1	
part	 ->1	.->1	e->31	i->86	n->28	s->1	
parå	d->1	
pas 	-->2	a->60	b->4	c->1	d->4	e->5	f->18	g->3	h->2	i->12	j->10	k->8	l->3	m->9	n->6	o->9	p->10	r->2	s->15	t->2	u->1	v->13	å->1	
pas,	 ->5	
pas.	-->1	D->4	J->1	K->1	P->1	V->2	
pas:	 ->1	
pas?	S->1	
pass	 ->4	a->18	e->3	i->3	n->4	u->1	
past	 ->9	e->2	
pat 	-->1	d->1	e->3	f->1	m->1	n->2	s->4	t->1	
pat.	F->1	
pat:	 ->1	
pate	t->1	
pati	 ->4	e->5	o->1	s->3	
patj	ä->1	
patr	i->1	
pats	 ->8	.->1	
pava	l->3	
paya	n->2	
pbac	k->1	
pbri	n->3	
pbyg	g->20	
pbär	a->1	
pbåd	a->1	
pdat	e->3	
pdel	n->3	
pdra	g->22	
pe i	 ->1	
pe p	å->1	
pean	u->1	
peau	"->1	
peci	a->14	e->42	f->29	
peda	g->1	
pedi	t->1	
pedo	f->1	
pegl	a->11	i->1	
pegn	a->1	
pehå	l->13	
peis	e->2	k->710	
peka	 ->20	,->1	d->10	n->9	r->12	s->4	t->14	
pekt	 ->27	:->1	a->6	e->68	i->38	r->2	ö->6	
peku	l->4	
pel 	-->2	B->1	N->1	R->1	a->2	b->2	d->1	e->1	f->11	g->2	h->6	i->6	m->1	n->2	o->4	p->20	r->1	s->7	t->2	u->1	v->1	ä->2	
pel,	 ->7	
pel.	D->1	I->1	J->1	M->1	V->1	
pel:	 ->3	
pel;	 ->1	
pela	 ->14	?->1	d->1	r->24	s->1	t->5	
pele	n->1	t->1	
pell	 ->1	
peln	i->1	
pelp	l->1	
pelr	e->4	u->1	
pelv	i->28	
pen 	"->3	(->2	-->1	D->4	E->2	N->2	T->1	U->2	a->24	b->6	d->1	e->4	f->10	g->5	h->12	i->14	k->8	m->19	n->6	o->38	p->4	s->16	t->4	u->4	v->7	ä->16	å->3	
pen,	 ->26	
pen.	 ->1	.->1	D->6	E->1	H->3	J->7	K->1	M->2	N->3	P->1	S->3	T->2	V->1	Ä->1	
pen:	 ->2	
pen?	.->1	
penN	ä->1	
penb	a->36	
penc	e->1	
pend	e->5	i->1	
peng	a->55	
penh	a->2	e->60	
peni	n->1	
penn	d->1	i->10	
pens	 ->84	a->3	e->8	i->14	p->1	
pent	e->1	
penu	t->1	
per 	E->1	a->6	b->3	c->10	d->6	e->6	f->8	h->4	i->10	j->1	k->3	l->2	m->5	n->1	o->13	p->2	r->3	s->16	t->3	u->6	v->2	ä->5	å->3	
per,	 ->9	
per.	A->1	E->2	F->3	G->1	I->1	N->1	O->1	V->2	
per:	 ->2	
pera	 ->1	d->2	h->1	s->1	t->17	
pere	r->1	t->1	
perf	e->7	
peri	f->6	n->2	o->86	
perl	i->1	
perm	a->8	
pern	 ->1	a->49	
pero	n->1	
perr	o->1	
pers	 ->1	l->1	o->104	p->17	
pert	e->20	g->3	i->3	k->17	r->2	u->1	
pes 	e->1	r->1	
pesk	å->1	
pess	i->2	
pest	 ->1	e->4	
pet 	"->3	(->1	-->2	a->3	b->2	d->3	e->2	f->9	g->1	h->3	i->5	j->1	k->13	l->2	m->7	n->2	o->16	p->6	r->1	s->10	t->4	v->4	ä->1	ö->1	
pet)	 ->1	
pet,	 ->18	
pet.	H->1	J->1	M->2	N->1	O->1	P->1	
pet?	R->1	
pete	n->11	
peti	t->1	
pets	 ->15	.->1	f->1	
pfal	l->1	
pfan	n->1	
pfat	t->51	
pfyl	l->54	
pföd	n->1	
pföl	j->10	
pför	a->12	s->1	
pgic	k->3	
pgif	t->77	
pgod	k->1	
pgra	d->1	
pgå 	t->1	
pgåe	n->7	
pgån	g->2	
pgår	 ->5	
pgör	e->2	
phar	m->1	
pher	d->3	
phet	 ->2	,->1	s->1	
phov	 ->8	s->5	
phta	l->1	
phän	t->1	
phäv	a->3	s->2	
phål	 ->1	:->1	e->1	
phöj	s->1	
phör	 ->3	a->5	t->1	
pia 	t->1	
pic 	B->1	
pice	 ->1	
piel	l->8	
pien	 ->1	,->2	
pier	a->1	
pill	o->1	
pilo	t->4	
pin 	h->1	
pini	o->4	
pion	j->1	
pira	t->1	
pire	r->3	
pisk	a->2	
pit 	o->1	s->1	
pita	 ->6	,->1	.->3	l->17	
pite	l->6	
pitu	l->2	
pjak	t->1	
pkay	 ->3	,->3	.->1	D->1	b->1	s->2	
pkol	l->1	
pkom	m->6	
pkra	f->1	
pla 	s->1	
plac	e->17	
plad	e->1	
plan	 ->19	,->2	.->4	:->1	N->1	d->2	e->100	t->3	
plar	i->2	
plas	 ->2	t->6	
plat	s->44	t->1	
plem	e->11	
plen	 ->3	a->4	u->5	
plet	 ->3	t->14	
plev	a->7	d->1	e->4	s->2	t->3	
plex	 ->1	.->1	a->1	t->1	
plic	e->12	i->1	
plig	 ->18	,->2	.->1	a->44	h->4	t->35	
plik	t->33	
plim	a->3	e->1	s->1	
plin	 ->4	,->1	e->3	f->1	g->3	r->1	ä->4	
plit	t->4	
pliv	a->1	
plom	a->11	
plos	i->2	
plun	d->1	
plur	a->1	
plus	 ->2	
plys	a->2	n->2	
pläd	e->2	
plåd	e->11	
plåg	e->1	
plån	a->1	b->1	i->1	
plös	a->1	e->1	n->1	t->1	
plöt	s->4	
pman	a->51	i->7	
pmju	k->2	
pmun	t->21	
pmär	k->53	
pmät	t->2	
pmöt	e->12	
pna 	d->1	f->2	g->1	m->1	o->1	p->2	r->1	
pna,	 ->2	
pnad	e->3	
pnar	 ->2	e->1	
pnas	 ->2	
pnen	 ->2	
pnin	g->119	
pnå 	d->11	e->21	f->2	g->1	m->3	n->1	p->2	r->1	s->1	v->4	y->1	ö->1	
pnå,	 ->1	
pnå.	 ->1	F->1	J->1	S->1	
pnåd	d->6	
pnår	 ->13	
pnås	 ->5	.->2	
pnåt	t->13	
po, 	s->1	
poet	 ->1	
pok 	i->1	
pok,	 ->1	
poke	n->2	
pol 	a->2	i->2	m->2	o->6	s->2	t->1	
pol,	 ->3	
pol-	f->1	
pol.	E->1	H->1	
pol;	 ->1	
pola	v->1	
pole	 ->1	m->1	
polf	r->1	ö->2	
poli	c->4	n->1	s->18	t->534	
polk	o->1	
pols	 ->3	i->1	
pond	e->1	
pone	n->5	r->7	
pons	 ->1	r->1	
pont	a->4	
pool	,->1	
popu	l->7	
por,	 ->1	
pord	f->1	
porn	o->2	
pors	l->1	
port	 ->83	)->1	,->9	-->3	.->3	N->1	a->1	b->2	d->1	e->109	f->3	g->1	i->9	k->2	m->2	n->1	o->3	p->1	s->8	u->73	v->1	
porä	r->2	
pos 	b->1	
posi	t->87	
post	 ->7	.->1	e->6	v->1	
pote	n->6	s->1	t->1	
poti	s->5	
pots	 ->1	
poul	o->5	
poän	g->12	
pp (	k->2	
pp -	 ->2	
pp E	u->1	
pp T	i->1	
pp a	l->5	n->5	t->3	v->11	
pp b	e->2	i->1	å->1	
pp d	e->40	o->1	ä->1	
pp e	f->3	l->1	n->10	t->6	x->1	
pp f	o->1	r->11	u->1	ö->12	
pp g	e->2	r->1	
pp h	a->6	e->1	u->1	ä->3	ö->1	
pp i	 ->22	d->1	g->4	n->3	
pp k	a->1	o->6	
pp l	a->1	i->1	ä->3	
pp m	e->8	å->1	
pp n	a->1	y->1	å->3	
pp o	c->6	l->1	m->2	r->2	
pp p	o->1	r->3	å->12	
pp r	e->2	ä->3	ö->1	
pp s	a->1	i->2	k->3	o->7	t->2	ä->2	å->1	
pp t	i->11	o->1	r->1	v->1	y->2	
pp u	n->2	t->7	
pp v	a->3	i->2	ä->2	
pp ä	n->2	r->7	
pp, 	E->1	a->2	b->1	d->1	e->4	f->1	h->2	i->1	j->1	m->2	n->1	o->2	r->1	s->3	v->1	
pp..	(->1	
pp.A	h->1	
pp.D	e->5	
pp.F	a->1	
pp.J	a->7	
pp.M	e->1	
pp.P	å->1	
pp.V	i->3	
pp.Ä	n->1	v->1	
pp?H	u->1	
ppa 	a->1	e->2	i->6	m->1	r->1	s->1	t->4	ö->1	
ppad	e->8	
ppan	d->2	
ppar	 ->3	a->1	
ppas	 ->96	,->4	t->9	
ppba	c->1	
ppbr	i->3	
ppby	g->20	
ppbä	r->1	
ppbå	d->1	
ppda	t->3	
ppde	l->3	
ppdr	a->22	
ppe 	i->1	
ppeh	å->13	
ppel	l->1	
ppen	 ->61	,->4	.->4	b->36	h->60	s->13	
pper	 ->32	,->4	.->5	:->1	a->1	e->1	i->2	l->1	n->21	s->2	
ppet	 ->32	,->2	.->1	
ppfa	n->1	t->51	
ppfy	l->54	
ppfö	d->1	l->10	r->13	
ppgi	c->3	f->77	
ppgr	a->1	
ppgå	 ->1	n->2	r->5	
ppgö	r->2	
pphe	t->4	
ppho	v->13	
pphä	n->1	v->5	
pphö	j->1	r->9	
ppja	k->1	
ppko	l->1	m->6	
ppla	 ->1	d->1	n->2	s->2	
pple	v->17	
ppli	n->2	v->1	
pply	s->4	
pplå	d->11	
pplö	s->4	
ppma	n->58	
ppmj	u->2	
ppmu	n->21	
ppmä	r->53	t->2	
ppmö	t->12	
ppna	 ->8	,->2	d->1	r->3	s->2	
ppni	n->17	
ppnå	 ->49	,->1	.->4	d->6	r->13	s->7	t->13	
ppon	e->3	
ppor	d->1	t->114	
ppos	i->2	
ppre	n->2	p->52	
ppri	k->6	
ppro	p->5	
ppru	s->1	
ppry	c->1	
pprä	c->2	k->1	t->36	
pprö	r->5	
pps 	u->1	v->3	
ppsa	m->4	t->3	
ppsb	r->1	y->1	
ppsk	a->23	j->4	o->2	
ppsp	å->2	
ppsr	e->2	ä->1	
ppss	t->1	ä->2	
ppst	o->4	ä->3	å->32	
ppsv	a->2	
ppsä	g->1	t->2	
ppt 	e->2	i->1	s->1	t->1	
ppta	g->7	r->1	s->2	
ppte	 ->1	s->2	
ppti	l->1	
ppto	g->2	
pptr	ä->10	
pptä	c->11	
ppun	d->1	
ppve	r->2	
ppvi	g->1	s->5	
ppvä	g->1	r->1	
ppy 	e->1	
prac	k->1	
prag	m->1	
prak	t->33	
pran	a->1	
prat	.->1	a->4	
prax	i->8	
prec	i->43	
pref	e->3	
prej	u->4	
prel	i->3	
prem	i->10	
pren	s->2	ö->3	
prep	a->51	n->1	
prer	o->1	
pres	e->47	i->9	s->21	t->4	
pric	k->3	
prid	a->4	e->5	i->1	n->8	s->2	
prik	t->6	
pril	 ->2	.->1	
prim	i->1	
prin	c->194	i->1	
prio	r->38	
pris	 ->4	.->1	a->1	e->19	n->1	s->1	u->1	
priv	a->21	i->7	
prob	l->174	
proc	e->201	
prod	u->76	
prof	e->7	i->3	
prog	r->238	
proj	e->62	
prok	l->1	
prom	i->22	
pron	a->1	
prop	 ->3	,->1	.->1	a->4	o->9	å->1	
pros	t->1	
prot	e->13	o->24	
prov	 ->9	i->5	k->1	s->3	
prun	g->19	
prus	t->1	
pryc	k->1	
präc	k->2	
präg	l->5	
präk	n->1	
prän	t->1	
prät	t->36	
pråk	 ->5	.->1	a->9	e->3	l->3	o->2	t->1	
prån	g->2	
prör	a->3	d->2	
pröv	a->9	n->5	o->1	
ps a	v->1	
ps f	a->1	
ps u	t->1	
ps v	ä->3	
ps- 	o->1	
ps.J	u->1	
ps.M	e->1	
psam	l->4	
psat	t->3	
psav	t->2	
psbe	f->1	g->1	s->2	
psbr	o->1	
psby	g->1	
psdi	r->1	
psfr	å->1	
psin	i->7	n->1	s->6	t->1	
psis	 ->1	
pska	t->23	
pskh	e->1	
pskj	u->4	
psko	n->3	v->2	
pskä	l->2	
psla	g->5	
psma	s->2	
psme	d->1	
psmä	n->16	
psmå	l->1	
psni	v->11	
pson	 ->1	
psor	g->1	
pspe	l->2	
pspo	l->2	
pspr	o->3	
pspå	r->2	
psra	m->1	
psre	d->2	g->9	
psrä	t->9	
psst	r->1	ä->1	ö->2	
pssy	s->1	
pssä	t->2	
psto	d->4	
pstä	l->3	
pstå	 ->3	:->1	n->1	r->16	t->11	
psva	r->2	
psyk	o->1	
psäg	n->1	
psät	t->2	
psåt	g->2	
pt b	e->2	
pt d	e->1	i->1	
pt e	n->1	t->1	
pt f	o->1	
pt i	 ->2	n->1	
pt k	o->1	
pt o	r->1	
pt s	e->1	k->1	
pt t	i->1	r->1	
pt u	t->5	
pt v	a->1	
pt ö	v->1	
pt.D	e->1	
pt.H	a->1	
pta 	k->1	v->1	
pta.	D->1	
ptab	e->27	l->10	
ptag	a->3	e->2	n->2	
ptan	s->7	
ptar	 ->1	
ptas	 ->1	.->1	
pte 	d->1	f->1	l->1	t->1	u->2	
ptem	b->15	
pten	 ->3	,->1	
pter	a->45	
ptes	 ->2	
ptet	 ->3	
ptik	e->3	
ptil	l->1	
ptim	a->3	i->4	
ptio	n->14	
ptis	k->5	
ptog	a->2	s->2	
ptom	 ->1	
pträ	d->9	t->1	
ptäc	k->11	
publ	i->26	
pula	r->1	
puli	s->4	
puls	 ->2	e->4	
pulä	r->2	
pump	a->2	
pund	 ->2	.->1	a->1	
punk	t->342	
puri	t->1	
pus 	j->5	
pver	k->2	
pvig	l->1	
pvil	l->1	
pvis	.->1	a->4	
pväg	a->1	
pvär	d->1	
py e	n->1	
pyra	m->1	
pyri	g->1	
pänn	a->4	i->7	
pärr	 ->1	a->2	
på -	 ->5	
på 1	0->1	3->2	4->1	
på 2	0->3	2->1	
på 3	3->1	4->1	7->1	
på 4	0->1	
på 5	 ->1	0->2	
på 7	,->1	5->1	
på 8	0->2	6->1	
på 9	0->1	5->1	
på A	l->2	t->1	
på B	S->1	a->5	e->1	
på C	E->1	S->1	
på E	G->3	U->4	r->1	u->10	
på F	ö->1	
på G	e->1	o->1	
på H	o->1	
på I	S->1	n->6	r->1	s->1	
på M	a->1	
på O	l->1	
på P	a->1	
på R	i->2	o->1	
på T	y->1	
på V	ä->2	
på a	c->1	k->1	l->29	n->16	r->11	s->1	t->145	v->1	
på b	a->4	e->8	i->5	l->1	o->3	r->7	ä->9	å->3	
på c	e->1	i->1	r->1	
på d	a->8	e->292	i->2	j->7	u->4	y->1	
på e	f->2	g->3	k->2	l->1	m->1	n->55	r->5	t->142	u->12	x->1	
på f	a->3	e->4	i->2	l->3	r->12	y->2	ä->6	ö->64	
på g	a->1	e->16	l->1	o->2	r->79	ä->1	å->5	ö->1	
på h	a->5	e->1	j->1	u->14	ä->1	ö->1	
på i	 ->4	c->1	l->1	n->19	t->1	
på j	a->1	o->1	u->2	ä->3	
på k	a->5	l->2	n->1	o->37	r->1	u->1	v->1	ä->1	ö->1	
på l	a->12	i->3	o->3	ä->6	å->9	ö->1	
på m	a->12	e->19	i->28	o->6	y->2	ä->1	å->5	ö->4	
på n	a->4	e->1	o->4	y->26	ä->8	å->21	
på o	b->2	c->4	l->4	m->19	n->2	r->2	s->5	
på p	a->1	e->3	l->9	o->1	r->9	
på r	a->2	e->26	i->2	y->1	ä->11	å->7	
på s	a->22	e->11	i->31	j->1	k->6	l->1	m->1	n->1	o->1	p->10	t->13	u->2	v->1	y->4	ä->5	å->16	
på t	a->7	e->4	i->10	j->1	o->10	r->10	v->7	ä->1	
på u	n->8	p->3	t->5	
på v	a->16	e->8	i->16	ä->34	å->16	
på y	t->1	
på z	i->1	
på Ö	s->2	
på ä	n->6	r->3	
på å	h->1	r->1	t->5	
på ö	k->1	n->1	p->5	v->1	
på, 	e->2	f->1	h->1	l->1	m->3	n->1	o->5	v->1	ä->1	
på.B	e->1	
på.D	e->3	o->1	
på.E	n->1	u->1	
på.J	a->3	
på.N	o->1	
på.O	r->1	
på.U	n->1	
på.V	i->1	
på.Ä	r->2	
på: 	f->2	Ö->1	
på?.	 ->1	
på?J	a->1	
påbj	u->1	
påbö	r->11	
pådr	a->1	
påfr	e->1	
påfö	l->4	
pågi	c->3	
pågå	 ->1	e->6	r->10	t->1	
påla	g->1	
påle	n->1	
påli	t->1	
pålä	g->1	
påmi	n->30	
påpe	k->50	
pår 	a->1	h->1	i->1	t->1	
pår,	 ->2	
påra	 ->2	n->1	s->1	
påre	n->1	
pårn	i->2	
påsk	y->7	
påst	r->1	å->20	
påta	g->4	l->5	
påtr	y->3	
påtv	i->4	
påve	r->37	
påvi	s->3	
pé o	c->1	
péer	 ->4	,->2	n->3	
péry	s->1	
pöke	 ->1	.->1	n->1	
pöks	t->1	
qal 	f->1	ä->1	
qua 	n->2	
qual	 ->6	"->1	,->1	
que 	k->1	
que,	 ->1	
ques	 ->4	"->1	
quie	r->1	
quin	s->1	
quio	l->1	
quis	i->1	
quit	a->1	
quo 	s->1	
quo,	 ->1	
quqa	l->2	
r "K	u->1	
r "a	n->2	
r "f	o->1	
r "i	n->1	
r "k	r->1	
r "n	a->1	
r "ö	v->1	
r (C	5->4	
r (F	I->1	
r (a	r->1	
r (i	 ->1	
r - 	1->2	a->11	c->1	d->12	e->5	f->2	g->1	h->3	i->8	j->1	k->4	l->1	m->2	n->2	o->9	s->10	t->1	u->1	v->3	ä->6	ö->1	
r -,	 ->1	
r 1 	4->1	f->1	
r 1,	2->1	4->1	
r 1/	3->1	
r 10	 ->3	0->1	
r 12	 ->1	4->1	
r 13	0->1	
r 15	 ->2	
r 16	7->1	
r 17	4->1	6->2	
r 19	2->1	3->1	7->1	8->2	9->67	
r 2 	b->1	
r 20	 ->4	0->58	1->2	
r 25	 ->1	
r 26	2->1	
r 27	 ->2	
r 28	 ->1	
r 29	 ->3	
r 3 	0->1	
r 3-	4->1	
r 30	 ->2	
r 31	 ->1	
r 32	 ->1	.->1	
r 33	 ->2	2->1	
r 35	 ->2	
r 36	 ->1	
r 37	 ->1	
r 38	 ->1	
r 39	 ->1	
r 4 	0->1	
r 40	 ->4	
r 41	 ->1	
r 42	 ->1	
r 43	.->1	
r 44	 ->1	
r 45	 ->1	
r 46	 ->1	
r 5 	f->1	m->1	å->1	
r 5,	8->1	
r 50	 ->2	
r 6 	f->1	
r 60	 ->1	
r 7 	g->1	p->1	
r 7.	F->1	
r 73	,->1	
r 75	 ->1	
r 76	 ->1	
r 8 	f->1	
r 80	 ->4	
r 81	 ->1	
r 9 	f->1	
r 90	 ->2	
r 97	.->1	/->1	
r Ag	r->1	
r Al	a->1	b->1	s->1	t->5	
r Am	o->2	
r An	t->1	
r Ar	a->1	
r Az	o->1	
r BN	I->1	P->1	
r BS	E->1	
r Ba	r->13	
r Be	l->1	r->5	
r Bi	s->1	
r Bo	l->1	u->2	w->2	
r Br	e->3	o->2	y->1	
r CE	N->1	
r CS	U->1	
r Ce	n->2	
r Co	c->1	n->1	x->3	
r Da	n->3	
r De	u->1	
r Do	r->1	
r Du	h->1	
r EC	H->1	
r EG	-->5	.->1	:->1	
r EM	U->2	
r EU	 ->2	,->1	-->4	.->2	:->9	
r Eg	y->1	
r Eh	u->1	
r Ek	o->1	
r El	s->1	
r Er	i->3	
r Eu	r->112	
r Ev	a->3	
r Ex	x->1	
r FN	.->1	:->2	
r FP	Ö->2	
r Fa	r->1	
r Fi	n->1	
r Fl	o->1	
r Fo	U->1	l->1	
r Fr	a->1	u->1	
r Fö	r->6	
r GA	S->1	
r Ga	m->2	
r Ge	n->1	
r Go	l->3	m->1	
r Gr	a->1	e->1	
r Gu	s->1	t->1	
r Ha	i->1	
r He	l->1	
r Hi	m->1	
r Hä	n->2	
r I 	o->1	
r I-	p->1	
r II	 ->1	-->2	I->1	
r IM	O->1	
r IN	T->1	
r In	t->2	
r Is	r->5	
r It	a->1	
r Ja	p->1	
r Jo	n->2	s->1	
r Jö	r->2	
r Ka	n->3	
r Ki	n->11	
r Ko	c->1	s->1	u->1	
r Ku	l->2	m->1	
r Kv	i->1	
r Ky	o->1	
r La	a->7	n->3	
r Le	i->1	
r Li	s->1	
r Lo	t->2	
r Lu	x->1	
r Ly	n->2	
r Ma	a->2	r->2	
r Me	l->1	
r Mo	n->16	r->1	
r Na	t->1	
r Ne	d->1	
r Ni	e->1	k->2	
r No	g->1	
r OF	S->1	
r OL	A->2	
r Or	a->1	
r Os	l->1	
r PP	E->1	
r PV	C->1	
r Pa	c->1	l->3	p->1	t->18	
r Po	e->3	h->1	m->1	n->1	o->1	r->3	
r Pr	e->1	o->1	
r RE	P->1	
r Ra	p->1	s->1	
r Re	d->2	
r Rh	ô->1	
r Ro	t->1	
r Ru	s->1	
r Rå	d->1	
r Sa	v->2	
r Sc	h->6	
r Se	a->1	g->2	i->2	
r Sh	a->1	
r Sk	o->1	
r So	l->2	
r Sp	e->1	
r Sw	o->1	
r Sy	r->2	
r Sã	o->1	
r Ta	c->1	m->1	n->1	
r Te	s->1	
r Th	e->1	
r Ti	b->6	
r To	r->1	
r Ts	a->2	
r Tu	r->4	
r UC	L->1	
r UN	M->1	
r US	A->1	D->1	
r Ur	q->1	
r Vi	t->5	
r Vo	l->1	
r WT	O->1	
r Wa	l->3	s->1	
r Wy	n->1	
r [S	E->1	
r ab	s->14	
r ac	c->6	
r ad	m->1	
r ag	e->1	
r ai	d->1	
r ak	t->12	
r al	d->9	l->282	
r am	b->3	e->1	
r an	a->8	b->1	d->25	f->2	g->9	h->1	k->1	l->5	m->3	n->13	o->3	s->85	t->22	v->18	
r ar	b->35	r->1	t->7	
r as	"->1	y->4	
r at	t->1979	
r au	c->1	
r av	 ->177	.->1	b->2	d->1	f->4	g->14	h->1	i->2	l->2	s->41	t->2	u->1	v->4	
r ba	k->8	l->1	n->2	r->30	s->3	
r be	a->5	d->13	f->17	g->24	h->32	k->16	l->2	m->1	r->48	s->41	t->57	v->13	
r bi	d->11	f->1	l->28	n->1	s->6	
r bj	u->1	
r bl	.->2	a->6	i->31	o->2	y->2	
r bo	m->3	r->10	s->3	t->1	v->1	
r br	a->21	e->1	i->15	o->7	u->2	y->1	å->4	ö->2	
r bu	d->21	s->1	
r by	g->6	r->2	x->1	
r bä	r->1	s->3	t->12	
r bå	d->11	
r bö	j->1	r->29	
r ca	p->10	
r ce	n->4	
r ch	o->2	
r ci	r->3	t->2	v->3	
r co	p->1	r->1	
r da	g->15	n->2	t->1	
r de	 ->396	,->2	b->32	c->3	f->5	l->38	m->58	n->471	r->27	s->111	t->1069	
r di	a->1	p->1	r->12	s->25	t->2	v->1	
r dj	u->9	ä->1	
r do	c->33	k->2	l->6	m->7	
r dr	a->13	i->2	o->1	
r du	 ->2	b->2	g->1	m->1	
r dy	k->1	n->1	
r dä	r->105	
r då	 ->22	l->7	
r dö	d->3	l->2	r->2	t->1	
r ec	u->2	
r ed	 ->1	
r ef	f->12	t->34	
r eg	e->16	n->1	o->1	
r ej	 ->5	,->1	.->2	
r ek	o->28	
r el	e->2	l->59	v->1	
r em	e->28	o->9	
r en	 ->587	.->1	a->2	b->4	d->12	e->15	g->3	h->9	i->2	k->5	l->20	o->6	s->9	
r er	 ->34	,->10	.->4	a->7	f->2	h->2	i->2	k->4	s->2	t->9	
r et	a->4	n->1	t->308	
r eu	r->31	
r ev	i->3	
r ex	a->2	c->1	e->7	i->1	p->7	t->9	
r fa	c->1	k->15	l->22	m->1	n->1	r->19	s->15	t->7	
r fe	d->1	l->10	m->5	
r fi	c->2	n->33	s->7	
r fj	o->1	
r fl	a->1	e->17	i->1	o->2	y->7	ä->1	
r fo	d->3	l->7	n->1	r->49	
r fr	a->99	e->10	i->17	u->1	ä->14	å->155	
r fu	l->17	n->9	
r fy	l->1	r->2	s->1	
r fä	r->1	s->1	
r få	 ->10	,->2	.->1	r->12	t->28	
r fö	g->1	l->14	r->745	
r ga	g->3	m->1	n->7	r->4	
r ge	 ->2	m->30	n->62	r->2	s->2	t->12	
r gi	l->1	v->14	
r gj	o->49	
r gl	a->12	o->1	ä->2	ö->4	
r go	d->27	l->1	t->1	
r gr	a->11	i->1	u->37	ä->13	å->1	
r gu	d->2	
r gy	n->3	
r gä	l->5	r->3	
r gå	 ->1	n->4	r->12	t->11	
r gö	m->2	r->25	
r ha	 ->15	d->1	f->16	k->1	l->6	m->3	n->62	r->112	v->2	
r he	d->2	l->104	m->5	n->10	r->1	t->1	
r hi	n->2	s->5	t->12	
r hj	ä->10	
r ho	m->2	n->15	p->1	r->1	s->7	t->6	
r hu	m->1	n->2	r->36	v->12	
r hy	s->2	
r hä	l->3	m->1	n->17	r->30	s->1	v->3	
r hå	l->12	r->2	
r hö	g->12	j->1	r->15	
r i 	-->1	2->1	A->1	B->4	C->1	D->2	E->41	F->4	I->3	K->7	L->1	M->1	O->1	P->1	S->5	T->1	U->2	W->1	a->28	b->10	d->121	e->30	f->45	g->12	h->8	i->3	j->2	k->22	l->2	m->23	n->6	o->13	p->25	r->14	s->52	t->7	u->13	v->24	Ö->7	ä->1	å->1	ö->5	
r i.	A->1	
r ia	n->1	
r ib	l->3	
r ic	k->2	
r id	e->5	é->2	
r if	r->6	
r ig	e->12	n->1	
r ih	o->4	
r ik	r->1	
r il	l->4	
r im	m->1	
r in	 ->11	b->3	c->2	d->14	f->37	g->59	i->6	k->5	l->10	n->21	o->56	r->15	s->22	t->443	v->13	
r ir	l->1	
r is	c->1	r->1	
r it	u->6	
r iv	ä->1	
r ja	,->1	g->284	
r jo	r->17	
r ju	 ->34	,->2	d->1	l->1	r->5	s->16	
r jä	m->5	r->3	
r ka	l->5	m->8	n->60	p->1	r->3	t->12	
r ke	m->1	
r kl	a->28	i->2	o->5	y->1	
r kn	a->5	u->3	
r ko	a->1	l->9	m->332	n->98	r->14	s->14	
r kr	a->14	e->1	i->12	y->1	ä->11	
r ku	b->1	l->27	n->16	r->1	s->3	
r kv	a->6	e->2	i->10	ä->2	
r kä	m->2	n->13	r->8	
r kö	l->1	r->2	
r la	g->53	n->7	s->3	
r le	 ->1	d->32	g->6	t->7	v->3	
r li	d->3	g->7	k->29	s->2	t->19	v->22	
r lo	b->1	g->2	k->4	t->1	v->5	
r lu	f->1	g->2	r->1	
r ly	c->17	f->1	s->5	
r lä	c->1	g->11	k->1	m->20	n->22	r->1	s->4	t->9	
r lå	n->32	s->1	t->4	
r lö	j->2	n->5	p->4	s->4	
r ma	i->3	j->4	k->1	l->2	n->175	r->9	s->2	t->4	
r me	d->293	k->1	l->18	n->21	r->31	s->3	t->4	
r mi	g->99	l->46	n->66	s->5	t->10	
r mo	b->1	d->5	g->1	n->1	r->7	t->39	
r mu	n->1	t->1	
r my	c->104	n->5	
r mä	n->32	
r må	l->9	n->40	r->1	s->45	
r mö	j->44	t->2	
r na	k->1	m->1	r->1	t->44	
r ne	d->6	g->2	j->3	k->1	r->4	
r ni	 ->51	,->3	v->2	
r no	g->3	r->10	t->7	
r nu	 ->40	,->2	.->2	:->1	m->1	
r ny	 ->3	a->16	c->1	h->1	l->2	t->4	
r nä	m->13	r->85	s->12	
r nå	g->106	t->4	
r nö	d->38	j->7	
r oa	c->7	v->2	
r ob	a->1	e->5	s->1	
r oc	h->570	k->162	
r oe	n->2	r->6	t->1	
r of	f->9	r->1	t->23	u->2	ö->4	
r oj	ä->1	
r ok	l->3	u->1	
r ol	a->1	i->9	j->4	y->4	ö->1	
r om	 ->253	,->5	.->6	b->1	f->11	k->9	l->1	p->1	r->13	s->2	v->1	ö->3	
r on	ö->2	
r op	i->1	
r or	d->28	i->1	o->13	s->5	ä->4	
r os	s->132	t->1	ä->1	å->1	
r ot	i->3	r->1	å->1	
r ou	m->1	n->2	t->2	
r ov	a->1	ä->1	
r oö	v->1	
r pa	p->1	r->58	s->3	
r pe	k->3	n->11	r->33	s->1	
r pl	a->10	e->2	i->2	u->1	
r po	l->23	s->9	t->1	ä->1	
r pr	a->3	e->16	i->10	o->56	ä->1	ö->2	
r pu	n->10	
r på	 ->302	,->3	.->3	b->4	f->1	l->1	m->2	p->7	s->1	t->4	v->6	
r ra	d->2	k->2	m->1	p->4	s->3	t->5	
r re	a->6	c->1	d->35	f->13	g->71	h->1	j->2	k->7	l->6	n->4	p->4	s->23	t->2	v->4	
r ri	g->1	k->11	m->4	n->1	s->13	
r ro	l->5	p->1	s->2	
r ru	i->1	m->2	n->1	s->1	t->1	
r ry	c->1	
r rä	d->4	k->7	t->66	
r rå	d->50	
r rö	r->11	s->15	
r sa	d->2	g->20	k->9	m->75	n->9	t->6	
r se	 ->8	d->29	g->3	k->4	n->14	r->6	s->1	t->9	x->4	
r si	d->2	g->126	k->1	n->58	s->5	t->26	
r sj	u->3	ä->29	ö->1	
r sk	a->84	e->6	i->9	j->5	o->5	r->14	u->24	y->18	ä->5	ö->2	
r sl	a->3	u->13	ä->3	
r sm	u->1	å->8	
r sn	a->12	e->2	ä->1	
r so	c->4	l->3	m->636	v->1	
r sp	a->3	e->18	i->1	o->1	r->4	ä->2	å->1	
r st	a->44	e->4	i->2	o->56	r->24	u->3	y->4	ä->13	å->22	ö->38	
r su	b->5	n->1	
r sv	a->11	å->19	
r sy	d->1	f->4	m->4	n->8	s->26	
r sä	g->4	k->48	l->1	m->1	n->1	r->37	t->3	
r så	 ->61	,->3	d->10	l->19	s->4	v->7	
r sö	d->1	n->3	
r t.	e->3	
r ta	 ->9	c->1	g->26	l->338	n->4	r->2	s->2	
r te	k->6	m->2	n->1	x->2	
r ti	b->2	d->18	l->413	o->4	t->2	
r tj	u->1	ä->14	
r to	b->1	g->2	l->5	n->2	p->1	r->3	t->3	
r tr	a->26	e->15	o->15	y->3	ä->8	å->2	ö->1	
r tu	n->2	r->3	s->2	
r tv	e->3	i->8	u->5	ä->3	å->21	
r ty	c->1	d->15	n->2	p->11	v->7	
r tä	n->6	r->1	t->1	
r tå	g->1	
r un	d->67	g->9	i->45	
r up	p->129	
r ur	 ->7	s->2	v->1	
r ut	 ->24	,->3	.->3	?->1	a->51	b->8	e->8	f->20	g->8	i->4	k->2	l->2	m->2	n->4	o->3	p->1	r->8	s->37	t->11	v->43	ö->7	
r va	d->36	g->1	k->5	l->10	n->5	r->116	t->2	
r ve	c->2	d->1	k->1	l->1	m->1	r->46	t->23	
r vi	 ->426	,->5	d->31	g->1	k->64	l->50	n->1	r->1	s->44	t->9	
r vo	l->1	n->1	t->1	
r vu	n->2	x->1	
r vä	c->5	g->5	l->39	n->7	r->15	s->4	x->2	
r vå	l->1	r->89	
r yn	g->1	
r yp	p->1	
r yr	k->2	
r yt	t->16	
r ÖV	P->1	
r Ös	t->7	
r äg	n->5	t->3	
r äl	d->4	
r äm	n->3	
r än	 ->59	d->38	g->1	n->17	
r är	 ->145	a->2	e->1	l->2	
r äv	e->35	
r å 	a->1	e->1	
r åk	l->1	
r ål	a->1	
r år	 ->27	,->1	e->7	t->1	
r ås	a->1	i->3	k->1	t->1	
r åt	 ->8	a->4	e->33	f->1	g->6	m->3	s->2	t->2	
r öa	r->1	
r öd	e->1	
r ög	o->7	
r ök	a->13	
r ön	s->7	
r öp	p->16	
r ör	e->2	
r ös	t->3	
r öv	a->1	e->92	r->29	
r! 1	9->1	
r! A	v->1	
r! B	e->1	l->1	
r! C	e->1	
r! D	e->19	i->1	
r! E	f->4	r->1	t->1	u->4	
r! F	ö->8	
r! G	o->1	r->1	
r! H	i->1	
r! I	 ->9	
r! J	a->25	ä->1	
r! K	a->1	
r! L	å->4	
r! M	e->1	
r! N	i->1	ä->2	å->1	
r! O	m->1	
r! P	P->1	å->1	
r! S	o->3	
r! T	a->2	i->3	
r! U	n->2	
r! V	i->10	å->1	
r! Ä	v->3	
r! Å	r->1	
r!"D	e->1	
r!"O	m->1	
r!.H	e->1	
r!De	 ->3	t->4	
r!Ef	t->1	
r!Er	i->1	
r!Ja	g->5	
r!Me	d->1	
r!Mi	n->1	
r!My	c->1	
r!Ti	l->1	
r!Vi	 ->2	
r" h	a->1	
r" m	å->2	
r" o	c->1	
r" s	o->2	
r"),	 ->1	
r", 	s->1	
r".D	e->1	
r".J	a->1	
r".O	m->1	
r) B	o->1	
r) V	i->1	
r) o	c->3	
r).)	B->1	
r)? 	H->1	
r)Fr	u->2	
r)Ja	g->1	
r)Ko	n->1	
r)Ta	c->1	
r, "	n->1	
r, (	B->1	
r, 1	6->1	
r, B	u->1	
r, E	u->1	
r, G	a->1	
r, M	a->1	
r, P	a->1	
r, T	h->1	y->1	
r, W	a->1	
r, a	c->1	d->1	l->9	n->6	r->1	t->37	v->5	
r, b	a->1	e->5	i->1	l->6	o->1	r->1	ä->3	å->3	
r, d	e->19	i->1	j->1	v->8	ä->11	å->7	ö->1	
r, e	f->10	l->5	n->17	r->1	t->3	x->2	
r, f	i->2	o->1	r->16	å->1	ö->36	
r, g	a->1	e->7	y->1	å->1	ö->2	
r, h	a->10	e->18	o->1	u->2	ä->2	ö->1	
r, i	 ->19	b->1	c->1	n->29	
r, j	a->10	ä->2	
r, k	a->7	o->19	r->4	u->1	ä->18	
r, l	a->1	e->2	i->8	o->1	ä->2	å->2	
r, m	a->3	e->75	i->10	o->2	y->2	ä->5	å->6	
r, n	a->1	e->2	i->2	o->1	y->2	ä->11	å->6	
r, o	a->1	c->111	l->1	m->17	r->4	
r, p	e->1	l->1	r->5	å->7	
r, r	e->3	o->1	ä->3	å->1	ö->1	
r, s	a->8	e->1	i->2	j->1	k->5	m->1	n->3	o->69	p->1	t->3	v->2	ä->7	å->20	
r, t	a->2	i->17	j->3	r->6	u->1	y->2	
r, u	n->10	p->4	t->29	
r, v	a->6	e->3	i->32	ä->4	å->1	
r, ä	n->3	r->26	v->8	
r, å	t->7	
r, ö	v->1	
r- o	c->4	
r- s	o->1	
r-bi	l->1	
r-ko	m->1	
r-na	t->1	
r-pr	o->11	
r-re	g->1	
r. (	F->1	
r. A	l->1	
r. D	e->7	
r. E	f->1	n->3	u->1	
r. F	r->1	
r. H	e->1	
r. J	a->2	
r. M	a->1	e->2	
r. N	i->1	
r. S	y->1	å->1	
r. T	i->1	
r. V	i->1	å->1	
r. i	n->1	
r. Ä	n->1	
r.(A	p->1	
r.(I	T->1	
r.(L	i->1	
r.) 	H->1	
r.)S	ä->1	
r.- 	(->3	H->1	
r.. 	(->4	
r..(	E->2	N->1	
r...	(->1	H->1	
r..H	e->1	
r..V	i->1	
r.90	 ->1	
r.Al	l->3	t->1	
r.Am	e->1	
r.An	t->1	
r.At	t->4	
r.Av	 ->4	
r.Ba	r->2	
r.Be	d->2	f->1	t->4	
r.Bl	a->2	
r.Bo	s->1	
r.Br	e->1	
r.CS	U->1	
r.Da	g->1	
r.De	 ->31	n->42	s->8	t->145	
r.Di	r->1	
r.Do	m->1	
r.Dä	r->14	
r.Då	 ->2	
r.EU	-->2	
r.Ef	t->5	
r.En	 ->10	b->1	l->3	
r.Er	f->1	
r.Et	t->6	
r.Eu	r->7	
r.Ex	e->1	
r.FP	Ö->1	
r.Fe	m->1	
r.Fo	l->1	
r.Fr	a->1	e->1	i->1	u->7	å->3	
r.Få	r->1	
r.Fö	r->43	
r.Ge	m->2	n->5	
r.Gö	r->1	
r.Ha	n->1	
r.He	r->25	
r.Hu	r->2	v->1	
r.Hä	n->2	r->6	
r.I 	E->1	H->1	I->3	R->1	a->2	b->1	d->6	e->3	f->1	g->1	j->1	m->1	r->3	s->2	v->3	
r.In	d->1	g->3	o->3	r->1	t->1	
r.It	a->1	
r.Ja	c->1	g->118	
r.Ka	n->2	r->1	
r.Ki	n->1	
r.Ko	d->1	m->21	n->5	
r.Kr	a->1	
r.Kv	i->1	
r.Kä	r->1	
r.La	n->1	
r.Li	k->3	
r.Ly	c->1	
r.Lå	t->6	
r.Ma	n->5	r->1	
r.Me	d->7	l->1	n->20	r->1	
r.Mi	n->4	
r.My	l->1	
r.Mä	n->1	
r.Na	t->4	
r.Ni	 ->1	v->1	
r.Nu	 ->1	
r.Ny	a->1	
r.Nä	r->10	
r.Nå	g->1	
r.Ob	e->1	
r.Oc	h->7	k->1	
r.Om	 ->16	r->1	
r.Or	d->1	o->1	
r.Pa	r->2	
r.Pl	a->1	
r.Pr	o->3	
r.Pu	n->1	
r.På	 ->3	
r.Ra	s->1	
r.Re	d->1	f->1	n->1	v->2	
r.Ri	s->1	
r.Rä	k->1	
r.Rå	d->3	
r.Sa	m->5	
r.Se	d->2	
r.Sk	u->1	
r.Sl	u->2	
r.So	m->7	
r.St	a->1	o->1	r->1	ö->2	
r.Så	 ->2	d->1	l->2	
r.Ta	c->5	
r.Te	r->1	
r.Ti	l->15	
r.Tr	o->1	
r.Ty	 ->1	v->2	
r.Un	d->6	i->1	
r.Ut	e->1	
r.Va	d->8	l->1	r->5	
r.Ve	m->2	
r.Vi	 ->85	d->1	s->2	
r.Vå	r->5	
r.ko	m->1	
r.Än	d->5	
r.Är	 ->3	
r.Äv	e->5	
r.Å 	a->2	
r.ÖV	P->1	
r: "	J->1	
r: A	n->1	
r: D	e->3	
r: F	i->1	r->1	ö->1	
r: I	n->1	
r: K	ä->1	
r: O	m->1	
r: P	å->1	
r: V	i->2	
r: a	n->2	t->2	
r: d	e->8	
r: e	n->2	
r: f	ö->3	
r: h	u->1	
r: i	n->1	
r: k	o->1	
r: n	u->1	
r: o	m->1	p->1	
r: t	i->1	
r: u	t->1	
r: v	e->1	i->4	
r: Ä	r->1	
r; a	t->1	
r; d	e->3	å->1	
r; e	n->1	
r; i	 ->1	n->1	
r; j	a->1	
r; m	e->1	
r; o	c->2	
r; v	i->2	
r?, 	r->1	
r?- 	(->1	
r?. 	(->1	
r?Bo	r->1	
r?De	t->2	
r?Dä	r->1	
r?Eu	r->1	
r?Fr	u->1	å->1	
r?Ha	r->2	
r?He	r->3	
r?Hu	r->1	
r?I 	e->1	m->1	
r?Ja	g->3	
r?Ka	n->1	
r?Ko	m->2	
r?Me	n->2	
r?Na	t->1	
r?Ni	 ->1	
r?Nä	s->1	
r?På	 ->1	
r?So	m->1	
r?Ta	c->1	
r?Ve	m->1	
r?Vi	 ->2	
r?Är	 ->2	
r?Äv	e->1	
rHer	r->1	
rJag	 ->1	
rMed	 ->1	
rNäs	t->2	
ra "	b->1	u->1	
ra -	 ->6	
ra 1	 ->1	0->1	5->1	6->1	
ra 2	 ->1	5->1	
ra 5	 ->1	5->1	
ra 7	0->1	
ra A	t->1	
ra B	a->1	
ra D	a->1	
ra E	E->1	U->4	u->13	
ra F	N->1	r->1	
ra I	n->1	s->2	
ra J	e->1	
ra L	i->2	o->1	
ra R	i->1	o->1	
ra T	y->2	
ra a	d->1	f->2	g->1	k->2	l->18	m->3	n->24	r->17	s->5	t->101	u->1	v->53	
ra b	a->8	e->50	i->6	l->2	o->1	r->6	u->1	y->1	ä->7	å->2	ö->2	
ra c	e->4	
ra d	a->9	e->260	i->9	j->2	o->1	r->3	u->1	y->1	ä->1	ö->1	
ra e	f->8	g->7	k->5	l->5	m->1	n->168	r->23	t->69	u->11	x->8	
ra f	a->22	e->5	i->1	l->6	o->6	r->54	u->4	ä->1	å->3	ö->163	
ra g	a->1	e->20	i->5	j->1	l->2	o->4	r->24	ä->7	å->13	ö->3	
ra h	a->13	e->20	i->3	o->6	u->16	ä->6	å->5	ö->2	
ra i	 ->43	a->1	c->1	d->3	f->1	g->2	h->1	l->2	n->53	
ra j	a->1	o->1	u->2	ä->2	
ra k	a->10	e->1	i->1	l->8	n->1	o->137	r->8	u->5	v->6	ä->4	
ra l	a->13	e->7	i->14	o->2	ä->29	ö->4	
ra m	a->6	e->92	i->41	o->9	y->22	ä->7	å->30	ö->10	
ra n	a->9	e->2	u->1	y->16	ä->14	å->33	ö->8	
ra o	b->5	c->56	f->4	k->1	l->11	m->54	n->1	p->2	r->29	s->11	t->1	
ra p	a->12	e->9	l->4	o->18	r->37	u->13	å->44	
ra r	a->10	e->44	i->9	o->2	u->2	ä->5	å->4	ö->1	
ra s	a->29	e->9	i->74	j->2	k->22	l->8	m->4	n->5	o->18	p->3	t->39	u->5	v->5	y->14	ä->27	å->27	
ra t	a->10	e->3	i->77	j->4	o->3	r->13	u->1	v->12	y->3	
ra u	n->23	p->17	r->3	t->26	
ra v	a->25	e->17	i->38	o->1	ä->25	å->8	
ra y	t->7	
ra Ö	s->3	
ra ä	g->2	n->22	r->30	
ra å	 ->1	r->33	t->19	
ra ö	g->3	k->1	n->1	p->1	r->1	s->2	v->19	
ra! 	D->1	
ra!M	ä->1	
ra".	.->1	D->1	
ra, 	1->1	a->9	b->1	d->5	e->1	f->5	g->2	h->4	i->6	k->2	m->8	o->9	p->1	s->5	u->4	v->5	ä->4	å->1	
ra. 	M->1	
ra.A	l->1	v->1	
ra.B	a->1	
ra.D	e->13	ä->3	
ra.E	G->1	n->5	
ra.F	ö->2	
ra.H	e->2	ä->1	
ra.I	 ->2	n->1	
ra.J	a->15	
ra.L	ä->1	å->2	
ra.M	e->3	i->1	å->1	
ra.N	a->1	u->1	ä->2	
ra.O	c->1	
ra.P	a->1	e->1	å->2	
ra.S	o->1	ä->1	
ra.U	n->1	
ra.V	a->1	i->4	
ra: 	I->1	V->1	g->1	r->1	s->1	u->1	Ä->1	
ra; 	f->2	
ra?A	n->1	
ra?D	e->1	
ra?J	a->1	
rabb	a->50	
rabe	h->5	
rabi	s->6	
rabl	a->1	
rabr	e->1	
rabs	t->2	
rabv	ä->1	
raca	 ->3	
rack	a->1	
raco	-->1	
rad 	A->1	a->14	b->6	d->3	e->6	f->10	g->2	i->14	k->7	m->8	n->1	o->5	p->8	r->2	s->11	t->6	u->2	v->4	y->1	ä->2	ö->9	
rad,	 ->3	
rad.	D->1	H->1	K->1	M->3	U->1	V->1	
rade	 ->201	,->6	.->11	n->3	r->12	s->26	t->3	
radi	k->16	o->2	t->19	
rado	x->6	
radv	i->3	
rael	 ->22	,->4	-->1	.->3	?->1	e->5	i->15	k->1	s->6	
raf 	o->1	
rafa	t->1	
raff	 ->2	,->1	-->2	a->4	b->1	l->1	p->2	r->28	
rafi	 ->1	.->2	k->9	n->1	s->10	
rafr	y->2	
raft	 ->38	,->9	.->5	?->2	e->26	f->12	i->34	s->10	t->5	v->8	
rag 	-->1	a->6	d->2	e->1	f->6	h->1	i->6	k->2	m->1	o->3	s->12	t->14	v->1	ä->3	å->2	
rag,	 ->2	
rag.	B->1	D->1	H->1	R->1	V->2	
rag:	 ->1	
raga	.->1	n->114	
rage	d->4	l->1	n->29	t->121	
ragi	s->6	t->12	
ragm	a->1	
ragn	a->1	i->48	
ragr	a->3	
rags	a->2	f->1	g->8	m->1	n->1	r->2	s->1	t->2	ä->3	
raha	n->1	
rahu	s->1	
rain	e->2	
rak 	h->2	i->1	k->1	l->1	m->1	s->2	v->1	ö->1	
rak,	 ->1	
rak.	D->2	T->1	
rak?	N->1	
raka	 ->2	m->1	s->1	
rake	l->1	t->2	
raki	s->1	
rako	p->5	
rakr	y->1	
raks	 ->3	
rakt	 ->5	.->1	:->1	a->35	e->3	f->1	i->39	ä->9	
ral 	I->2	b->1	d->1	f->1	p->2	r->2	s->3	å->1	
ral,	 ->1	
ral-	 ->6	
ral.	F->1	H->1	
rala	 ->36	,->2	s->6	t->1	
ralb	a->8	
rald	e->1	i->17	
rale	n->2	r->3	u->1	
ralf	ö->1	
rali	b->1	s->43	
rall	e->5	t->10	
rals	e->2	
ralt	 ->10	,->1	
ram 	"->1	-->4	8->1	D->1	a->6	b->3	d->19	e->56	f->41	g->2	h->8	i->15	k->4	l->3	m->13	n->6	o->10	p->6	r->5	s->26	t->47	u->2	v->7	ä->4	å->1	ö->2	
ram,	 ->28	
ram.	.->1	D->5	F->4	G->2	H->2	J->2	K->2	M->2	N->1	O->1	R->1	S->3	T->1	V->2	
ram?	J->1	V->1	
rama	n->1	r->8	t->6	v->3	
rame	n->60	t->2	
ramf	a->1	ö->145	
ramg	i->1	å->52	
ramh	ä->5	å->17	ö->2	
rami	d->1	
ramk	a->1	o->10	
raml	a->13	ä->8	
ramm	e->109	
ramn	i->2	
ramp	 ->2	e->3	l->8	r->12	
ramr	u->1	
rams	k->2	t->48	
ramt	 ->1	a->5	i->107	r->2	v->2	
ramu	t->1	
ramv	e->1	i->3	
ramå	t->22	
ramö	v->2	
ran 	H->1	a->10	f->5	g->1	h->1	i->1	j->1	m->1	o->8	s->2	t->3	u->1	v->1	ö->1	
ran,	 ->4	
ran-	 ->1	
ran.	)->1	D->2	F->1	N->2	
ran?	F->1	O->1	
rana	t->1	
ranb	i->8	
ranc	,->1	a->1	e->2	i->1	
rand	 ->4	.->1	a->2	e->777	i->2	m->1	o->14	r->10	s->1	
rang	e->6	
rani	n->1	u->2	
rank	r->43	
ranl	e->2	
rann	a->5	h->1	l->2	s->2	
rano	i->1	
rans	 ->4	,->3	.->3	c->7	e->2	i->7	k->90	l->2	m->5	p->108	v->6	
rant	 ->10	.->2	e->59	i->34	ö->3	
ranv	a->4	ä->18	
ranz	 ->3	
ranç	o->1	
raor	d->1	
rape	r->1	
rapp	o->109	
rapr	o->1	
rar 	-->1	1->1	3->1	E->3	I->1	P->1	R->1	S->1	a->42	b->5	d->70	e->25	f->20	g->2	h->16	i->42	j->15	k->11	l->2	m->27	n->12	o->24	p->17	r->4	s->24	t->28	u->5	v->20	y->1	ä->6	å->1	ö->4	
rar!	 ->18	J->1	M->1	T->1	
rar,	 ->31	
rar.	.->1	A->1	D->1	F->3	H->1	J->1	N->1	R->1	S->1	V->2	
rar:	 ->1	
rar;	 ->1	
rara	 ->1	
rarb	e->2	
rare	 ->38	,->4	.->3	n->1	s->1	
rark	i->4	
rarl	ä->1	
rarn	a->17	
rars	 ->1	
rart	,->1	e->1	r->1	
rarv	 ->1	,->2	.->1	e->1	
ras 	4->1	E->1	a->47	b->6	c->2	d->8	e->14	f->32	g->8	h->5	i->39	j->2	k->7	l->5	m->19	n->9	o->25	p->14	r->9	s->30	t->15	u->12	v->7	y->1	ä->3	å->3	ö->5	
ras!	D->1	G->1	
ras,	 ->23	
ras.	 ->2	A->1	B->1	D->10	E->2	F->4	G->2	I->4	J->3	M->3	N->1	P->2	S->3	U->1	V->8	Y->1	
ras;	 ->1	
rasa	d->2	s->1	t->1	
rasb	o->5	
rasc	h->3	
rase	r->1	
rash	a->1	
rasi	l->1	s->26	
rask	a->1	
rasm	a->1	
rass	l->1	o->1	t->1	
rast	 ->12	.->1	e->7	i->3	r->15	
rat 	-->3	A->1	E->2	F->1	S->1	a->10	b->5	d->14	e->9	f->10	g->1	h->6	i->8	k->5	l->2	m->6	n->3	o->9	p->3	r->1	s->15	t->4	v->6	å->1	
rat,	 ->14	
rat.	 ->1	.->1	B->1	D->3	E->1	H->1	J->3	K->1	T->1	V->1	
rat;	 ->1	
rata	 ->3	l->6	r->1	
rate	g->63	n->2	r->24	s->1	t->12	
rati	 ->14	"->1	,->3	.->9	e->3	f->14	n->24	o->69	r->1	s->95	v->24	
rato	g->2	m->4	r->3	
rats	 ->33	,->6	.->5	?->1	
ratt	a->1	r->1	
ratu	l->37	r->13	s->3	
ratö	r->2	
raum	a->1	
rav 	-->1	4->1	8->1	b->1	d->2	e->1	f->5	g->1	i->1	l->1	n->1	o->3	p->17	s->9	t->1	u->1	v->1	
rav,	 ->4	
rav.	(->1	.->1	D->2	E->1	R->1	
rav?	V->1	
rava	 ->1	l->1	r->1	
rave	n->27	r->5	t->16	
ravt	 ->1	
rax 	a->1	e->1	i->1	
raxi	s->8	
ray,	 ->1	
raça	 ->5	
rb, 	e->1	
rba-	,->1	
rbal	a->1	
rban	"->1	d->2	i->1	
rbar	 ->3	.->1	a->8	h->1	i->2	m->1	t->4	
rbas	t->1	
rbay	e->1	
rbed	ö->1	
rbeg	r->1	
rbeh	å->6	
rbel	a->3	
rbem	a->1	
rber	 ->2	,->3	a->1	e->27	n->2	
rbes	t->2	
rbet	a->134	e->214	s->221	t->1	ä->6	
rbi 	d->1	
rbif	a->2	
rbig	å->6	
rbih	a->1	
rbil	d->1	
rbin	d->22	
rbis	e->1	k->6	
rbju	d->33	
rbjö	d->1	
rble	v->1	
rbli	 ->8	c->1	r->6	
rblå	s->2	
rbri	n->1	t->14	
rbro	t->1	
rbru	k->1	
rbry	g->3	t->2	
rbrä	n->2	
rbud	 ->11	,->2	.->3	e->8	s->2	
rbun	d->12	
rbät	t->78	
rböl	d->1	
rbör	a->1	l->10	
rce 	b->1	
rcel	o->2	
rcen	t->1	
rcou	r->1	
rcyk	l->4	
rd -	 ->1	
rd 2	 ->1	
rd C	o->1	
rd I	n->2	
rd K	o->1	
rd a	n->1	r->1	t->4	v->5	
rd b	l->1	r->1	
rd d	e->1	ä->1	
rd e	f->1	k->1	l->1	n->1	u->1	
rd f	r->1	ö->9	
rd g	r->1	
rd i	 ->4	n->2	v->1	
rd j	a->1	
rd k	a->2	o->2	r->1	u->1	
rd m	a->1	e->2	i->2	
rd n	ä->1	
rd o	c->16	m->3	
rd p	r->1	å->1	
rd s	i->1	j->1	k->1	o->9	
rd t	a->1	e->1	i->3	
rd u	r->1	
rd v	a->2	i->4	
rd),	 ->1	
rd, 	b->1	d->2	h->1	m->2	o->5	s->4	t->2	ä->1	
rd-a	f->1	
rd-f	ö->1	
rd.B	e->1	
rd.D	e->5	ä->1	
rd.E	u->1	
rd.H	e->1	
rd.I	 ->1	
rd.J	a->1	
rd.U	n->1	
rd.V	i->2	
rd: 	"->2	
rd; 	d->1	i->2	
rda 	a->6	d->2	e->5	f->3	g->1	h->2	k->8	l->2	m->3	n->3	o->2	p->7	r->4	s->7	t->2	u->2	v->4	ä->1	
rda,	 ->5	
rda.	D->1	H->2	O->1	
rda?	D->1	
rdad	.->1	e->2	
rdag	 ->1	,->1	e->3	l->2	
rdal	a->4	y->2	
rdam	 ->9	,->3	.->1	e->4	f->27	r->1	
rdan	 ->5	.->3	d->7	i->1	s->1	
rdar	 ->5	,->1	e->4	
rdas	 ->1	.->1	t->2	
rdat	 ->3	s->1	
rdbr	u->56	ä->1	
rdbä	v->10	
rde 	K->1	a->4	b->5	d->12	e->8	f->7	g->3	h->9	i->14	j->3	k->9	m->7	n->3	o->3	p->7	r->8	s->9	t->5	u->6	v->14	
rde,	 ->3	
rde-	 ->1	l->1	
rde.	D->2	G->1	J->2	L->1	N->1	T->1	
rdea	u->1	
rded	e->2	
rdef	u->7	
rdeg	e->3	
rdel	 ->3	,->2	.->2	a->15	e->1	n->23	ö->1	
rdem	o->1	
rden	 ->23	,->3	.->5	a->4	n->1	s->3	t->25	
rder	 ->167	,->13	.->21	?->1	a->21	i->44	l->5	n->22	
rdes	 ->14	,->1	.->1	s->2	
rdet	 ->25	.->2	
rdeu	r->1	
rdfö	r->223	
rdhe	t->1	
rdig	 ->6	.->1	a->11	h->18	s->1	t->4	
rdin	ä->1	
rdir	l->2	
rdis	e->9	k->4	
rdit	a->1	
rdju	p->11	
rdku	s->1	
rdla	d->1	
rdli	g->7	s->1	
rdmå	n->1	
rdna	 ->7	c->2	d->10	n->2	r->5	s->2	t->3	
rdni	n->155	
rdo 	R->1	
rdom	 ->6	,->1	a->1	l->1	s->2	
rdon	 ->32	,->8	.->9	?->1	N->1	e->7	s->7	
rdor	 ->1	n->1	
rdra	 ->3	g->164	n->7	r->2	s->5	t->1	
rdre	 ->1	
rdri	f->3	k->2	n->1	v->13	
rdrö	j->1	
rds 	r->1	
rds-	 ->1	
rdsb	u->1	
rdsk	a->1	
rdsl	i->1	ö->2	
rdsm	y->1	å->1	
rdso	m->1	
rdsp	a->2	l->3	r->1	u->1	
rdss	k->1	t->2	
rdst	o->3	
rdsu	t->1	
rdsv	i->1	
rdti	d->1	
rdty	s->1	
rdub	b->2	
rdun	k->1	
rdvr	ä->1	
rdvä	n->1	s->1	
rdär	v->4	
rdöm	a->13	e->5	t->2	
rdör	r->1	
re -	 ->5	
re 1	1->1	5->1	
re 2	0->1	1->1	
re 3	5->1	
re 4	,->1	
re A	m->1	
re B	N->1	
re D	e->1	i->1	
re E	u->2	
re H	i->1	
re K	i->1	
re a	d->1	k->1	l->4	m->1	n->17	r->1	t->28	v->11	
re b	a->2	e->27	i->3	l->4	o->1	r->1	y->4	ä->1	å->1	ö->2	
re c	h->1	
re d	a->2	e->20	i->3	o->1	u->1	y->1	ä->1	å->1	
re e	f->2	k->3	l->7	m->1	n->13	t->6	u->4	x->2	
re f	a->7	e->1	i->4	j->1	l->1	o->2	r->37	u->1	y->2	å->4	ö->67	
re g	e->6	j->1	o->2	r->8	å->3	ö->1	
re h	a->24	e->2	i->2	o->1	u->2	ä->1	å->1	ö->2	
re i	 ->40	d->1	n->17	t->1	
re j	o->1	ä->2	
re k	a->18	l->1	o->29	r->5	u->5	v->1	ä->2	
re l	a->3	e->1	i->1	ä->5	ö->1	
re m	a->71	e->19	i->6	o->4	y->3	å->16	ö->2	
re n	i->4	u->1	ä->9	å->4	
re o	c->48	l->2	m->16	r->5	s->1	v->2	
re p	a->2	e->6	l->2	o->2	r->10	u->2	å->18	
re r	e->12	i->2	o->3	ä->4	
re s	a->9	e->6	i->16	j->1	k->17	l->1	m->1	n->1	o->38	p->2	t->16	u->1	y->4	ä->12	å->2	
re t	a->8	i->29	j->4	o->3	r->1	v->3	y->3	
re u	n->2	p->8	t->23	
re v	a->18	e->5	i->14	o->1	ä->2	
re ä	n->48	r->10	
re å	r->6	t->3	
re ö	k->2	n->2	p->6	v->1	
re!S	k->1	
re" 	s->2	
re",	 ->1	
re, 	A->1	D->1	F->1	H->1	a->3	b->5	d->2	e->2	f->3	h->5	i->5	j->1	k->2	m->10	n->3	o->11	p->5	s->11	u->3	v->7	ä->4	å->2	
re-A	t->1	
re. 	D->1	O->1	Ä->1	
re.A	l->1	t->1	
re.B	å->1	
re.D	e->19	ä->2	å->2	
re.E	f->2	n->1	u->2	
re.F	ö->3	
re.H	e->1	
re.I	 ->4	m->1	
re.J	a->8	
re.K	o->2	
re.M	a->2	e->4	i->2	
re.N	u->1	ä->1	
re.P	r->1	å->1	
re.R	o->1	å->1	
re.S	o->3	
re.T	i->2	r->1	
re.U	r->1	
re.V	a->1	i->5	å->1	
re.Ä	n->2	r->1	v->2	
re: 	b->1	d->1	
re?D	e->1	
re?K	a->1	
re?O	c->1	
re?V	i->1	
rea 	b->1	o->3	
reag	e->16	
reak	t->21	
real	 ->1	,->1	i->16	
ream	i->8	
reat	i->2	ö->1	
rebe	f->2	h->1	
rebi	l->1	
rebo	a->1	
rebr	å->2	
reby	g->23	
reci	r->1	s->49	
reck	 ->1	
reco	v->1	
rect	n->1	
recy	c->1	
red 	b->1	d->1	e->1	i->6	l->1	m->1	o->7	v->1	
red,	 ->1	
red.	D->1	H->2	I->1	
reda	 ->15	,->2	k->1	n->158	r->9	s->2	
redd	 ->21	a->13	e->4	
rede	l->5	n->2	r->10	
redg	a->1	
redi	e->2	t->2	
redj	e->73	
redl	i->10	
redn	i->8	
redo	 ->3	g->10	v->4	
redr	a->165	o->1	
reds	 ->2	,->1	.->1	a->4	b->2	f->3	k->2	p->23	s->28	u->1	
redu	c->4	
redö	m->2	
ree-	f->1	l->1	
ree.	D->1	
reel	l->4	
refa	l->20	
refe	r->7	
refl	e->7	
refo	r->134	
reft	e->13	
refu	s->1	
refö	l->1	
rege	l->50	r->282	
regi	,->1	c->1	m->3	o->251	s->20	
regl	e->126	
regr	i->1	
regå	e->15	n->2	
reha	b->1	v->1	
reis	k->1	
reju	d->4	
rejä	l->3	
reke	r->1	
reki	s->6	
rekl	a->17	
reko	m->67	n->6	r->2	
rekr	y->1	
rekt	 ->50	,->2	.->8	;->1	a->10	i->194	o->18	ö->1	
rekv	e->1	
rela	 ->1	t->26	
rele	g->1	v->9	
reli	g->30	k->1	m->3	
rell	 ->13	a->28	t->15	
rels	e->28	
relä	g->2	
rema	 ->2	
reme	n->1	
remh	ö->14	
remi	s->11	ä->10	
remo	t->19	
rems	-->1	a->2	
remt	 ->4	
remå	l->13	n->1	
ren 	-->2	2->1	H->1	K->1	V->1	a->10	b->6	d->4	e->9	f->39	g->3	h->15	i->18	j->1	k->5	l->1	m->6	n->2	o->35	p->7	r->2	s->23	t->5	u->4	v->5	ä->12	å->1	ö->1	
ren)	.->1	J->1	
ren,	 ->41	
ren.	)->5	.->1	A->1	D->8	E->1	F->1	H->2	I->3	J->5	K->1	M->2	O->2	R->1	T->2	V->3	Ö->1	
ren;	 ->1	
ren?	I->1	V->1	Ä->1	
rena	 ->11	d->16	n->5	r->15	s->1	
rend	 ->5	!->2	,->2	-->1	a->3	b->1	e->21	s->2	t->7	
reng	u->2	ö->3	
renh	e->24	
reni	n->22	
renk	l->8	
renl	i->9	
reno	v->3	
rens	 ->102	!->1	,->12	-->2	.->10	/->1	:->1	?->2	a->4	b->9	d->5	e->168	f->8	h->4	i->2	k->60	m->11	n->9	o->3	p->80	r->20	s->27	u->2	v->11	ä->2	
rent	 ->22	a->29	e->1	i->5	s->1	
renz	 ->12	)->2	,->3	F->1	b->1	
renö	r->3	
rep 	m->1	
repa	 ->15	,->1	d->8	r->21	s->7	t->5	
repn	i->1	
repp	 ->10	,->1	a->1	e->11	s->2	
repr	e->24	i->2	
repu	b->18	
rer 	-->1	a->5	b->1	d->1	e->2	f->2	g->1	h->3	i->8	k->1	m->2	o->18	p->1	s->26	u->1	v->1	ä->2	å->1	
rer!	 ->1	
rer,	 ->17	
rer.	D->6	E->2	J->1	K->1	P->1	T->2	V->3	
rera	 ->40	d->13	r->12	s->15	t->8	
reri	n->19	
rern	a->41	
rero	g->1	
rers	 ->1	
rerö	v->1	
res 	a->2	d->1	e->1	f->1	i->2	l->4	n->1	o->2	p->1	r->4	v->1	å->1	ö->1	
res,	 ->3	
resa	 ->12	,->2	.->1	n->1	t->6	
rese	n->48	r->9	
resi	d->10	
resk	r->28	
resl	a->24	o->11	å->69	
reso	l->100	n->4	r->1	
resp	.->2	e->81	o->4	r->9	
ress	 ->4	a->24	e->108	i->4	k->2	m->1	n->1	
rest	 ->2	a->6	e->12	i->1	n->1	r->4	s->1	ä->9	å->6	
resu	l->111	r->50	
resä	t->1	
ret 	(->1	-->2	1->10	a->6	b->1	e->1	f->30	g->2	h->3	i->9	k->3	l->2	o->13	p->2	r->2	s->7	t->6	u->3	v->1	ä->7	å->1	ö->1	
ret,	 ->11	
ret.	 ->1	D->5	E->1	F->1	I->1	J->4	L->1	M->1	T->2	V->2	
ret:	 ->1	
reta	 ->36	,->2	g->207	n->1	r->3	
rete	r->2	s->12	
reti	s->4	
reto	r->3	
retr	o->11	ä->74	
rets	 ->8	,->1	a->3	e->2	l->2	
rett	 ->10	.->1	i->2	o->3	s->1	
reur	o->1	
reus	s->1	
reut	b->1	v->3	
rev 	d->2	f->1	i->1	n->1	o->1	s->1	t->2	u->1	
rev.	F->1	
revi	d->17	s->18	
revl	i->3	å->1	
revo	l->1	
revs	 ->3	
rext	r->6	
rey 	C->3	
reye	r->3	
rez,	 ->1	
rfal	l->3	s->1	
rfar	a->76	e->25	i->2	n->1	t->1	
rfat	t->7	
rfek	t->7	
rfin	i->1	n->3	
rfir	a->2	
rfis	k->1	
rfjo	l->1	
rflu	t->14	
rfly	t->6	
rflö	d->1	
rfod	e->4	
rfog	a->18	
rfon	d->58	
rfor	d->6	m->1	s->22	
rfry	s->1	
rfrå	g->13	
rfun	n->2	
rfäk	t->1	
rfär	a->1	g->1	l->1	
rfån	g->1	
rföl	j->8	l->2	
rför	 ->317	,->8	.->1	:->2	?->3	a->5	d->1	e->4	i->12	m->1	t->3	v->1	
rg H	a->14	
rg a	v->1	
rg f	i->1	ö->1	
rg g	j->1	
rg i	 ->1	
rg k	r->1	
rg m	e->2	
rg o	c->1	m->7	
rg s	a->1	
rg t	i->1	
rg u	t->1	
rg ö	p->1	
rg, 	B->1	I->1	f->1	j->1	k->1	s->1	
rg.D	e->1	
rg.J	a->1	
rg.L	e->1	
rg.V	i->1	
rga 	f->1	
rgad	 ->1	
rgan	 ->15	"->1	,->6	.->1	e->9	i->66	
rgar	 ->1	d->1	e->72	i->1	n->89	s->7	
rgav	s->2	
rge 	e->1	o->1	v->2	
rge,	 ->1	
rgen	 ->1	s->6	
rger	 ->15	,->2	.->2	M->1	b->1	i->1	l->3	
rges	 ->2	,->1	
rgh.	V->1	
rgi 	b->1	g->2	h->1	l->1	m->1	o->4	s->3	
rgi,	 ->2	
rgi-	,->1	
rgi.	A->1	E->2	F->1	M->1	
rgia	g->1	n->6	
rgib	e->3	
rgic	e->1	
rgie	f->4	
rgif	o->1	t->2	ö->4	
rgii	m->1	
rgik	a->1	o->1	ä->37	
rgim	i->1	y->1	
rgin	 ->3	,->1	a->6	
rgio	r->2	
rgip	o->2	r->5	
rgis	e->4	k->1	n->1	ä->7	
rgiv	e->4	l->1	n->3	
rgiz	i->5	
rgiä	k->1	
rgiå	t->1	
rgli	g->3	
rglö	m->2	
rgmä	s->2	
rgne	 ->1	
rgo 	s->1	
rgon	 ->27	,->2	.->6	d->2	
rgot	 ->1	
rgri	p->14	
rgru	n->3	p->1	
rgrä	v->4	
rgsf	u->1	
rgum	e->17	
rgäl	l->1	
rgäv	e->1	
rgå 	t->1	
rgån	g->12	
rgår	 ->6	
rgåt	t->1	
rgör	 ->2	a->13	s->2	
rhan	d->98	
rhas	t->3	
rhav	e->1	
rhea	d->1	
rhet	 ->145	,->12	.->27	?->3	J->1	e->57	s->63	
rheu	g->2	
rhin	d->31	
rhis	t->1	
rhol	k->4	
rhop	p->12	
rhun	d->7	
rhus	 ->1	,->1	e->1	
rhäm	t->2	
rhän	;->1	g->2	
rhåg	o->2	
rhål	l->70	
rhög	h->2	
rhöl	l->4	
rhör	d->3	t->9	
ri -	 ->1	
ri 1	9->4	
ri 2	0->5	
ri 8	 ->2	
ri L	a->3	
ri V	a->1	
ri a	v->1	
ri b	e->1	
ri d	i->1	
ri e	n->1	t->1	
ri f	r->1	ö->4	
ri i	 ->3	n->4	
ri k	o->3	
ri m	e->1	o->1	å->1	
ri n	ä->2	
ri o	c->11	m->1	
ri r	ö->8	
ri s	e->1	k->1	o->6	
ri v	a->2	
ri ä	r->2	
ri ö	k->1	p->1	
ri!H	e->1	
ri, 	d->1	e->1	l->2	m->4	n->1	o->5	s->3	t->2	u->1	v->1	
ri- 	o->10	
ri.B	å->1	
ri.H	u->1	
ri.J	a->1	
ri.L	i->1	
ri.M	a->1	
ri.V	i->1	
ria 	-->1	P->1	a->2	d->2	f->2	i->2	m->1	o->3	r->10	s->2	t->1	v->4	å->1	
ria,	 ->4	
ria.	D->1	Ä->1	
rial	 ->12	,->2	.->5	e->4	
rian	e->3	
rias	 ->3	
riat	 ->2	.->1	i->2	
ribe	k->4	
ribl	a->6	
ribu	t->1	
rich	t->6	
rici	o->1	t->1	
rick	a->1	e->3	f->1	n->1	s->1	
rid 	i->1	m->8	s->1	
rid,	 ->1	
rid.	E->1	
rida	 ->6	n->13	s->1	
ridd	 ->2	
ride	n->2	r->24	
ridi	g->1	s->30	t->1	
ridl	i->1	
ridn	i->15	
rido	r->2	
rids	 ->4	
rie 	C->1	
rie-	s->1	
rief	i->1	
riel	l->15	s->6	
rien	 ->21	,->4	.->6	f->1	s->3	t->6	
rier	 ->30	,->5	.->5	a->2	n->18	
ries	m->1	
riet	 ->5	"->1	,->2	.->3	s->2	
rife	r->6	
rifi	e->1	n->1	
rifr	å->6	
rift	 ->4	.->1	e->13	i->1	l->8	s->3	
rig 	a->5	b->1	d->1	f->17	h->3	i->3	k->5	m->7	o->2	p->2	r->1	s->4	t->3	v->3	ä->1	å->1	
rig"	.->1	
rig,	 ->4	
rig.	J->1	
riga	 ->64	,->3	.->4	
rige	 ->6	.->2	n->38	r->1	t->12	
righ	e->51	t->3	
rigi	n->2	
rigj	o->1	
rigo	r->4	
rigs	h->1	s->1	
rigt	 ->43	,->3	.->1	
rigö	r->5	
riha	n->2	
rihe	t->116	
rik 	e->1	i->3	n->2	p->1	
rik,	 ->2	
rik.	F->1	G->1	
rika	 ->36	,->8	-->1	.->5	n->17	r->10	s->11	
rike	 ->56	,->15	.->20	:->1	E->1	F->1	N->1	d->10	r->13	s->50	t->17	
riki	s->49	
rikl	i->2	
riko	m->1	n->1	
rikt	 ->15	,->1	.->2	a->60	i->50	l->70	n->50	p->2	
ril 	1->1	f->1	u->1	
ril.	J->1	
rila	g->1	n->1	
rili	k->1	
rilj	o->1	
rilo	b->1	
rimi	n->27	t->1	
riml	i->23	
rimm	a->1	
rims	a->2	b->2	p->1	r->2	å->1	
rimå	l->1	
rin 	a->3	b->1	e->2	f->5	h->1	i->4	k->3	l->1	m->1	o->6	p->1	s->9	v->2	ä->2	
rin!	H->1	
rin,	 ->15	
rin.	 ->2	D->3	H->1	I->1	J->2	N->1	S->2	V->3	
rin:	 ->1	
rin?	P->1	
rinc	i->194	
rind	u->2	
rinf	ö->4	
ring	 ->300	!->1	"->2	)->1	,->39	.->51	;->2	?->3	a->191	e->142	g->2	s->458	å->1	
rinh	o->6	
rini	p->1	
rinn	a->1	
rino	 ->3	,->1	.->2	s->1	
rinr	a->13	e->1	ä->1	
rins	 ->9	e->1	t->8	
rint	a->1	e->5	
rinä	r->3	
rio 	f->1	u->1	
riod	 ->23	,->5	.->2	?->1	e->41	i->14	
rior	.->1	i->39	
riot	 ->2	i->1	
ripa	 ->15	,->1	.->1	n->19	s->1	
ripe	n->1	r->15	t->3	
ripi	t->2	
ripl	i->6	
ripn	a->1	
ripo	l->3	
rips	 ->1	
rirr	a->1	
ris 	(->1	P->1	f->3	h->2	i->2	k->2	l->1	m->1	o->1	s->2	u->1	v->1	ä->2	å->1	
ris,	 ->2	
ris.	J->1	S->1	
ris:	 ->1	
ris?	Ä->1	
risa	 ->1	
risd	i->5	
rise	k->2	n->6	r->20	s->2	t->7	
risf	ö->1	
risk	 ->24	,->3	.->1	a->33	b->4	e->54	f->4	h->6	k->3	n->1	t->9	u->1	v->3	
risl	ä->2	
rism	 ->11	,->4	.->7	e->8	
risn	i->1	
riso	m->1	n->3	
riss	i->1	t->1	ä->1	
rist	 ->25	a->15	d->11	e->45	f->8	h->1	i->4	s->2	ä->1	å->1	
risu	t->1	
rit 	a->2	b->2	d->1	e->13	f->7	g->1	h->3	i->5	k->4	l->2	m->8	n->2	o->2	p->5	r->2	s->9	t->3	u->1	v->2	
rita	n->16	s->1	t->1	
rite	r->57	t->128	
riti	k->16	m->3	s->33	
ritl	e->1	
rito	r->17	
ritr	e->1	
ritt	 ->3	,->1	.->1	e->2	i->17	
rium	 ->4	,->3	.->5	
riut	s->1	
riva	 ->30	n->3	s->3	t->21	
rivb	o->1	
rive	l->5	n->9	r->22	t->7	
rivi	l->19	t->8	
rivk	r->3	
rivn	a->4	i->5	
rivs	 ->13	,->1	.->1	
riär	e->3	p->1	
rièr	e->1	
riös	 ->1	a->3	t->4	
rja 	a->7	d->1	e->2	f->8	k->2	m->37	o->1	p->3	r->1	s->1	t->3	u->1	å->1	
rjad	e->10	
rjan	 ->17	,->2	
rjar	 ->16	.->1	
rjat	 ->9	.->2	s->1	
rjde	 ->1	
rje 	1->1	E->1	a->3	b->3	d->9	e->7	f->15	g->5	h->2	i->3	k->2	l->9	m->11	o->1	r->3	s->6	å->10	
rjer	 ->2	
rjni	n->4	
rk -	 ->2	
rk a	t->1	
rk b	e->1	y->1	
rk d	a->1	
rk e	l->2	n->1	
rk f	i->1	å->1	ö->3	
rk g	e->1	
rk h	a->1	
rk i	 ->6	n->5	
rk k	a->1	o->3	ä->1	
rk l	y->1	
rk m	e->2	å->1	
rk o	c->6	f->1	
rk p	o->2	å->3	
rk s	e->1	k->2	o->5	å->1	
rk t	i->2	r->1	
rk u	t->1	
rk v	i->4	
rk ä	r->2	
rk, 	d->1	g->2	m->1	o->1	s->1	ä->1	
rk-d	a->1	
rk.B	e->1	
rk.D	e->2	å->1	
rk.F	r->1	
rk.J	a->1	
rk.S	y->1	
rk.V	a->1	
rk?R	e->1	
rka 	-->2	1->1	2->1	E->1	a->3	b->2	d->8	e->2	f->11	h->2	i->9	k->6	l->1	m->4	n->2	o->6	p->4	r->3	s->7	t->9	u->2	v->3	ä->1	å->1	
rka,	 ->5	
rka.	H->1	
rkad	e->2	
rkan	 ->23	,->1	.->1	d->3	e->4	s->1	t->3	
rkap	i->1	
rkar	 ->59	,->1	a->5	e->31	n->35	
rkas	 ->10	,->1	.->1	s->2	t->16	
rkat	 ->3	,->1	a->13	e->2	s->5	
rkba	r->3	
rkbo	r->1	
rkda	m->1	
rke 	i->2	m->1	t->5	
rkef	ö->1	
rkel	 ->1	s->5	
rken	 ->29	,->1	.->1	
rkep	o->1	
rker	 ->7	a->7	i->3	
rkes	a->1	e->1	f->1	k->2	l->4	m->1	u->7	v->1	
rket	 ->34	,->6	s->2	
rki.	D->1	
rkie	t->35	
rkil	t->1	
rkin	 ->1	.->1	
rkis	k->7	
rkiv	 ->1	e->1	
rkki	 ->2	
rkla	g->6	r->78	s->1	
rkli	g->210	
rkly	v->1	
rklä	g->1	
rkme	n->2	
rkna	d->191	
rkni	n->35	p->3	
rkog	å->1	
rkol	l->1	
rkom	a->1	m->6	s->1	
rkon	f->1	t->2	
rkop	 ->1	
rkor	 ->1	,->1	t->2	
rkot	i->7	
rkov	 ->1	
rkra	n->1	
rkro	m->1	
rkrä	v->1	
rks 	b->1	g->1	o->2	t->1	
rks.	D->1	O->1	V->1	
rksa	m->104	n->1	
rkst	ä->19	
rkt 	E->3	a->3	b->6	c->1	d->2	e->1	f->2	i->2	k->1	m->5	o->2	p->2	r->2	s->6	v->1	ö->3	
rkt,	 ->1	
rkt.	D->2	
rkta	 ->18	
rkts	 ->1	
rkty	g->8	
rkul	a->1	e->2	
rkun	n->2	
rkur	s->1	
rkän	d->5	n->35	t->2	
rköt	t->1	
rl H	e->1	
rl o	c->1	
rl v	o->3	
rl-H	e->1	
rlag	 ->4	,->1	.->2	d->1	e->1	o->2	t->3	
rlam	e->600	
rlan	d->25	g->6	
rld 	W->1	s->1	
rld,	 ->2	
rld.	J->1	
rlde	n->37	
rlds	d->1	e->1	f->1	h->4	k->6	l->1	m->1	n->1	o->1	
rled	a->1	i->1	
rleg	a->2	
rlek	e->2	
rlev	a->2	e->3	n->4	s->1	
rlig	 ->29	!->1	,->4	.->2	:->1	a->123	e->56	g->1	h->26	t->177	
rlik	a->2	n->44	
rlin	 ->4	,->2	.->1	g->2	
rlis	t->2	
rlit	a->6	l->4	
rliv	,->1	.->1	a->19	
rlor	a->20	
rlsr	u->2	
rlun	d->3	
rlus	t->10	
rlys	e->1	t->1	
rläg	g->9	s->2	
rläk	t->1	
rläm	n->18	
rlän	d->36	g->4	
rlär	l->1	
rlät	t->18	
rlåt	a->7	e->3	i->2	l->2	s->1	
rlös	t->2	
rløn	,->2	
rm a	t->2	v->24	
rm b	e->1	
rm d	a->1	ö->1	
rm e	l->5	
rm f	ö->3	
rm i	 ->3	
rm j	u->1	
rm k	a->1	o->3	
rm l	ö->1	
rm o	c->3	
rm p	å->1	
rm s	k->2	o->4	p->1	
rm v	i->2	ä->1	
rm ä	r->1	
rm ö	v->1	
rm, 	e->2	f->1	m->1	o->2	s->1	u->1	ä->1	
rm-e	l->1	
rm.D	e->1	
rm.E	G->1	
rm.M	e->1	
rm.N	u->1	
rm.S	a->1	
rm.V	i->1	
rm.Ä	r->1	
rm: 	e->1	
rma 	M->1	b->3	d->3	e->1	f->3	k->4	m->3	p->1	s->6	u->1	v->1	å->1	ö->1	
rma.	O->1	
rmac	e->1	
rmad	e->5	
rmaj	o->1	
rmak	o->1	
rmal	a->2	i->4	t->5	
rman	 ->1	.->1	d->6	e->8	s->2	
rmar	 ->12	b->3	e->15	n->13	
rmas	 ->3	t->13	
rmat	 ->8	e->1	i->74	s->1	
rmed	 ->47	,->2	l->3	
rmel	l->16	s->1	
rmen	 ->13	,->2	.->3	a->2	i->1	s->5	
rmer	 ->57	,->4	.->12	a->26	i->17	n->18	
rmfä	l->1	
rmfö	r->2	
rmid	d->12	
rmin	e->1	i->10	n->1	
rmis	.->1	t->1	
rmni	n->31	
rmo,	 ->1	
rmod	 ->1	i->1	l->12	
rmon	b->1	i->18	
rmor	g->1	
rmou	t->1	
rmpa	k->1	
rmpr	o->14	
rmra	p->2	
rmsi	g->2	
rmst	a->1	ä->1	
rmt 	a->3	d->1	e->2	h->1	m->1	o->3	t->5	u->1	v->2	
rmul	e->18	
rmyn	d->15	
rmäs	s->1	
rmå 	b->1	r->1	
rmåg	a->31	
rmål	i->1	
rmån	 ->11	e->2	s->1	
rmår	.->1	
rmåt	g->1	
rmé 	o->1	
rmén	 ->1	.->1	
rmög	n->1	
rmöt	e->2	
rn (	f->1	
rn -	 ->4	
rn E	r->2	
rn b	i->1	ö->1	
rn d	e->1	ä->1	
rn e	l->1	n->2	
rn f	i->1	o->1	r->1	ö->7	
rn g	r->1	
rn h	a->3	
rn i	 ->4	n->2	
rn k	a->1	o->4	
rn l	i->2	
rn m	e->1	
rn n	y->1	
rn o	c->14	m->2	
rn p	å->1	
rn r	e->1	
rn s	a->2	k->3	o->3	t->1	ä->1	å->2	
rn t	a->1	o->1	
rn u	n->2	
rn v	a->1	i->1	
rn ä	r->3	
rn).	D->1	
rn, 	B->1	R->1	a->1	e->1	f->1	h->1	i->5	j->1	m->4	o->3	s->3	v->2	
rn- 	o->2	
rn.)	 ->1	
rn..	 ->1	
rn.D	e->7	ä->1	
rn.F	ö->3	
rn.H	e->2	
rn.J	a->1	u->1	
rn.K	o->1	
rn.M	i->1	
rn.O	m->1	
rn.V	i->1	
rn.Ö	g->1	
rn/N	o->2	
rn?A	n->1	
rna 	(->1	-->18	1->5	3->1	6->1	8->8	A->1	I->1	P->1	T->1	a->95	b->33	d->28	e->27	f->187	g->30	h->60	i->205	j->3	k->48	l->10	m->75	n->14	o->184	p->34	r->12	s->129	t->55	u->39	v->35	ä->53	å->3	ö->8	
rna!	D->1	H->1	O->1	
rna"	.->2	i->1	
rna,	 ->221	
rna.	 ->5	(->1	)->1	-->1	.->1	A->9	B->2	D->63	E->11	F->15	G->2	H->9	I->15	J->24	K->10	L->4	M->19	N->7	O->5	P->5	R->1	S->11	T->4	U->5	V->35	Ä->3	Å->1	
rna/	s->1	
rna:	 ->3	
rna;	 ->4	
rna?	E->1	H->2	I->1	J->2	M->1	V->4	Ä->1	
rnaH	e->1	
rnad	e->1	
rnag	e->1	
rnal	i->2	
rnam	n->1	
rnan	 ->6	
rnar	 ->4	d->1	e->1	
rnas	 ->216	,->2	.->1	
rnat	i->94	
rnba	r->1	
rnd 	L->3	
rne 	o->1	
rne,	 ->1	
rnea	r->1	
rned	r->2	
rnek	a->8	
rnen	e->8	
rner	 ->1	i->2	n->1	
rnet	 ->4	,->4	.->3	
rnfr	e->1	å->2	
rnhi	l->1	
rnie	r->14	
rnin	g->27	
rnis	e->24	
rnit	i->1	
rniv	å->1	
rnié	 ->1	
rnka	t->1	
rnkr	a->22	
rnog	r->2	
rnpo	r->2	
rnpr	i->2	
rnpu	n->2	
rns 	a->1	d->1	f->3	h->1	n->1	o->2	p->3	s->4	u->1	v->1	
rnst	e->1	r->1	
rnsä	k->3	
rnt 	s->3	u->1	
rnt.	S->1	
rnte	k->2	n->1	
rntu	n->1	
rnuf	t->14	
rnva	p->8	
rnvä	g->15	
rnya	 ->1	n->1	r->1	s->1	
rnyb	a->39	
rnye	l->6	
rnät	e->1	
rnöd	v->1	
rnör	,->1	
ro -	 ->2	
ro 1	9->1	
ro E	u->1	
ro a	t->4	
ro b	e->1	l->1	
ro d	e->1	i->1	
ro f	u->1	ö->10	
ro h	a->1	
ro i	 ->6	
ro l	e->1	
ro m	e->1	å->1	
ro n	ä->2	å->3	
ro o	c->5	m->1	
ro p	e->2	å->4	
ro s	o->12	
ro t	i->2	r->1	
ro u	n->1	
ro v	a->1	
ro ä	r->3	v->1	
ro ö	v->1	
ro!A	l->1	
ro, 	d->1	f->2	h->1	k->1	o->3	s->4	t->1	v->1	ä->1	
ro-r	å->1	
ro.A	t->1	
ro.B	e->1	
ro.D	e->2	ä->1	
ro.F	l->1	ö->1	
ro.H	u->1	
ro.J	a->2	
ro.K	n->1	
ro.N	ä->1	
ro.O	m->1	
ro.S	e->1	
ro.T	r->1	
ro.V	i->3	
roa 	f->1	o->1	s->1	
road	 ->3	e->2	
roak	t->12	
roan	d->9	s->1	
roar	 ->5	
roat	e->1	
robl	e->183	
roce	d->1	n->94	s->109	
rock	s->1	
roda	c->5	s->4	
rodd	a->1	e->8	
rode	r->2	
rodi	 ->17	,->1	.->2	;->1	s->7	
rodu	c->31	k->53	
roed	t->14	
roek	o->5	
roen	d->127	
rof 	-->1	a->1	e->2	f->5	h->2	i->3	k->1	l->1	o->2	s->4	u->1	ä->1	
rof,	 ->4	
rof.	D->2	E->1	J->1	
rofa	l->1	
rofd	r->1	
rofe	d->1	n->20	r->31	s->7	
rofh	j->1	
rofi	l->3	n->1	
rofs	i->1	t->3	
rofö	r->1	
rog 	a->1	f->1	s->1	t->2	
roga	n->2	t->1	
rogb	e->1	
roge	n->1	r->1	t->1	
rogk	u->1	
rogr	a->238	e->1	u->1	
rogs	 ->2	
rois	k->1	
roje	k->64	
rojk	a->1	
roju	s->6	
rok 	d->1	f->2	g->1	o->1	s->1	
rok,	 ->3	
roki	g->2	
rokl	a->1	
rokr	e->2	
rol,	 ->1	
rol.	M->1	
role	u->1	
roli	g->18	
roll	 ->87	!->1	,->19	-->1	.->25	:->1	a->1	e->86	f->1	m->4	o->2	s->3	u->14	v->1	
rolä	m->2	
rom 	d->1	g->1	
rom,	 ->1	
roma	d->1	
rome	r->9	t->1	
romi	s->22	
romr	å->3	
roms	 ->1	a->4	v->1	
ron 	-->1	a->4	e->1	f->2	o->1	p->1	s->1	ä->1	ö->1	
ron,	 ->3	
ron-	 ->1	
rona	z->1	
rong	e->1	
roni	.->1	k->1	s->10	
ronj	u->1	
ronm	ä->2	
rono	d->3	m->1	
rons	 ->3	
ront	a->1	e->3	
room	r->1	
rop 	o->2	s->1	
rop,	 ->1	
rop.	S->1	
ropa	 ->141	!->2	"->1	,->36	.->60	;->1	?->3	N->1	d->2	g->5	k->1	m->1	n->1	p->166	r->4	s->48	t->1	v->3	
rope	i->712	t->1	
ropo	l->16	r->9	
ropp	e->2	
ropr	o->1	
ropå	 ->1	
ropé	 ->1	e->9	
ror 	-->1	a->81	d->8	e->1	f->2	g->1	i->14	j->24	k->2	m->5	n->5	o->7	p->11	s->5	t->2	u->2	v->3	ä->4	ö->1	
ror,	 ->4	
ror.	J->1	N->1	S->1	V->2	
ror?	H->1	
rord	a->2	n->47	
rore	n->28	
rori	s->10	
rorn	a->6	
rors	a->6	
ros 	f->1	m->1	o->1	s->1	
rosa	t->1	
rose	n->1	
rosk	e->3	
rosm	o->4	
ross	a->1	e->2	t->1	
rost	a->2	b->1	i->1	
rot.	J->1	
rota	 ->3	d->2	r->2	s->5	t->1	
rote	k->4	s->9	
rotf	ä->1	
roth	e->1	
rotn	i->17	
roto	k->26	
rots	 ->63	y->1	
rott	 ->14	,->9	.->5	a->2	e->4	m->1	s->27	
rotu	l->1	r->1	
rouk	 ->1	
roup	 ->1	
roux	-->1	
rov 	f->4	o->2	p->9	s->1	
rov"	,->1	
rov,	 ->1	
rov.	 ->1	D->1	
rova	n->3	
rove	r->4	t->3	
rovi	c->1	n->3	s->2	
rovk	a->1	o->1	
rovs	i->1	k->2	t->1	
rovä	c->3	r->15	
rpa 	a->1	b->1	d->1	h->1	k->1	t->1	
rpac	k->5	
rpar	l->1	t->2	
rpas	 ->1	?->1	s->1	
rpeg	n->1	
rper	s->1	
rpet	 ->2	
rpla	n->1	
rpli	k->21	
rpni	n->1	
rpol	-->1	i->20	
rpop	u->1	
rpos	t->2	
rpre	s->1	
rpri	s->1	
rpro	g->3	j->1	
rpt 	d->1	f->1	
rpta	 ->2	
rpus	 ->5	
rpå 	k->1	t->1	
rqui	o->1	
rr A	l->1	
rr B	a->2	e->5	o->3	
rr C	o->3	
rr E	v->2	
rr F	r->1	
rr G	o->1	r->1	
rr H	ä->2	
rr J	o->1	
rr K	i->4	o->2	
rr L	a->1	
rr M	o->1	
rr N	o->1	
rr P	a->3	o->5	
rr R	a->1	
rr S	c->2	e->2	p->1	
rr W	y->1	
rr a	l->1	
rr b	a->1	l->1	ö->1	
rr d	e->3	å->1	
rr e	l->2	
rr f	i->1	o->1	ö->6	
rr g	e->1	ö->1	
rr h	a->6	
rr i	 ->1	n->4	
rr k	a->2	o->83	
rr l	e->15	
rr m	i->2	
rr n	ä->1	
rr o	c->1	f->1	r->5	
rr p	a->3	
rr r	å->12	
rr s	a->1	e->1	t->1	ä->1	
rr t	a->319	j->1	
rr v	a->3	
rr ä	n->1	r->3	v->1	
rr å	t->1	
rr ö	p->1	
rr, 	i->2	m->1	ä->1	
rr.V	i->1	
rr?V	i->1	
rra 	T->1	d->2	k->6	m->2	o->1	p->2	r->1	s->1	v->13	å->19	
rrad	 ->1	e->1	
rrai	n->2	
rran	d->3	g->6	
rrar	 ->10	!->20	,->16	.->1	;->1	n->2	
rras	 ->1	,->1	k->1	
rrat	.->1	i->2	s->1	
rre 	-->2	a->7	b->4	d->3	e->2	f->4	h->2	i->3	j->2	k->2	l->2	m->4	o->6	p->4	r->4	s->10	t->1	u->8	v->6	ä->3	ö->6	
rre,	 ->1	
rrec	t->1	
rref	o->1	
rreg	e->3	l->3	
rrek	t->27	
rren	 ->2	,->3	s->278	t->2	
rrep	a->1	r->2	
rrer	a->5	
rres	 ->1	p->1	t->4	
rrey	 ->3	
rrez	,->1	
rrgå	n->1	r->3	
rrid	o->2	
rrik	a->7	e->74	i->49	
rrin	g->9	
rris	 ->1	
rrit	a->1	e->3	o->17	
rriä	r->4	
rrog	a->2	
rron	g->1	
rror	.->1	i->10	
rrum	p->2	
rrup	t->7	
rrva	r->1	
rräd	e->1	
rrän	 ->4	
rrät	t->2	
rråd	 ->1	,->1	e->13	
rrón	 ->3	
rrör	 ->4	
rrös	t->1	
rs 1	9->1	
rs 2	0->1	
rs E	G->1	U->1	
rs a	l->1	n->8	r->3	t->1	v->18	
rs b	a->1	e->13	i->1	r->1	u->3	y->1	
rs d	e->6	u->1	ö->2	
rs e	f->1	k->3	n->5	r->2	t->2	
rs f	l->5	o->1	r->7	u->4	ö->8	
rs g	i->1	o->1	r->1	
rs h	a->7	j->1	ä->4	
rs i	 ->16	n->7	
rs j	u->1	
rs k	a->4	o->5	
rs l	e->2	i->3	ä->1	ö->1	
rs m	e->3	o->1	å->4	
rs n	a->2	e->1	i->1	
rs o	a->1	c->7	f->1	k->1	l->1	r->1	
rs p	a->6	l->1	o->1	r->2	å->5	
rs r	a->1	e->2	o->1	ä->4	
rs s	a->1	i->2	k->4	o->4	t->3	y->1	ä->2	å->2	
rs t	a->1	i->6	o->1	r->1	y->1	
rs u	n->1	p->2	t->8	
rs v	a->2	ä->1	
rs y	r->1	
rs ä	g->1	r->2	
rs å	s->1	t->1	
rs ö	k->1	p->1	v->3	
rs, 	L->1	a->2	e->1	f->2	i->1	k->2	m->2	o->6	p->1	s->1	ä->1	
rs-b	i->1	
rs. 	E->1	
rs..	(->1	
rs.D	e->9	
rs.H	e->1	
rs.J	a->3	
rs.M	e->1	
rs.N	u->1	
rs.O	n->1	
rs.T	y->1	
rs.U	t->1	
rs.V	i->3	å->1	
rsaf	t->1	
rsai	l->1	
rsak	 ->1	.->2	a->18	e->17	
rsal	m->1	
rsam	l->13	m->7	t->1	
rsan	a->1	
rsat	t->5	
rsav	g->1	
rsbe	f->2	l->1	r->1	s->1	
rsbr	i->1	
rsbu	d->1	
rsch	e->1	
rsda	g->8	
rse 	d->1	f->2	k->1	o->2	s->1	
rse,	 ->1	
rse.	D->1	V->1	
rsei	l->1	
rsek	t->5	
rsel	!->1	l->3	
rsen	 ->6	,->1	a->14	i->13	
rser	 ->28	,->3	.->7	n->17	
rses	 ->1	
rsfr	i->43	å->4	
rsfu	l->4	
rsfö	r->5	
rshi	p->1	
rsie	l->9	
rsif	i->2	
rsik	t->85	
rsin	r->1	
rsio	n->13	
rska	l->4	p->33	r->5	s->1	
rski	l->161	n->2	
rskj	u->1	
rskn	i->35	
rsko	n->1	t->2	
rskr	i->19	o->2	ä->4	
rskt	 ->1	
rsku	l->2	
rskä	m->1	n->3	
rskå	d->6	r->1	
rsla	g->494	n->1	
rsli	n->1	
rslu	n->1	
rsma	k->1	
rsme	d->1	
rsmi	n->1	
rsmä	n->1	
rsmå	l->1	
rsom	 ->189	,->1	r->7	
rson	 ->6	,->1	a->24	e->43	i->4	l->34	s->1	
rsor	d->1	
rsot	 ->1	
rspe	g->3	k->17	r->3	
rspo	l->4	r->1	s->1	
rspr	o->1	u->19	
rspå	r->1	
rsra	p->2	
rssk	i->2	
rssl	ö->1	
rst 	a->9	c->1	d->3	e->4	f->1	g->2	h->2	i->5	j->1	k->2	m->4	n->3	o->23	p->1	r->3	s->13	t->3	u->1	v->14	
rst.	M->2	
rsta	 ->229	,->10	:->5	;->2	b->1	d->1	g->1	i->22	k->1	t->5	
rste	 ->1	
rsti	d->2	g->5	l->1	
rstk	l->1	
rsto	d->3	l->1	
rstr	e->1	y->27	ä->12	ö->2	
rstä	d->2	l->41	r->29	
rstå	 ->20	,->1	.->2	d->2	e->14	n->9	r->42	s->4	t->10	
rstö	d->9	r->21	
rsum	b->1	m->8	
rsun	d->3	
rsva	g->21	r->41	
rsvi	n->15	
rsvu	n->4	
rsvä	m->7	
rsvå	r->2	
rsyd	d->1	
rsyn	 ->1	t->1	
rsäk	r->44	t->15	
rsäl	j->5	
rsäm	r->10	
rsän	d->1	k->1	
rsät	t->35	
rsåg	s->1	
rsåt	e->1	
rsök	 ->5	,->2	a->41	e->20	n->23	t->18	
rsör	j->4	
rsöv	e->1	
rt -	 ->6	
rt C	a->1	
rt D	u->1	
rt E	G->1	u->4	
rt F	P->1	
rt G	o->1	
rt a	g->2	l->1	n->16	r->10	t->89	v->33	
rt b	a->1	e->12	i->3	l->1	o->1	r->1	u->1	ä->2	ö->2	
rt d	e->23	j->1	r->2	y->1	ä->1	
rt e	g->5	k->4	l->1	m->2	n->13	r->3	t->10	u->3	x->1	
rt f	a->6	i->3	r->11	å->2	ö->50	
rt g	e->8	o->1	r->3	å->2	
rt h	a->5	e->1	i->1	o->3	u->3	ä->1	å->1	
rt i	 ->13	f->1	n->23	
rt k	a->2	l->2	n->1	o->9	r->4	u->3	ä->1	
rt l	a->3	i->1	o->1	y->1	ä->3	ö->2	
rt m	a->4	e->20	o->2	y->2	å->8	ö->1	
rt n	e->1	u->1	y->2	ä->2	å->8	
rt o	c->41	l->1	m->15	r->6	s->2	
rt p	a->14	e->2	o->4	r->6	å->9	
rt r	e->6	i->1	ä->1	
rt s	a->12	e->5	i->11	k->7	l->1	o->24	p->2	t->14	v->8	y->3	ä->10	å->4	
rt t	a->10	e->2	i->4	o->2	r->1	y->1	
rt u	n->5	p->2	t->21	
rt v	a->2	e->3	i->8	ä->2	å->1	
rt y	t->2	
rt Ö	s->1	
rt ä	m->1	n->2	r->6	
rt å	t->1	
rt ö	g->1	v->2	
rt!H	e->1	
rt!J	a->1	
rt) 	t->1	
rt, 	a->1	b->2	c->1	d->2	e->4	g->2	h->6	i->1	k->2	l->1	m->7	n->1	o->6	p->1	s->3	t->3	v->4	ä->2	
rt- 	o->1	
rt-s	t->2	
rt. 	7->1	I->1	
rt.A	r->1	
rt.D	e->7	i->1	å->1	
rt.E	n->1	
rt.F	r->1	ö->1	
rt.H	ä->1	
rt.I	 ->2	
rt.J	a->6	u->1	
rt.K	o->3	
rt.L	å->1	
rt.M	e->2	
rt.N	i->1	
rt.O	c->1	
rt.R	i->1	
rt.S	a->1	l->1	t->1	
rt.U	t->1	
rt.V	a->1	i->6	
rt.Ä	v->1	
rt: 	E->1	e->1	
rt?J	a->1	
rtNä	s->1	
rta 	a->1	d->1	e->1	f->4	k->1	m->1	o->3	p->1	r->1	s->1	t->1	u->1	ä->1	
rtab	l->1	
rtad	 ->2	e->3	
rtag	,->1	a->8	n->1	
rtal	 ->3	a->1	e->4	
rtam	e->1	
rtan	d->1	k->3	n->3	s->2	
rtar	 ->2	,->1	.->2	
rtas	 ->3	t->1	
rtat	 ->10	,->1	.->2	:->1	s->2	
rtbe	s->2	
rtbi	l->1	
rtdi	r->1	
rtec	k->24	
rtel	l->15	
rtem	e->9	
rten	 ->43	,->3	.->5	:->1	d->1	s->3	
rter	 ->37	,->7	.->12	a->22	i->1	n->30	
rtet	 ->15	.->1	s->3	
rtex	t->3	
rtfa	l->6	r->89	t->2	
rtfe	d->1	
rtfr	å->1	
rtfö	r->1	
rtgr	u->4	
rtgå	.->2	e->3	
rthe	t->1	
rthu	 ->1	
rthy	 ->1	
rti 	a->1	d->1	f->2	h->2	i->4	k->1	m->1	p->1	s->7	t->2	å->1	
rti,	 ->7	
rti.	.->1	D->1	H->1	K->1	
rtid	 ->66	,->3	s->6	
rtie	l->2	r->10	t->30	
rtif	i->8	
rtig	h->1	
rtii	n->1	
rtik	a->3	e->95	l->15	r->1	
rtil	e->1	l->3	
rtin	e->1	o->1	
rtio	 ->3	n->10	s->1	
rtip	r->2	
rtis	 ->2	,->1	.->1	k->3	p->1	
rtju	s->1	
rtjä	n->20	
rtko	m->17	s->2	
rtle	v->1	
rtli	g->7	
rtlä	g->1	
rtma	r->1	
rtmo	n->1	
rtne	r->28	
rtni	n->2	
rtnä	t->1	
rtog	 ->1	
rtom	 ->15	!->1	,->3	.->1	r->3	
rton	 ->8	d->1	e->1	h->1	
rtpl	a->1	
rtpr	i->1	o->1	
rtra	k->1	m->1	n->1	p->1	r->1	
rtre	g->1	
rtro	e->56	g->1	s->2	t->1	
rtry	c->2	
rträ	d->6	f->3	n->1	
rtrö	t->1	
rts 	"->1	a->13	c->1	d->3	e->2	f->6	h->4	i->6	m->2	n->1	o->6	p->2	s->1	t->1	u->1	v->2	
rts,	 ->6	
rts.	D->1	J->2	S->1	T->1	V->1	
rtsa	m->1	t->12	
rtse	 ->4	r->1	t->1	
rtsi	f->1	k->4	n->1	
rtsk	r->1	
rtsm	e->1	y->1	
rtso	r->2	
rtss	e->3	
rtsä	k->7	t->82	
rtug	a->26	i->70	u->1	
rtun	i->2	
rtus	e->3	
rtut	s->2	
rtvi	n->1	v->1	
rtyd	l->3	
rtyg	 ->28	)->1	,->3	.->4	;->1	a->34	e->24	s->12	
rtyr	e->1	
rtz 	o->1	s->1	
rtz,	 ->1	
rtäc	k->1	
rtän	k->2	
ru A	h->2	n->1	
ru B	e->1	
ru F	r->1	
ru L	y->1	
ru M	c->1	
ru P	e->1	l->1	
ru R	e->3	
ru S	c->3	u->1	
ru T	h->1	
ru W	a->1	
ru k	o->46	
ru l	e->2	
ru t	a->83	
ru, 	s->1	
ruar	i->16	
rubb	a->3	
rubr	i->2	
ruck	i->1	n->1	
ruer	a->5	
ruhe	 ->1	,->1	
ruin	e->1	
ruk 	a->1	m->1	o->5	p->1	s->1	
ruk!	A->1	
ruk,	 ->9	
ruka	d->2	r->14	s->1	
ruke	n->1	t->19	
ruki	t->1	
rukn	i->1	
ruks	e->1	f->2	l->1	o->2	p->9	r->2	s->6	
rukt	 ->1	.->1	a->11	b->2	e->1	i->30	u->153	ö->3	
rull	a->3	s->3	
rum 	e->1	f->7	h->2	i->18	m->1	o->4	p->3	u->2	y->1	å->1	
rum!	M->1	
rum,	 ->5	
rum.	 ->1	D->1	M->1	O->1	
rume	n->52	t->3	
rump	e->2	
runa	 ->1	
rund	 ->107	,->1	.->1	?->1	a->30	b->1	e->38	f->4	k->1	l->90	o->1	p->2	r->2	s->2	t->1	v->25	
rung	 ->2	.->2	e->2	l->12	s->1	
runk	n->3	
runo	 ->1	
runt	 ->4	.->1	a->3	o->1	p->1	
rupp	 ->56	,->9	.->2	?->1	b->12	e->120	k->1	l->1	o->1	r->7	s->7	t->12	u->1	v->1	
rupt	i->7	
rusa	 ->1	l->2	r->2	
rust	a->3	b->1	e->4	n->5	r->2	
rut 	a->1	o->1	
rut.	D->1	
ruta	l->2	
rutb	e->1	i->2	
rute	a->3	n->1	t->1	
rutg	i->1	
ruti	n->8	t->2	
ruto	m->15	
ruts	a->1	e->8	k->1	ä->54	
rutt	e->1	n->2	o->1	
rutv	a->2	e->2	
rutö	v->1	
ruva	 ->1	
ruvi	d->15	
rv f	å->1	
rv o	c->2	
rv, 	a->1	e->1	s->1	
rv."	D->1	
rv.B	a->1	
rv.E	n->1	
rva 	d->1	f->1	n->1	o->1	p->1	r->1	
rvad	e->1	
rvak	a->14	n->11	
rval	 ->3	e->1	s->1	t->49	
rvan	d->4	s->2	
rvar	a->42	e->1	n->1	o->4	r->1	
rvat	 ->1	i->9	s->1	t->17	ö->1	
rvbr	i->1	
rvec	k->1	
rven	 ->3	.->3	e->2	t->5	
rver	 ->3	a->2	k->23	
rvet	 ->3	,->1	e->1	
rvhe	t->1	
rvic	e->7	
rvid	 ->8	l->1	
rvin	n->74	
rvir	r->12	
rvis	 ->1	a->2	s->8	
rvju	 ->2	a->1	
rvli	g->2	
rvri	d->1	
rvrä	n->1	
rvsa	r->3	
rvsi	n->1	
rvss	t->2	
rvt 	p->2	
rvtr	u->1	
rvun	n->3	
rväg	 ->5	,->4	.->2	a->25	d->1	e->7	r->3	t->2	
rväl	d->3	
rvän	d->3	t->29	
rvär	d->5	l->2	r->4	t->1	v->7	
rvån	a->6	
rwel	l->1	
ry F	o->1	
ry o	c->1	
ry, 	H->1	
ry.D	e->1	
ryck	 ->24	,->2	.->1	a->23	b->1	e->19	l->13	n->5	s->3	t->14	
ryft	a->1	
rygg	a->6	e->3	h->6	r->1	
rygt	 ->3	
ryk.	H->1	
ryka	 ->23	,->2	s->4	
ryke	r->2	
ryks	 ->2	
rykt	a->1	b->1	e->7	
rymd	 ->1	e->1	
rymm	a->1	e->11	
ryms	 ->1	
rymt	 ->1	
ryos	t->1	
ryph	å->3	
ryps	.->1	
rypt	o->2	
ryr 	e->1	j->1	
rys 	o->1	
rysa	 ->2	
rysk	 ->1	a->1	
rysn	i->1	
ryss	a->2	e->19	
ryta	 ->6	n->1	s->1	
ryte	l->2	r->7	
rytn	i->2	
rytt	e->2	
rzwa	l->1	
rä u	t->1	
rä ö	v->1	
räck	 ->1	a->13	e->22	h->1	l->77	n->31	s->2	t->3	v->3	
räd 	b->1	f->1	h->2	u->1	
räd,	 ->1	
räd.	D->1	
räda	 ->10	,->1	n->10	r->57	
rädd	 ->5	,->1	a->14	e->7	n->4	
räde	 ->15	.->3	H->1	P->1	l->5	n->4	r->16	s->9	t->12	
räds	 ->2	l->9	
räff	a->115	l->2	
räft	a->29	e->1	
räga	r->1	
räge	r->36	
rägl	a->5	i->1	
räke	n->9	
räkn	a->39	e->2	i->14	
räkt	a->1	s->1	
räl 	g->1	i->1	
räl,	 ->1	
rämb	e->1	
rämd	 ->1	
räme	l->1	
rämj	a->62	
räml	i->35	
rämm	a->3	e->2	
räms	t->48	
rän 	m->2	n->1	s->1	å->2	
räna	 ->3	
ränd	a->2	e->4	r->73	
räng	 ->4	a->18	d->2	e->5	n->35	t->5	
räni	n->1	t->12	
ränk	a->2	b->1	e->5	n->13	s->3	t->7	
ränn	a->3	i->2	
räns	 ->2	a->62	e->34	f->2	k->7	l->7	n->12	o->1	p->1	v->1	ö->12	
ränt	a->1	
räpn	i->1	
räpr	o->1	
rär 	o->1	
rärt	 ->1	
räsc	h->2	
räsk	.->1	
räta	s->1	
räto	r->1	
rätt	 ->112	,->10	.->7	?->2	a->114	e->90	f->8	h->9	i->122	m->1	n->2	s->204	v->72	ä->1	
räva	 ->33	d->4	n->17	r->4	s->9	t->1	
rävd	e->4	
räve	r->45	
rävi	g->1	
rävs	 ->52	,->3	
rävt	 ->1	s->1	
rå s	o->1	
rå v	a->1	
rå ä	r->1	
råd 	(->1	-->1	a->1	b->1	f->3	i->1	n->1	o->5	s->3	
råd,	 ->4	
råd.	D->1	J->1	K->1	L->1	M->1	
råd?	Ä->1	
råda	 ->9	n->4	r->3	
rådd	e->1	
råde	 ->57	,->14	.->23	:->1	;->1	?->1	n->134	r->24	t->396	
rådf	r->6	
rådg	i->26	ö->1	
råds	b->1	k->20	l->3	m->3	o->19	r->1	t->1	
råer	,->1	
rået	.->1	
råga	 ->232	!->1	,->24	.->40	:->7	?->1	d->8	n->203	r->20	s->20	t->6	v->1	
råge	k->1	s->10	t->2	
rågn	i->8	
rågo	r->275	
råk 	f->1	p->3	t->1	
råk.	 ->1	
råka	 ->1	r->9	
råke	t->4	
råki	g->3	
råkl	i->3	
råko	m->2	
råkr	a->30	
råkt	a->1	
råld	r->3	
rålk	a->1	
råln	i->3	
råls	k->1	
rån 	(->21	-->1	1->7	2->1	3->1	5->3	8->1	9->1	A->10	B->5	C->3	D->2	E->29	F->6	G->4	H->2	I->5	J->1	K->5	L->3	M->1	N->3	O->1	P->7	R->1	S->6	T->6	U->2	V->1	W->2	a->35	b->13	d->94	e->43	f->33	g->4	h->6	i->1	j->4	k->37	l->8	m->21	n->6	o->22	p->18	r->17	s->25	t->25	u->22	v->19	Ö->1	ä->1	å->1	ö->4	
rån,	 ->3	
rån.	D->1	Ä->1	
rång	 ->1	,->2	e->1	l->1	m->1	å->1	
rånk	o->3	
rånt	a->2	o->1	
rånv	a->8	ä->1	
råol	j->1	
råps	l->1	
råri	g->12	
rås 	f->2	
råt 	k->1	
råtg	ä->1	
rått	o->1	
råzo	n->1	
rébe	t->1	
réfé	r->1	
rêts	 ->1	
rínc	i->1	
rón 	C->2	i->1	t->1	v->1	
röd.	-->1	D->2	
röda	 ->2	n->3	
röde	l->2	r->1	
rödg	r->1	
rödo	r->1	
rögh	e->1	
röja	 ->5	.->1	r->1	s->1	
röjd	e->1	
röje	r->3	
röjo	r->1	
röjs	m->2	
röjt	s->1	
rök 	b->1	
rök,	 ->1	
röks	,->1	
röm 	a->2	b->1	i->1	
röm,	 ->1	
röm:	 ->1	
römm	a->4	e->4	
römn	i->6	
römt	 ->1	
römv	ä->1	
rön 	v->2	
röna	 ->12	/->1	r->1	s->2	
rönb	o->1	
röni	t->1	
rönt	 ->1	
rör 	E->1	P->1	a->3	b->1	d->6	f->6	i->1	j->1	k->1	o->3	p->3	s->17	t->2	u->3	v->1	
röra	 ->3	n->24	s->2	
rörd	 ->2	a->19	e->2	h->1	
röre	l->9	
röri	g->2	
rörl	i->24	
rörs	 ->8	
rört	 ->3	s->2	
rös 	o->1	p->1	r->1	
rösa	 ->3	
rösk	e->3	
röst	 ->13	,->2	.->2	a->90	e->5	f->7	n->57	r->3	t->1	v->3	
röt 	h->1	t->4	
röts	 ->2	
rött	 ->1	.->1	a->2	e->4	
röva	 ->4	d->1	r->4	s->4	t->1	
röve	r->1	
rövn	i->5	
rövo	å->1	
rövr	a->2	
rövs	t->1	
s "B	i->1	
s "g	e->1	
s (P	P->1	
s (f	i->1	
s (u	n->1	
s - 	a->2	b->1	e->1	f->1	h->1	i->2	j->1	m->1	n->1	o->7	s->1	t->1	
s -,	 ->1	
s 19	5->1	6->1	9->3	
s 2 	4->1	
s 20	 ->1	0->1	
s 24	 ->1	
s 28	:->1	
s 3,	8->1	
s 40	0->1	
s 80	 ->1	
s Ad	o->1	
s Al	g->1	
s BN	I->2	P->1	
s Ba	l->1	r->2	
s Bl	o->1	
s CE	N->1	
s Da	m->1	
s De	l->3	
s EG	-->2	
s EU	-->2	
s Eu	r->13	
s FP	Ö->1	
s Ge	n->1	
s Gi	l->1	
s Go	l->1	
s He	l->1	
s Is	r->1	
s Le	i->1	
s Mi	t->1	
s Oz	,->1	
s Pa	c->1	
s RE	P->1	
s Ru	i->1	
s SO	L->1	
s Sj	ö->2	
s Sp	a->3	
s VD	 ->1	
s Vi	c->1	
s Wi	e->1	
s Wu	r->1	
s XX	V->1	
s ab	s->3	
s ad	m->1	
s ag	e->3	
s ak	t->1	
s al	b->1	d->1	k->1	l->44	t->1	
s am	b->3	
s an	 ->3	a->3	d->11	f->2	g->5	h->1	i->1	l->2	m->4	n->1	p->1	s->57	t->5	v->3	
s ar	b->36	g->2	k->1	t->2	
s at	t->174	
s au	k->3	t->1	
s av	 ->272	d->1	g->6	s->7	t->1	v->1	
s ax	l->1	
s ba	c->1	k->1	r->4	s->2	
s be	f->12	g->12	h->14	k->2	l->1	n->1	r->3	s->36	t->59	v->3	
s bi	d->4	l->4	s->1	
s bl	.->2	a->4	i->7	o->2	
s bo	r->8	
s br	a->2	i->4	u->1	y->1	å->1	
s bu	d->15	
s by	g->1	r->3	
s bä	r->1	s->3	t->3	
s bå	d->4	
s bö	r->1	
s ce	n->7	
s ci	r->1	
s co	s->1	
s da	 ->5	g->16	t->1	
s de	 ->24	b->7	f->3	l->24	m->13	n->27	r->2	s->3	t->101	
s di	m->2	p->2	r->18	s->3	t->1	
s dj	u->1	
s do	c->2	g->1	k->4	m->6	
s dr	a->2	
s du	 ->1	b->1	
s dä	r->31	
s då	 ->3	
s dö	d->5	
s ef	f->6	t->18	
s eg	e->12	n->6	
s ek	o->30	
s el	l->23	
s em	b->1	e->5	o->2	
s en	 ->94	d->9	e->2	h->9	l->6	o->1	s->2	v->1	
s er	f->2	s->1	
s et	 ->1	t->42	
s eu	r->3	
s ev	e->1	
s ex	a->1	e->3	i->3	k->1	p->2	t->2	
s fa	b->1	k->4	l->5	m->3	n->1	r->6	s->4	v->1	
s fe	l->2	m->2	
s fi	l->1	n->6	s->4	
s fj	o->1	
s fl	a->5	e->9	o->1	y->1	
s fo	l->6	n->2	r->17	t->2	
s fr	a->55	e->2	i->9	ä->5	å->42	
s fu	l->13	n->8	
s fy	l->1	r->2	s->1	
s få	 ->8	r->2	
s fö	l->4	r->298	
s ga	l->1	n->1	r->3	s->1	
s ge	 ->1	m->26	n->36	o->1	r->1	
s gi	l->4	v->1	
s gj	o->1	
s go	d->8	
s gr	a->4	u->21	ä->5	ö->1	
s gu	v->1	
s gä	l->1	r->2	
s gå	 ->1	n->2	r->1	
s gö	r->4	
s ha	 ->3	d->4	f->1	m->4	n->9	r->33	v->5	
s he	k->1	l->4	t->1	
s hi	n->1	s->7	t->4	
s hj	ä->5	
s ho	p->2	s->3	t->1	
s hu	r->3	v->4	
s hy	c->1	
s hä	l->8	n->6	r->20	
s hå	l->2	r->5	
s hö	g->2	j->1	
s i 	2->1	A->4	B->2	D->1	E->12	F->3	G->2	I->1	J->1	K->5	L->2	M->3	P->1	S->8	T->3	U->1	a->8	b->9	d->56	e->19	f->27	g->6	h->9	j->1	k->9	l->2	m->7	n->5	o->6	p->12	r->18	s->24	t->5	u->2	v->16	Ö->1	ä->3	å->1	ö->3	
s id	e->2	é->2	
s ig	e->4	
s ih	o->1	
s ik	r->2	
s il	l->2	
s im	m->1	
s in	 ->8	,->3	b->2	d->3	f->5	g->29	i->6	k->4	l->4	n->15	o->15	r->12	s->28	t->88	v->3	
s ir	r->1	
s ja	g->11	
s jo	r->2	
s ju	 ->2	d->1	r->11	s->5	v->1	
s jä	m->1	
s ka	b->1	l->3	n->10	p->3	t->1	
s ke	m->1	
s kl	.->6	a->6	i->1	
s ko	l->4	m->42	n->41	p->1	r->5	
s kr	a->8	e->1	i->3	ä->1	
s ku	l->4	m->2	n->3	s->5	
s kv	a->10	i->1	o->1	
s kä	l->1	n->2	r->2	
s kö	p->1	
s la	g->18	n->7	
s le	 ->1	d->15	g->7	t->1	v->3	
s li	b->2	g->1	k->12	l->1	n->1	t->1	v->10	
s lj	u->1	
s lo	b->1	g->2	p->2	v->1	
s lu	c->1	g->1	
s lä	g->2	m->2	n->6	r->1	s->1	
s lå	n->1	
s lö	f->2	p->1	
s ma	k->5	n->6	r->2	s->1	t->1	
s me	d->168	l->15	n->4	r->7	s->3	t->3	
s mi	g->1	l->12	n->10	s->1	
s mo	n->2	r->1	t->18	
s my	c->17	
s mä	n->4	r->2	
s må	l->12	n->20	s->9	
s mö	j->15	r->1	t->3	
s na	c->2	m->6	t->16	
s ne	d->5	g->4	
s ni	 ->2	o->1	v->4	
s no	g->1	r->1	
s nu	 ->7	v->9	
s ny	a->6	f->1	l->4	s->1	
s nä	m->4	r->17	s->1	
s nå	g->33	
s nö	d->3	
s oa	c->1	n->2	
s ob	e->3	l->3	
s oc	h->189	k->39	
s od	i->1	j->1	
s oe	n->1	
s of	f->5	t->2	ö->3	
s oh	j->1	ö->1	
s oi	n->5	
s ok	u->1	
s ol	a->1	i->6	j->1	y->1	ä->1	
s om	 ->70	)->1	,->1	.->6	b->1	f->5	r->7	s->1	v->1	
s or	d->40	g->5	i->1	o->10	s->1	
s os	s->3	ä->2	
s ot	i->3	r->1	v->1	
s ov	a->1	
s pa	p->1	r->22	s->1	t->1	
s pe	l->1	n->3	r->6	
s ph	a->1	
s pl	a->5	e->1	
s po	l->24	p->1	r->3	s->4	t->1	ä->1	
s pr	a->1	e->7	i->13	o->20	
s pu	b->1	n->1	
s på	 ->157	,->1	.->1	p->3	t->1	
s qu	o->2	
s ra	d->1	m->3	n->1	p->15	s->3	t->1	
s re	a->2	d->7	f->5	g->40	k->3	l->1	p->1	s->23	t->1	
s ri	g->1	k->8	s->4	
s ro	,->1	c->1	l->10	t->1	
s ru	n->3	t->1	
s ry	k->2	
s rä	d->1	k->10	t->40	
s rå	d->4	
s rö	r->3	s->2	t->1	
s sa	d->3	k->7	m->35	t->1	
s sc	i->1	
s se	 ->3	d->4	g->1	k->3	m->1	n->2	r->1	s->2	x->1	
s si	d->26	f->1	k->1	n->4	s->1	t->7	
s sj	ä->15	
s sk	a->21	e->1	i->3	o->5	r->2	u->24	y->3	ä->3	ö->3	
s sl	a->4	o->2	u->13	
s sm	å->2	
s sn	a->6	
s so	c->12	l->3	m->107	
s sp	e->9	å->1	ö->1	
s st	a->10	e->2	o->4	r->30	u->2	y->2	ä->9	å->14	ö->17	
s su	b->2	v->6	
s sv	a->5	å->5	
s sy	f->2	n->8	
s sä	g->2	k->10	l->1	n->1	r->8	t->4	
s så	 ->17	d->1	l->4	r->1	v->1	
s sö	n->2	
s ta	 ->3	c->1	k->2	l->6	n->2	p->1	
s te	k->2	n->2	r->5	x->4	
s ti	d->13	l->142	o->2	
s tj	o->1	u->1	ä->11	
s to	g->1	t->2	
s tr	a->2	e->4	o->13	
s tu	l->1	r->3	
s tv	i->5	ä->2	å->5	
s ty	d->6	p->3	v->1	
s un	d->43	i->1	
s up	p->71	
s ur	 ->2	s->6	
s ut	 ->12	,->4	.->5	a->10	b->3	f->7	g->4	i->3	m->7	n->1	r->5	s->7	t->25	v->23	ö->1	
s va	c->1	d->5	l->3	n->1	p->2	r->30	t->3	
s ve	c->1	r->29	t->2	
s vi	 ->9	a->1	c->1	d->23	k->9	l->17	n->1	s->6	t->5	
s vo	l->1	t->1	
s vu	x->1	
s vä	c->2	g->22	k->1	l->4	n->3	p->1	r->7	s->1	
s vå	n->1	r->3	
s yr	k->2	
s yt	a->1	t->18	
s äg	a->6	g->1	
s än	 ->2	d->12	n->7	
s är	 ->50	
s äv	e->7	
s ål	d->5	
s år	 ->2	.->1	h->1	l->4	
s ås	i->8	t->3	
s åt	 ->17	,->1	.->1	a->2	e->5	g->10	m->2	
s öd	e->5	
s ög	o->2	
s ök	a->5	
s öm	s->1	t->1	
s ön	s->2	
s öp	p->2	
s ör	e->2	o->1	
s öv	e->37	r->1	
s! J	a->1	
s! V	a->1	
s!De	t->1	
s!Eu	r->1	
s!Fö	r->1	
s!Ge	n->1	
s!He	r->1	
s!Vi	 ->1	
s".D	e->1	
s".J	a->1	
s".K	a->1	
s) f	ö->1	
s) o	c->1	
s, 1	2->1	
s, E	v->1	
s, L	u->1	
s, M	i->1	
s, S	t->1	
s, T	o->1	
s, W	u->1	
s, a	l->2	n->3	t->12	v->1	
s, b	e->3	l->1	ä->1	ö->1	
s, d	e->7	i->1	v->1	ä->4	å->3	
s, e	f->8	l->2	n->6	t->3	u->1	
s, f	o->1	r->7	ö->15	
s, g	e->2	i->1	ö->1	
s, h	a->3	e->2	u->2	ä->1	
s, i	 ->6	n->8	
s, j	a->3	o->1	
s, k	a->1	o->6	
s, l	e->1	
s, m	e->25	i->2	o->1	y->1	ä->2	å->1	
s, n	ä->7	å->2	
s, o	c->44	m->8	
s, p	a->1	å->6	
s, r	e->1	
s, s	a->1	k->2	o->10	p->2	ä->2	å->15	
s, t	.->1	i->1	r->3	y->1	
s, u	n->1	p->1	r->1	t->8	
s, v	a->4	i->9	ä->1	å->1	
s, ä	r->4	v->2	
s, å	t->4	
s- f	ö->1	
s- o	c->42	
s-, 	u->1	
s-Ca	r->1	
s-Jø	r->2	
s-be	l->1	s->1	
s-bi	l->1	
s-de	-->1	
s-fö	r->1	
s-in	t->2	
s-no	t->1	
s-ny	t->1	
s-pr	o->1	
s-si	t->1	
s. 1	1->2	
s. D	e->3	
s. E	q->1	u->1	
s. M	e->2	
s. P	a->1	
s. W	a->1	
s. a	r->1	t->10	
s. d	e->4	
s. e	n->1	r->1	t->1	
s. f	o->1	ö->2	
s. g	r->1	
s. h	o->1	u->1	
s. i	 ->1	d->1	n->3	
s. j	a->1	
s. m	a->2	e->1	i->1	
s. n	ä->1	
s. o	m->2	
s. p	å->1	
s. s	p->1	
s. v	a->1	i->1	
s.(E	N->1	
s.)Å	t->1	
s.- 	(->1	
s..(	F->1	
s.Al	l->3	
s.An	h->1	t->1	
s.At	t->1	
s.Be	t->3	v->1	
s.Bl	a->2	
s.Ce	n->1	
s.Da	g->1	
s.De	 ->4	n->15	s->2	t->62	
s.Di	r->1	
s.Dä	r->12	
s.Då	 ->4	
s.Ef	t->2	
s.Ek	o->1	
s.En	 ->5	d->1	l->2	
s.Er	t->1	
s.Et	t->5	
s.Eu	r->3	
s.Fa	c->1	
s.Fl	o->2	
s.Fr	u->5	å->2	
s.Fö	r->8	
s.Ge	n->4	
s.Gr	e->1	
s.Ha	n->1	
s.He	l->1	r->10	
s.Hi	s->1	t->1	
s.Ho	p->1	
s.Hu	r->1	v->1	
s.Hä	r->1	
s.I 	a->2	d->3	e->1	k->1	l->1	r->1	s->2	ö->1	
s.In	g->1	o->1	t->1	
s.Ja	g->28	
s.Jo	n->1	
s.Ju	s->1	
s.Jä	m->1	
s.Ko	m->6	n->1	s->1	
s.La	n->1	
s.Le	d->1	
s.Lå	t->2	
s.Ma	n->3	
s.Me	d->3	l->1	n->9	
s.Mi	n->2	
s.My	n->1	
s.Mä	n->1	
s.Må	n->1	
s.Ni	 ->1	
s.Nu	 ->2	
s.Nä	r->4	
s.Nå	g->1	
s.OL	A->1	
s.Oa	v->1	
s.Om	 ->2	
s.On	ö->1	
s.Pa	r->3	
s.Pe	r->1	
s.Pr	e->1	o->1	
s.På	 ->2	
s.Ra	p->1	
s.Re	a->1	d->1	s->2	
s.Rå	d->1	
s.Sa	m->2	n->1	
s.Se	d->1	
s.Sl	u->5	
s.Sn	a->1	
s.So	m->2	
s.Så	 ->1	
s.Ta	c->1	l->1	n->1	
s.Ti	l->1	
s.Ty	v->1	
s.Un	d->4	
s.Ut	f->1	m->1	
s.Va	d->4	r->2	
s.Vi	 ->29	d->1	l->1	
s.Vå	r->3	
s.Yt	t->2	
s.k.	 ->4	
s.Än	d->2	n->1	
s.Äv	e->2	
s.Åt	a->1	g->1	
s/de	n->1	
s/in	t->1	
s: a	n->1	t->1	
s: e	n->1	
s: f	ö->1	
s: h	ö->1	
s: k	o->1	
s: v	a->1	
s; a	t->1	
s; b	)->1	
s; d	e->1	
s; e	n->1	
s; o	c->1	
s; v	i->1	
s?. 	(->1	
s?.H	e->1	
s?De	n->1	
s?Et	t->1	
s?Fr	å->1	
s?Ha	r->1	
s?I 	s->1	
s?Ja	,->1	
s?Jo	,->1	
s?Ko	m->1	
s?Oc	h->1	
s?Sk	u->1	
s?Ti	l->1	
s?Vi	l->2	
s?Är	 ->1	
sNäs	t->1	
sa (	a->1	
sa -	 ->1	
sa 1	0->1	
sa 2	5->3	
sa 3	5->1	
sa P	P->1	
sa R	y->1	
sa a	l->4	m->1	n->14	r->5	s->2	t->7	v->23	
sa b	e->14	i->5	l->2	r->3	å->4	ö->1	
sa c	e->1	
sa d	a->1	e->23	i->1	o->2	r->1	
sa e	f->2	g->1	l->1	n->3	r->2	
sa f	a->11	e->1	i->2	o->6	r->23	u->1	ö->22	
sa g	a->1	e->6	o->2	r->6	
sa h	a->4	e->1	i->7	o->1	u->2	ä->2	ö->1	
sa i	 ->11	n->20	
sa k	a->7	l->1	o->16	r->4	u->1	v->3	
sa l	a->3	i->1	ä->13	ö->2	
sa m	a->4	e->17	i->8	o->3	ä->1	å->13	ö->2	
sa n	i->2	o->1	y->1	å->1	
sa o	b->1	c->18	k->1	l->1	m->21	r->4	s->1	
sa p	a->5	e->10	i->1	l->3	o->1	r->22	u->5	å->14	
sa r	e->22	i->9	u->1	ä->1	
sa s	.->1	a->8	e->2	i->13	j->1	k->8	l->2	m->2	o->4	p->5	t->13	v->1	y->1	ä->3	å->1	
sa t	a->2	e->2	i->15	o->2	r->8	v->4	y->1	
sa u	n->5	p->11	r->1	t->5	
sa v	a->7	e->2	i->6	ä->8	å->2	
sa ä	m->2	n->26	r->7	v->1	
sa å	r->1	t->8	
sa ö	v->3	
sa!L	å->1	
sa, 	5->1	b->1	d->3	e->1	f->5	g->1	h->1	l->1	m->2	o->1	s->2	u->1	v->1	å->1	
sa..	.->1	
sa.A	n->1	
sa.B	a->1	l->1	
sa.D	e->4	ä->2	
sa.E	u->1	
sa.F	r->1	ö->1	
sa.H	e->1	
sa.I	 ->2	
sa.J	a->3	
sa.K	ä->1	
sa.M	a->1	e->2	i->1	
sa.R	å->1	
sa.S	a->1	
sa.U	p->1	
sa.Å	r->1	
sa?P	r->1	
sabe	l->2	t->1	
sabl	a->1	
sabo	n->8	
saca	 ->1	
sace	 ->1	.->2	
sad 	a->1	d->2	e->2	g->1	h->1	o->3	s->2	t->6	
sad,	 ->2	
sad.	D->1	J->1	V->1	
sade	 ->84	,->14	.->6	:->1	s->3	
sadö	r->1	
safe	t->1	
saff	ä->2	
saft	o->1	
sag 	i->1	
sage	r->1	
sagt	 ->28	,->8	.->1	s->12	
sail	l->1	
sak 	a->4	b->2	g->3	h->3	j->1	k->1	m->4	n->1	s->9	t->3	u->1	v->5	ä->2	
sak,	 ->2	
sak.	A->1	D->1	E->1	N->1	T->1	
sak:	 ->1	
saka	 ->5	d->3	r->4	s->2	t->6	
sake	n->15	r->45	
sakf	ö->1	
sakk	u->2	
sakl	i->11	
sakn	a->39	
sako	m->2	
sakp	r->1	
sakr	e->1	
sakt	 ->2	.->1	e->3	i->2	ö->1	
sala	 ->1	
sale	m->2	
sali	n->1	
salm	e->1	
salt	e->1	
salu	f->1	
sam 	a->4	b->3	c->1	d->5	e->3	f->4	g->1	h->2	i->2	l->2	m->6	n->1	o->3	p->5	r->6	s->10	t->3	u->2	v->3	å->2	ö->2	
sam,	 ->2	
sam.	I->1	
sama	r->83	
samb	a->47	
same	x->2	
samf	i->1	u->5	ö->7	
samh	e->97	ä->47	
samk	a->3	
saml	a->20	e->1	i->25	
samm	a->492	e->1	
samo	r->37	
samr	ä->1	å->9	
sams	t->4	y->3	
samt	 ->99	,->2	.->3	a->16	i->53	l->25	y->6	
samv	e->5	
san 	h->1	i->2	o->2	t->1	ä->1	
san,	 ->2	
san.	M->1	S->1	V->1	
sana	l->6	
sand	a->4	e->16	
sanf	ö->1	
sank	t->8	
sanl	ä->9	
sanm	ä->1	
sann	 ->1	a->1	e->4	i->3	o->8	
sans	 ->1	a->2	p->1	t->1	v->1	
sant	 ->24	!->1	,->3	.->2	:->1	a->5	
sar 	a->10	d->6	e->6	f->3	h->2	i->5	j->2	k->3	m->3	n->2	o->6	p->9	r->2	s->5	t->9	u->2	v->8	ä->3	å->1	
sar!	D->1	
sar,	 ->4	
sar.	D->1	S->1	
sarb	e->27	
sare	 ->4	.->1	
sarg	u->1	
sarn	a->1	
sart	i->3	
sas 	a->1	b->2	d->2	e->1	i->3	k->1	m->2	o->4	p->1	s->3	t->10	v->1	
sas,	 ->1	
sas.	D->1	
sasp	e->3	
sat 	a->10	b->1	d->2	e->5	f->1	h->1	i->2	m->2	n->1	o->2	p->4	s->9	t->1	v->1	
sat,	 ->1	
sat.	D->2	F->1	H->1	N->1	
sate	l->1	
sati	o->46	
sato	r->3	
sats	 ->24	,->5	.->3	a->13	e->85	f->1	n->4	o->3	s->3	
satt	 ->21	,->3	.->2	a->27	e->9	s->3	
saur	o->1	
savb	r->1	
savg	i->1	r->1	å->1	ö->5	
savi	 ->1	
savt	a->15	
savv	e->1	
sban	k->2	
sbar	 ->1	a->1	t->3	
sbas	.->1	e->1	
sbed	r->2	ö->2	
sbef	o->3	r->6	
sbeg	r->4	
sbeh	a->3	o->1	
sbek	ä->3	
sbel	a->4	o->2	ä->1	
sber	ä->2	
sbes	k->2	l->7	t->23	ä->1	
sbet	a->2	o->1	ä->2	
sbev	a->1	i->6	
sbid	r->2	
sbil	d->7	
sbis	t->2	
sbol	a->3	
sbor	d->3	
sbou	r->5	
sbri	s->2	
sbro	t->2	
sbru	k->16	
sbud	g->3	
sbur	n->1	
sbus	s->1	
sbut	i->1	
sbyg	d->43	g->1	
sbåd	a->1	
sbör	d->12	
scay	a->6	
scen	 ->1	a->5	e->1	s->1	t->7	
scer	t->1	
sch 	f->1	i->1	o->1	s->1	
sch!	 ->1	
sch.	E->1	
sch?	F->1	
scha	b->1	
sche	 ->1	f->12	m->1	n->5	r->4	
schh	o->1	
schl	e->4	
schw	i->1	
scie	n->1	
scip	l->14	
scis	m->3	t->9	
scor	e->1	
scyk	e->3	
sdag	 ->8	.->4	:->1	e->1	s->1	
sdeb	a->3	
sdel	 ->4	.->1	a->8	e->1	
sdep	a->1	
sdig	r->2	
sdik	t->5	
sdim	e->1	
sdir	e->7	
sdok	u->6	
sdom	 ->1	i->1	s->2	
sdra	b->4	
sdrä	n->1	
sdug	l->5	
sduk	a->1	
sdöm	d->1	t->1	
se (	a->1	
se -	 ->3	
se G	r->1	
se a	n->1	r->1	t->38	v->14	
se b	a->1	e->1	
se d	e->16	o->1	
se e	l->1	n->3	t->3	
se f	o->1	r->10	ö->22	
se g	e->2	i->1	
se h	a->3	o->2	u->4	ä->1	
se i	 ->9	n->2	
se j	a->2	u->1	
se k	a->2	o->5	
se l	y->1	
se m	e->20	o->1	y->1	
se n	o->2	ä->3	
se o	c->15	l->1	m->13	
se p	e->1	å->11	
se r	e->2	i->1	
se s	a->2	i->1	k->2	n->2	o->17	p->1	t->1	ä->1	å->1	
se t	a->1	i->70	
se u	n->1	p->2	t->3	
se v	a->4	e->1	i->10	
se ä	n->1	r->3	
se ö	v->14	
se",	 ->1	
se, 	d->3	e->3	i->3	j->1	k->1	l->1	m->3	s->1	t->1	u->1	v->1	
se- 	o->1	
se-N	o->1	
se.B	e->1	
se.D	e->6	
se.E	f->1	n->2	t->1	
se.F	ö->1	
se.J	a->3	
se.K	o->1	
se.L	å->1	
se.M	a->1	e->1	i->2	
se.N	i->1	
se.O	m->1	
se.S	a->1	k->1	
se.V	a->1	i->2	
se; 	j->1	
se?E	n->1	
seak	t->1	
seba	l->1	
seby	g->1	
sed 	s->1	
seda	n->104	
sedd	 ->2	a->3	
sede	r->1	
seen	d->60	
seff	e->7	
sefu	l->11	
seg 	t->1	
segd	r->1	
sege	r->4	
segl	a->13	
segr	a->3	
sehi	n->1	
seil	l->1	
seis	m->2	
seke	l->4	
sekl	e->2	
seko	n->26	
sekr	e->16	
sekt	i->2	o->89	
seku	n->3	
sekv	e->61	
sel 	f->2	i->1	k->2	m->1	n->1	o->5	v->1	ä->1	å->1	
sel!	 ->1	T->1	
sel,	 ->5	
sel-	 ->1	I->2	
sel.	D->1	F->1	S->1	
selb	y->1	
sele	d->2	k->1	
self	e->1	
sell	 ->2	a->1	
selo	d->1	
sels	a->1	ä->102	
selö	s->3	
seme	l->3	s->4	
semi	n->1	t->3	
semö	n->1	
sen 	"->1	(->2	-->6	1->2	2->1	E->2	M->1	a->49	b->10	d->6	e->2	f->16	g->3	h->10	i->39	k->7	l->3	m->23	n->3	o->26	p->5	r->1	s->32	t->11	u->6	v->7	ä->10	ö->1	
sen!	N->1	
sen,	 ->44	
sen.	 ->3	A->4	D->17	E->1	F->4	G->1	H->7	I->3	J->9	K->1	L->1	M->3	N->2	O->4	P->1	R->2	S->5	T->1	V->14	Ä->1	
sen;	 ->1	
sen?	F->2	
senN	ä->2	
sena	 ->6	,->1	d->10	r->30	s->68	t->1	
senb	e->3	
send	e->9	
senf	ä->1	
senh	e->4	
seni	n->13	
senl	i->3	
senr	ö->1	
sens	 ->29	,->1	i->1	
sent	 ->3	,->1	.->4	a->33	e->24	l->26	
seom	r->1	
sepa	r->1	
sept	e->15	
ser 	-->4	4->1	A->1	E->1	a->132	b->7	d->34	e->12	f->59	g->3	h->9	i->30	j->38	k->11	l->1	m->13	n->5	o->46	p->10	r->5	s->53	t->16	u->12	v->31	ä->5	å->1	ö->4	
ser!	D->1	
ser,	 ->40	
ser.	 ->2	(->1	-->1	.->1	9->1	A->1	B->1	D->11	E->1	F->1	H->2	I->4	J->3	K->5	O->1	S->1	T->1	V->5	
ser:	 ->1	
ser?	E->1	M->1	V->1	
sera	 ->59	.->1	d->43	n->3	r->23	s->19	t->15	
serb	,->1	e->7	i->6	j->1	
seri	 ->2	.->1	e->1	k->1	n->90	ö->7	
serl	i->13	
sern	a->140	
sers	 ->1	
serv	a->11	e->4	i->7	t->1	
ses 	d->2	f->1	g->1	i->1	m->3	p->1	s->4	t->1	u->1	v->2	ö->5	
ses.	A->1	
sesi	d->5	
sess	i->6	
set 	-->2	a->6	b->2	e->2	f->6	h->1	i->4	k->2	m->2	o->1	p->3	u->1	
set,	 ->1	
set.	D->1	F->1	J->1	
seta	p->1	
seti	k->1	
sets	 ->1	
sett	 ->58	,->3	.->5	:->1	s->2	
setê	t->2	
seur	o->1	
seut	v->1	
sevi	s->2	
sevä	r->14	
sewi	e->1	
sex 	a->2	e->1	m->11	p->1	t->1	ö->1	
sex,	 ->1	
sexi	s->1	
sexm	å->1	
sexp	o->1	
sext	o->1	
sexu	e->3	
sexv	ä->1	
sfak	t->1	
sfal	l->6	
sfar	a->2	
sfas	,->1	e->4	t->1	
sfat	t->11	
sfel	,->1	e->1	
sfie	n->31	
sfin	a->1	
sfis	k->3	
sfla	g->15	
sflo	t->2	
sfly	g->1	
sfon	d->22	
sfor	d->1	m->4	s->1	u->2	
sfos	t->1	
sfri	 ->3	a->2	h->45	s->10	
sfrä	m->4	
sfrå	g->44	n->1	
sful	l->16	
sfun	k->2	
sfär	e->1	
sfäs	t->1	
sfån	g->1	
sför	b->1	d->13	e->5	f->16	h->20	k->5	l->2	m->8	o->3	s->219	
sgar	a->3	
sgas	e->4	
sgem	e->1	
sgil	l->1	
sgiv	a->15	n->1	
sgra	d->5	
sgre	n->2	
sgru	n->1	p->10	
sgrä	n->3	
sgyn	n->7	
sgå 	K->1	d->1	
sgås	:->1	
sgör	 ->1	
sh P	e->1	o->1	
sh, 	a->1	
shal	l->1	
shan	d->13	t->2	
shat	e->1	
shau	s->1	
shav	e->1	
shem	 ->1	
sher	r->1	
shet	 ->15	,->4	.->4	e->25	s->3	
shin	d->11	g->3	
ship	 ->1	
shjä	l->2	
shop	,->1	
shot	a->1	
shus	.->1	h->1	
shäm	m->2	
shän	s->1	
shål	l->1	
sias	m->3	
siat	i->2	
sibi	l->1	
sida	 ->13	,->9	.->8	?->1	n->46	r->1	
side	n->9	s->2	
sidi	a->21	g->13	ä->1	
sidk	a->1	
sido	e->1	r->6	
sidu	e->1	
siel	l->37	
sien	 ->4	,->1	.->1	s->1	
sier	a->16	i->34	
siff	r->22	
sifi	c->9	e->5	
sifu	l->1	
sig 	E->1	O->1	a->44	b->12	d->14	e->18	f->36	g->4	h->4	i->39	j->1	k->3	l->2	m->27	n->7	o->34	p->27	r->2	s->25	t->26	u->9	v->11	ä->5	å->13	ö->4	
sig,	 ->8	
sig.	A->1	B->1	D->2	E->2	H->2	J->2	K->1	M->1	S->1	T->1	V->3	Ä->1	
sig;	 ->1	
siga	 ->14	,->2	
sign	a->14	e->2	
sigt	 ->13	.->1	
sik 	i->1	m->1	
sike	.->1	n->1	r->1	
sikt	 ->69	,->9	.->6	a->2	e->48	i->76	l->4	n->2	s->3	
sil 	e->1	
sila	 ->2	
sili	e->1	
silv	e->3	
simi	s->2	
simm	a->1	
simu	l->2	
sin 	a->5	b->10	d->6	e->14	f->12	g->2	h->19	i->4	k->3	l->3	m->6	n->8	o->7	p->9	r->17	s->19	t->6	u->9	v->5	w->1	ä->1	å->2	ö->1	
sin.	B->1	
sina	 ->138	
sind	u->8	
sine	 ->3	
sinf	o->2	r->1	
sing	f->20	
sini	t->9	
sinn	a->1	e->6	i->1	
sino	m->1	
sinr	i->4	
sins	a->4	e->3	p->2	t->13	
sint	e->3	r->1	
sion	 ->51	)->2	,->4	.->10	?->3	e->937	s->44	ä->248	
sis 	a->2	n->1	o->1	
sis,	 ->1	
sisk	 ->6	,->1	a->83	e->2	t->6	
sism	 ->6	,->2	.->4	e->3	
sist	 ->8	,->4	.->1	a->44	e->7	i->11	n->2	
site	t->1	
siti	o->15	v->75	
sitl	a->2	ä->1	
sitr	u->1	
sitt	 ->94	,->1	a->1	e->8	n->2	r->1	
situ	a->126	
siv 	a->1	b->1	k->1	m->1	r->1	s->2	t->1	
siv.	.->1	
siva	 ->7	r->1	
sive	 ->17	
sivt	 ->11	
siär	a->1	e->1	
sjov	i->17	
sju 	g->1	i->1	m->1	p->1	r->1	
sju,	 ->1	
sjuk	.->1	a->1	d->1	f->1	h->6	v->3	
sjun	d->4	k->9	
sjur	i->2	
sjut	t->2	
själ	,->1	.->2	e->2	v->168	
sjät	t->19	
sjöf	a->8	
sjöm	ä->2	
sjön	.->1	k->4	
sjös	s->4	
sjöt	r->1	
sjöv	ä->1	
sk -	 ->1	
sk T	V->1	
sk a	 ->1	g->1	l->7	n->5	r->3	s->1	t->2	
sk b	a->4	e->7	i->4	l->1	o->1	r->1	y->2	ö->1	
sk c	i->2	
sk d	a->1	e->7	i->7	
sk e	k->1	n->1	r->1	
sk f	e->1	i->2	l->2	o->3	r->4	y->1	ö->6	
sk g	e->4	l->1	r->3	
sk h	a->5	j->2	ä->1	
sk i	 ->1	d->1	m->1	n->10	
sk j	o->1	u->2	ä->2	
sk k	a->9	l->1	o->23	u->3	v->1	
sk l	a->5	e->5	i->5	ä->1	ö->1	
sk m	a->6	e->3	i->3	o->1	y->2	
sk n	a->3	i->14	j->1	ä->1	
sk o	c->21	f->3	j->1	m->1	p->1	
sk p	a->2	e->2	l->2	o->16	r->5	u->1	
sk r	a->2	e->9	i->1	o->5	ä->1	å->1	ö->1	
sk s	i->5	k->1	m->1	o->5	t->12	y->6	
sk t	e->1	i->6	r->2	y->1	
sk u	n->7	p->3	r->1	t->12	
sk v	e->1	i->1	ä->2	
sk ä	n->1	
sk å	k->13	
sk ö	v->3	
sk, 	e->2	f->1	k->1	m->2	s->1	
sk-b	r->1	
sk-f	r->1	
sk-i	s->1	
sk-s	k->1	
sk. 	J->1	
sk.D	e->1	
sk.H	e->4	
sk.I	 ->2	n->1	
sk.J	a->1	
sk.M	e->1	
sk.O	m->1	
sk.V	i->1	
ska 	"->1	E->3	F->1	K->1	P->1	T->1	a->45	b->62	c->3	d->38	e->26	f->110	g->47	h->25	i->85	j->3	k->150	l->38	m->88	n->13	o->149	p->79	r->110	s->136	t->28	u->273	v->38	ä->2	å->18	ö->5	
ska,	 ->18	
ska.	D->1	E->3	F->1	H->1	J->2	P->1	V->3	
ska:	 ->2	
skab	e->1	
skad	 ->6	a->25	e->16	l->10	o->25	
skaf	f->26	
skak	a->2	
skal	:->1	a->3	d->1	i->3	l->670	v->1	
skam	 ->2	!->1	l->2	m->2	p->3	
skan	 ->16	,->1	.->1	a->3	d->31	s->2	
skap	 ->75	"->3	,->16	.->17	:->1	a->180	e->244	i->2	l->37	s->92	
skar	 ->31	,->2	.->3	a->1	e->6	n->2	p->2	r->1	t->1	
skas	 ->14	,->1	.->1	t->1	
skat	 ->8	,->1	.->2	s->3	t->66	
skbe	d->4	s->4	
ske 	-->1	I->1	a->2	b->3	d->4	e->3	f->4	g->3	h->2	i->13	k->7	l->5	m->3	n->3	o->8	p->8	r->2	s->4	t->3	u->6	v->5	ä->6	
ske!	Ä->1	
ske)	 ->2	
ske,	 ->6	
ske.	-->1	D->1	
sked	 ->3	.->1	a->4	e->7	
skek	v->1	
skel	n->3	
skem	å->3	ö->4	
sken	 ->17	,->1	
skeo	m->2	
skep	p->8	s->1	t->8	
sker	 ->41	,->1	.->6	a->18	e->1	i->5	n->6	ä->1	
skes	e->1	
sket	 ->3	,->1	r->3	s->1	t->15	
skev	a->2	
skfa	k->1	
skfr	i->1	
skfy	l->1	
skfö	r->1	
skha	n->6	
skhe	t->1	
skic	k->17	
skie	n->2	
skif	t->6	
skil	d->62	j->21	l->47	t->129	
skin	 ->3	e->3	g->3	l->1	
skip	a->3	n->9	
skis	k->4	s->4	
skju	t->31	
skka	p->1	
skko	m->2	
skla	n->22	r->1	u->2	
skli	g->43	m->2	
skni	n->77	v->1	
skoa	l->2	
skoe	f->1	
skof	ö->2	
skog	 ->3	a->10	e->5	r->1	s->19	
skoh	a->3	
skol	a->6	i->3	l->1	o->3	
skom	m->43	n->3	
skon	a->2	c->3	f->144	k->1	s->2	t->18	
skop	,->3	
skor	 ->40	,->3	.->1	n->24	s->14	t->2	
skos	l->1	t->10	
skot	t->166	
skou	r->1	
skov	 ->1	e->1	
skra	f->48	r->1	t->2	v->10	
skre	t->1	v->8	
skri	d->21	f->22	g->6	k->1	m->20	s->4	t->5	v->61	
skro	t->27	v->15	
skrä	c->9	d->1	m->5	n->11	p->1	
skt 	E->3	K->1	M->1	a->12	b->20	c->1	d->3	e->8	f->24	g->6	h->8	i->14	j->1	k->12	l->4	m->13	n->3	o->22	p->10	r->4	s->41	t->10	u->12	v->15	ä->5	å->1	ö->2	
skt!	N->1	
skt,	 ->7	
skt.	(->1	A->1	B->1	D->4	G->1	J->2	S->1	Å->1	
skta	l->1	
skug	g->3	
skul	d->3	l->496	t->9	
skun	n->1	
skup	p->1	
skur	 ->1	a->1	s->6	
skus	 ->1	s->61	
skut	a->6	e->78	
skva	,->1	l->7	
skvo	t->3	
skvä	r->13	
sky 	f->1	
skyd	d->108	
skyf	a->1	
skyh	ö->1	
skyl	d->29	l->5	
skym	t->1	
skyn	d->15	
skyv	ä->1	
skäl	 ->35	,->1	.->4	e->11	i->1	
skäm	d->1	m->2	t->1	
skän	k->2	n->1	s->2	
skär	 ->2	n->3	p->11	s->1	
skåd	a->3	l->6	n->1	
skål	e->1	
skår	,->1	
skön	h->1	
sköp	a->1	
skör	.->1	a->2	d->3	t->1	
sköt	 ->2	a->7	e->1	s->8	t->5	
sköv	l->1	
sla 	-->1	a->7	f->1	g->1	h->1	m->5	o->2	
sla"	.->1	
sla,	 ->2	
sla.	B->1	
slad	e->1	
slag	 ->331	,->33	.->39	;->1	?->3	a->1	e->138	i->16	n->33	r->1	s->27	
slak	t->1	
slam	 ->1	
slan	 ->4	d->17	
slap	p->3	
slar	 ->5	
slat	 ->1	
slav	a->1	i->1	
sled	a->39	
slen	,->1	.->1	
sler	 ->1	
sles	k->1	n->4	
slib	e->1	
slie	r->1	
slig	 ->29	a->84	h->13	t->32	
slin	g->2	j->2	s->1	
slip	p->2	
slir	a->1	
slis	t->48	
slit	a->1	
sliv	e->14	
slo 	o->1	
slo,	 ->2	
slob	b->1	
slog	 ->14	i->2	s->4	
slol	a->1	
slom	ä->1	
slop	p->2	
slor	 ->4	.->1	
slot	t->1	
slov	e->1	
sluk	a->3	
slum	p->4	r->1	
slun	t->1	
slus	s->2	
slut	 ->102	,->14	.->12	;->1	a->131	e->77	f->9	g->8	h->1	i->4	k->1	l->38	n->42	p->1	r->2	s->72	v->1	ä->5	
slyc	k->18	
släc	k->3	
släg	e->8	r->1	
släk	a->1	t->3	
släm	n->2	
slän	d->34	g->1	
släp	a->1	p->20	
slå 	E->1	a->6	e->4	f->6	i->1	k->4	m->2	n->1	p->1	r->1	s->2	v->4	
slåd	a->1	
slåe	n->1	
slån	g->1	
slår	 ->43	"->1	.->2	?->1	
slås	 ->25	.->1	s->1	
slöj	a->6	
slös	 ->2	a->9	e->3	h->39	n->2	t->3	
slöt	 ->3	
sm -	 ->1	
sm e	l->2	t->1	
sm f	ö->1	
sm h	ä->1	
sm i	n->1	
sm m	å->1	
sm o	c->12	m->6	
sm p	å->2	
sm s	a->1	o->5	
sm u	n->1	
sm ä	n->1	r->1	
sm ö	v->1	
sm, 	a->1	f->1	i->1	m->1	n->2	o->2	s->1	v->1	ä->1	
sm.D	e->6	ä->1	
sm.F	r->1	
sm.H	e->1	
sm.I	 ->2	
sm.J	a->1	
sm.M	e->1	
sm.N	ä->1	
sm.O	c->2	
sm.V	a->1	i->3	
sm?V	i->1	
smaj	o->1	
smak	t->4	ä->1	
sman	 ->1	.->1	n->14	
smar	k->15	
smas	k->2	
smat	t->1	
smed	b->9	d->2	e->95	i->3	l->5	v->2	
smek	a->2	
smen	 ->12	,->3	.->1	;->1	?->1	s->4	
smer	 ->4	.->2	n->3	
smet	o->6	
smid	i->3	
smil	j->5	
smin	i->16	
smis	k->2	
smit	a->1	n->1	t->1	
smod	e->2	
smol	n->1	
smom	e->5	
smon	o->1	
smot	o->1	
smug	g->1	
smul	a->1	
smus	s->1	
smut	s->3	
smyn	d->31	
smäd	e->1	
smäl	t->1	
smän	 ->16	g->2	n->15	
smär	k->1	r->1	t->2	
smäs	s->12	
små 	E->1	a->1	b->1	e->1	f->4	l->2	m->4	o->32	p->1	s->5	å->1	
små,	 ->2	
små.	D->1	
småf	ö->5	
småg	r->1	
smål	 ->7	.->2	e->2	s->1	
smån	i->4	
smås	k->1	
smöj	l->4	
smön	s->1	
smöt	e->2	
sna 	d->2	m->1	n->1	o->1	p->4	t->4	
sna,	 ->2	
snab	b->71	
snac	k->2	
snad	e->4	
snar	 ->5	.->2	a->36	k->1	l->1	t->27	
snat	 ->9	
sned	l->1	v->12	
snie	r->2	
snin	g->108	
snit	t->15	
sniv	å->33	
snor	m->7	
snyc	k->1	
snyh	e->1	
snäl	l->1	
snät	 ->1	e->2	
snäv	a->1	
snål	a->5	
snår	i->1	
snöj	d->2	e->1	
snöv	i->1	
so e	t->1	
so f	a->1	
so i	 ->1	
so o	c->1	
so ä	r->1	v->1	
so, 	d->1	
so- 	o->1	
soch	i->1	
soci	a->202	e->2	o->3	
sodl	i->1	
soef	f->1	
soff	e->2	
sofi	 ->2	,->1	n->1	s->1	
soft	 ->1	
sola	 ->1	
sold	a->2	
sole	r->7	
soli	d->33	
soll	m->1	
sols	k->1	
solu	t->140	
soly	c->1	
som 	"->4	-->3	1->1	2->1	3->1	4->2	A->5	B->10	C->3	D->5	E->41	F->6	G->3	H->3	I->2	J->3	L->4	M->2	N->1	O->1	P->4	R->3	S->3	T->4	W->2	a->131	b->154	c->5	d->254	e->158	f->280	g->126	h->289	i->216	j->115	k->183	l->97	m->184	n->94	o->67	p->66	r->103	s->268	t->99	u->88	v->317	y->1	Ö->1	ä->198	å->18	ö->14	
som,	 ->22	
somg	i->1	
soml	i->3	
somm	a->3	
somr	å->40	ö->1	
soms	p->1	
son 	a->1	f->1	h->3	i->3	k->1	o->1	s->2	v->1	
son,	 ->1	
son.	N->1	
sona	l->23	n->2	
sone	l->2	m->3	n->1	r->40	
song	s->1	
soni	 ->1	n->4	
sonl	i->34	
sons	 ->1	
sont	a->2	e->1	
sopa	 ->1	
sor 	M->2	T->3	e->1	m->1	o->1	
sor,	 ->4	
sor.	F->1	J->1	
sorb	e->1	
sord	f->21	n->15	
sore	l->1	
sorg	 ->9	a->11	l->3	s->1	
sori	e->1	s->3	
sorn	a->1	
sort	e->1	s->7	
sos 	o->2	
sos,	 ->1	
sosk	y->1	
sosä	k->2	
sot 	s->1	
sovj	e->1	
sovo	 ->25	,->11	.->12	?->2	N->1	k->2	s->7	
sovå	d->1	r->2	
sp",	 ->1	
sp. 	s->1	t->1	
spak	e->4	t->4	
span	e->1	j->1	s->10	
spar	a->7	i->3	k->5	l->1	s->1	t->4	
spat	i->2	
spec	i->85	
speg	l->12	
spek	t->148	u->4	
spel	 ->5	,->2	.->2	;->1	a->37	e->2	n->1	p->1	r->5	
spen	d->5	s->8	
sper	i->18	s->1	
spet	s->2	
spic	e->1	
spil	l->1	
spin	 ->1	
spir	e->3	
spis	k->1	
spla	c->3	n->31	t->9	
spli	k->7	t->4	
spo,	 ->1	
spol	i->128	
spon	d->1	s->2	t->4	
spor	t->110	
spos	 ->1	i->3	t->1	
spot	s->1	
spra	x->1	
spri	d->20	n->79	o->1	s->3	
spro	b->10	c->53	d->6	g->32	j->3	t->1	
spru	n->19	
språ	k->24	n->2	
spun	k->18	
spän	n->11	
spär	r->3	
spåf	ö->1	
spår	 ->4	,->2	a->4	e->1	n->2	
spök	e->3	s->1	
sque	,->1	
squi	n->1	
srad	 ->1	
srae	l->58	
sram	 ->1	,->1	a->4	e->2	
srap	p->6	
srea	k->1	
sred	a->2	
sref	o->2	
sreg	e->11	i->7	l->21	
srek	o->5	
srel	a->1	
srep	r->2	u->4	
sres	a->2	o->7	u->1	
srik	 ->5	,->1	a->5	t->6	
sril	a->1	
sris	k->3	
srol	l->1	
srub	r->1	
sruh	e->2	
srum	 ->1	
srun	d->2	
srut	i->1	
sryc	k->1	
srym	d->2	
sräd	s->1	
srät	t->61	
sråd	 ->2	,->1	.->2	e->4	g->14	
srör	e->2	
ss -	 ->1	
ss a	l->7	n->6	r->1	t->29	v->6	
ss b	a->1	e->6	i->1	r->2	u->1	
ss d	a->2	e->11	o->3	ä->6	å->2	
ss e	g->3	k->1	l->2	m->2	n->10	t->4	u->1	x->1	
ss f	l->1	o->5	r->5	u->3	å->1	ö->19	
ss g	e->5	j->1	r->2	ä->1	
ss h	a->4	e->1	i->1	o->1	u->1	ä->1	
ss i	 ->25	d->1	n->16	
ss k	a->1	l->1	o->7	v->1	
ss l	a->1	e->1	i->2	u->1	å->1	
ss m	a->2	e->14	i->1	o->3	y->3	ä->1	å->6	
ss n	a->2	e->2	y->2	ä->4	å->1	
ss o	a->1	c->14	d->1	e->1	f->1	m->19	r->7	s->1	
ss p	a->1	e->1	o->2	r->2	å->16	
ss r	a->1	e->5	y->1	ä->3	ö->1	
ss s	a->6	e->1	i->2	j->10	k->3	l->3	o->20	t->4	v->1	y->1	ä->1	å->3	
ss t	a->1	i->17	j->1	o->1	r->2	v->1	y->2	
ss u	n->4	p->1	t->8	
ss v	a->7	e->3	i->5	ä->3	å->1	
ss y	t->1	
ss ä	n->3	r->10	
ss å	s->2	t->14	
ss ö	d->1	m->1	r->1	v->3	
ss".	D->1	
ss) 	o->1	
ss, 	T->1	a->2	d->1	e->1	f->2	g->1	h->1	i->2	m->3	o->3	s->3	v->2	ä->1	å->1	
ss.A	l->1	
ss.D	e->6	i->1	ä->1	
ss.E	n->2	u->1	
ss.F	r->2	
ss.H	e->2	
ss.J	a->4	
ss.M	a->1	å->1	
ss.N	ä->1	å->1	
ss.S	l->1	
ss.V	a->1	i->5	å->1	
ss.Ä	v->2	
ss: 	k->1	
ss?.	 ->1	
ss?J	o->1	
ss?V	i->1	
ssa 	-->1	1->1	2->3	3->1	P->1	a->44	b->26	c->1	d->10	e->4	f->61	g->12	h->15	i->19	k->27	l->18	m->35	n->4	o->24	p->42	r->32	s->46	t->20	u->12	v->14	ä->32	å->9	ö->2	
ssa!	L->1	
ssa,	 ->4	
ssa.	B->1	D->2	I->1	J->1	M->3	
ssab	o->8	
ssad	 ->5	,->1	e->2	ö->1	
ssag	 ->1	e->1	
ssak	r->1	
ssal	a->1	
ssam	a->3	h->5	m->1	t->5	
ssan	d->3	k->1	t->21	
ssar	 ->4	,->1	b->3	n->1	
ssas	 ->7	
ssat	 ->1	
ssav	g->1	
ssbe	l->5	
ssbr	u->10	
ssch	e->1	
sse 	(->1	a->6	d->3	f->5	l->1	o->1	p->1	s->2	t->1	
sse,	 ->5	
sse-	N->1	
sse.	F->1	M->2	
sse?	E->1	
ssed	 ->1	
ssek	r->1	t->18	
ssel	 ->11	!->1	,->5	-->3	.->2	b->1	f->1	o->1	s->103	
ssen	 ->57	,->21	.->32	?->1	N->1	a->5	s->7	t->1	
sser	 ->5	,->2	a->19	i->1	l->13	n->8	v->1	
sset	 ->4	,->1	ê->2	
ssfa	l->1	
ssfo	r->1	s->1	
ssfö	r->4	
ssgy	n->7	
sshe	t->4	
sshu	s->1	
sshä	n->1	
ssid	a->1	
ssif	f->3	i->9	
ssig	 ->3	a->15	t->14	
ssil	 ->1	a->2	
ssim	i->2	
ssin	 ->1	
ssio	n->1223	
ssis	k->5	t->2	
ssit	u->4	
ssiv	 ->3	.->1	a->4	t->4	
ssjö	f->1	
sska	d->3	n->1	p->1	t->1	
sske	d->3	
sski	c->1	f->2	l->5	p->3	
ssko	n->2	
sskr	i->1	o->7	
ssky	d->3	l->2	
sskä	l->3	
sskö	t->6	
ssla	 ->1	d->1	n->6	r->5	t->1	
ssly	c->18	
sslö	s->2	
ssme	d->4	
ssna	 ->9	,->1	d->4	r->5	t->9	
ssni	n->7	
ssnö	j->3	
sso 	e->1	i->1	o->1	ä->2	
sso,	 ->1	
ssoc	i->1	
sson	i->1	
ssor	 ->7	,->2	
sspe	l->1	
sspr	i->1	å->1	
ssre	g->1	s->2	
ssrä	t->2	
sst 	b->1	d->1	f->1	j->1	k->2	m->1	n->1	
ssta	 ->1	d->3	g->8	n->7	r->3	t->293	v->1	
sste	 ->4	x->1	
ssti	l->1	
ssto	l->1	
sstr	a->11	o->3	u->5	ä->2	ö->4	
ssty	r->7	
sstä	l->24	m->21	n->4	
sstå	l->1	
sstê	t->1	
sstö	d->30	r->1	
ssue	l->1	
ssup	p->2	
ssus	e->1	
ssut	o->61	
ssvä	r->4	
ssvå	r->1	
ssyn	e->1	p->1	
ssys	 ->1	s->1	t->55	
ssäk	e->65	r->1	
ssäl	l->7	
ssän	k->1	
ssät	t->10	
st -	 ->3	
st 1	 ->1	0->1	2->1	
st 2	5->1	
st 3	 ->2	
st 4	0->1	
st 5	,->1	
st 7	0->1	
st 9	 ->1	
st D	a->1	
st E	u->3	
st I	n->1	
st M	i->1	
st P	e->1	
st a	c->2	k->1	l->4	n->9	r->3	t->12	v->16	
st b	e->11	i->1	l->1	
st c	a->1	
st d	a->1	e->25	r->4	y->1	ä->6	å->3	
st e	f->5	n->8	r->1	t->8	x->1	
st f	a->4	l->1	o->1	r->9	u->1	å->2	ö->28	
st g	e->6	j->3	l->2	r->1	ä->1	å->1	ö->2	
st h	a->20	ä->3	ö->1	
st i	 ->26	l->1	n->16	
st j	u->2	
st k	a->7	o->10	r->4	u->4	
st l	a->2	e->1	i->1	o->3	ä->3	å->2	ö->2	
st m	e->11	i->6	o->5	å->9	ö->3	
st n	e->1	i->1	o->2	u->10	y->1	ä->10	å->2	ö->1	
st o	b->1	c->34	f->1	l->1	m->11	p->1	r->1	v->1	
st p	e->5	l->1	o->3	r->6	å->30	
st r	a->1	e->5	i->2	u->1	ä->2	ö->3	
st s	a->7	e->4	i->1	k->15	l->1	o->7	t->7	v->3	y->2	ä->3	å->2	
st t	a->6	i->16	r->4	v->4	ä->1	
st u	n->1	p->3	t->13	
st v	a->7	e->1	i->37	ä->3	
st ä	r->11	
st å	r->1	t->4	
st ö	n->1	v->3	
st!D	ä->1	
st!T	v->1	
st, 	P->1	a->1	d->5	e->4	f->1	h->2	i->2	k->1	m->3	o->2	p->1	s->2	v->1	
st- 	o->1	
st-b	e->5	
st. 	A->1	
st.A	c->1	
st.D	e->3	
st.E	f->1	
st.F	ö->2	
st.G	i->1	
st.J	a->3	
st.K	o->1	ä->1	
st.M	e->1	i->1	
st.N	u->1	ä->1	
st.V	a->1	i->3	
st.Ä	r->1	
st: 	m->1	
st?N	e->1	
st?V	i->1	
sta 	a->17	b->23	c->1	d->29	e->12	f->52	g->40	h->33	i->15	k->15	l->4	m->39	n->7	o->17	p->52	r->34	s->51	t->20	u->8	v->18	ä->20	å->2	ö->4	
sta,	 ->16	
sta.	)->1	-->1	.->1	D->3	E->1	H->1	S->1	V->5	
sta:	 ->5	
sta;	 ->2	
sta?	N->1	
staN	ä->1	
staa	f->1	
stab	 ->1	e->1	i->22	u->1	
stac	k->1	
stad	 ->7	,->1	.->3	e->20	g->28	i->8	k->24	s->4	t->1	
stag	 ->2	,->1	.->3	a->52	e->2	n->2	
stai	n->22	
stak	,->1	a->5	l->1	
stal	i->2	l->3	t->1	
stam	p->1	
stan	 ->64	,->5	.->14	b->1	d->41	k->5	n->7	s->42	t->4	
star	 ->25	e->2	i->1	k->61	t->16	
stas	 ->5	,->1	i->1	t->1	
stat	 ->59	,->7	.->13	e->363	i->23	l->98	s->50	t->1	u->10	
stau	r->1	
stav	 ->1	l->1	
stba	n->4	
stbe	s->1	v->1	
stbi	l->1	
stbl	o->1	
stbr	i->1	
stde	m->11	
ste 	-->3	E->8	F->1	I->1	a->40	b->49	c->2	d->62	e->18	f->58	g->41	h->16	i->35	j->11	k->33	l->10	m->46	n->17	o->32	p->14	r->27	s->82	t->51	u->36	v->114	ä->13	å->22	ö->8	
ste,	 ->4	
ste.	D->1	F->1	V->1	
ste:	 ->1	
sted	t->4	
stee	n->5	r->1	
stef	e->1	r->1	ö->5	
steg	 ->55	,->3	.->2	e->7	
stei	n->1	
stek	n->2	
stel	a->2	e->1	s->5	t->1	
stem	 ->75	,->9	.->11	:->1	a->15	e->81	ä->37	
sten	 ->33	"->1	,->12	.->9	N->1	a->3	d->2	e->1	k->1	s->8	t->1	
step	r->1	
ster	 ->119	!->1	"->2	,->19	.->32	a->33	d->39	f->3	i->17	m->2	n->87	p->3	r->147	s->1	
stes	 ->2	e->2	t->1	
stet	 ->1	.->3	
steu	r->9	
stex	t->3	
stfl	i->1	
stfu	l->1	
stfä	l->8	
stfö	r->8	
stgr	u->3	
stgö	r->3	
stha	n->1	
stho	m->3	
sthä	l->1	
sthå	l->1	
stia	n->1	
stic	e->4	k->5	
stid	 ->2	,->1	e->6	n->2	s->3	
stie	r->1	
stif	t->128	
stig	 ->1	a->4	e->2	h->1	i->2	l->4	m->1	t->4	
stik	 ->3	e->3	
stil	 ->2	l->59	
stim	u->11	
stin	a->10	d->2	i->4	k->3	r->1	s->8	
stio	n->1	
stip	e->1	
stis	k->93	
stit	i->6	u->159	
stjä	n->7	r->2	
stkl	a->1	
stko	m->1	
stku	b->1	s->1	
stkä	l->1	
stla	g->1	n->2	
stli	g->1	n->2	
stlä	g->2	n->1	
stma	k->1	r->1	
stmy	n->3	
stmä	n->2	
stna	d->108	r->1	
stni	n->72	
stnä	m->2	
sto 	h->1	v->1	
stod	 ->15	o->1	
stol	 ->7	.->2	a->25	e->46	k->1	p->1	s->10	t->11	
stom	r->2	
ston	e->27	
stop	-->1	p->19	
stor	 ->103	,->1	.->1	a->157	d->2	e->4	f->2	h->1	i->36	k->1	m->27	s->4	t->41	
stow	n->3	
stpa	r->5	
stra	 ->8	d->1	f->40	k->1	m->3	n->1	r->17	t->91	x->2	
stre	a->8	c->1	g->1	r->15	s->2	t->1	
stri	 ->11	,->3	-->1	b->1	c->6	d->23	e->8	f->4	k->25	l->2	n->83	p->2	s->3	
stro	e->2	f->90	n->4	t->1	
stru	e->5	k->186	m->52	n->4	
stry	k->34	p->1	
strä	c->32	n->65	t->3	v->31	
strå	e->1	l->5	
strö	j->1	k->3	m->19	
sts 	p->1	v->1	
sts.	D->1	S->1	
stsa	m->2	
stse	k->2	
stsl	a->2	o->2	å->17	
stst	ä->51	
stsv	a->1	
stto	n->1	
stty	s->2	
stu 	m->1	
stud	e->5	i->9	
stug	o->1	
stul	l->1	
stum	 ->1	
stun	d->17	
stur	i->2	
stut	v->2	
stva	k->1	
stve	r->1	
stvi	k->3	s->1	
stvä	r->1	
styc	k->5	
stym	p->3	
styr	 ->1	a->11	e->15	k->17	n->7	s->2	
städ	a->2	e->19	
stäl	l->426	
stäm	d->19	m->186	n->2	p->2	s->1	t->16	
stän	 ->1	d->108	g->11	k->6	
stär	k->51	
stät	h->1	
stäv	 ->1	j->1	
stå 	a->16	d->3	e->1	f->21	h->2	i->5	k->4	n->2	o->3	s->1	t->1	u->2	v->4	
stå,	 ->3	
stå.	F->1	J->1	
stå:	 ->1	
ståd	d->2	
ståe	l->14	n->32	
stål	f->5	g->1	i->25	s->5	v->5	
stån	d->226	
står	 ->177	,->3	.->3	
stås	 ->6	
ståt	t->30	
stêt	e->1	
stöd	 ->157	,->14	.->38	;->1	?->1	d->2	e->119	j->72	m->2	n->1	p->1	r->2	s->12	å->5	
stöl	d->1	
stör	 ->4	a->5	d->3	e->5	i->2	n->5	r->73	s->37	t->3	
stöt	a->3	e->2	f->1	t->13	
sual	i->1	
subj	e->1	
subs	i->23	t->4	
subv	e->10	
succ	e->5	
sudd	a->1	
suel	l->2	
suga	r->1	
sul 	o->1	s->1	
sul.	V->1	
sule	r->3	
sult	a->111	b->1	e->9	
sum 	o->1	
sumb	a->1	
sume	n->61	
summ	a->6	e->6	o->8	
sumt	i->2	
sund	 ->1	a->4	e->3	i->3	
sune	r->1	
supp	e->1	f->3	g->1	s->1	
supr	a->1	
surd	 ->1	
surs	b->1	e->46	f->1	s->1	t->1	
surt	 ->2	
sus 	k->2	o->1	
suse	n->1	
susp	e->1	
suta	n->3	
sutb	i->9	y->6	
suto	m->61	
sutr	u->1	y->4	
suts	a->1	k->2	l->1	ä->2	
sutt	i->1	r->1	
sutv	e->2	ä->1	
sutö	v->1	
suve	r->17	
sv. 	M->1	V->1	m->1	
sv.,	 ->1	
sv.?	A->1	
sv.S	v->1	
svag	 ->3	a->28	h->12	n->1	
sval	,->1	
svan	s->2	
svar	 ->96	,->26	.->35	?->1	a->94	e->73	i->56	s->81	t->2	v->2	
svat	t->2	
svek	 ->2	
sven	s->2	t->1	
svep	 ->1	s->1	t->1	
sver	k->7	
svik	e->7	n->1	
svil	j->2	l->20	
svin	n->15	s->1	
svis	 ->25	,->6	.->1	
svun	n->4	
sväg	,->1	
sväl	t->2	
sväm	m->3	n->4	
svän	l->2	
svär	d->14	e->1	l->6	r->4	t->4	
sväs	e->6	
svät	s->1	
sväv	n->1	
svåg	 ->1	e->1	
svån	g->1	
svår	 ->5	a->25	b->2	d->1	i->31	l->2	t->28	ö->1	
swag	e->1	
sydd	a->1	
syde	u->1	
sydk	u->1	
sydv	ä->1	
sydö	s->1	
syft	a->36	e->38	
syko	l->1	
syl 	g->1	o->3	
syl,	 ->2	
syl-	 ->1	
syl.	D->1	J->1	V->1	
sylb	e->1	
sylf	ö->2	
sylr	ä->2	
syls	ö->6	
symb	o->9	
symp	a->8	t->1	
syn 	-->1	a->2	g->1	i->2	o->5	p->4	t->65	v->1	ä->2	
syn,	 ->2	
syn.	A->1	E->1	S->2	
syn;	 ->1	
syna	 ->1	s->3	
synd	 ->4	a->2	e->1	r->1	
syne	n->6	r->2	s->1	
synl	i->8	
synn	e->52	
syno	n->1	
synp	u->29	
syns	 ->1	t->2	ä->4	
synt	 ->2	,->1	e->1	
synv	i->12	
syra	 ->3	
syri	e->4	s->4	
sys 	f->1	
syss	e->103	l->6	
syst	e->191	
säg:	 ->1	
säga	 ->148	,->15	.->2	:->4	n->2	r->4	s->5	
säge	l->8	r->73	
sägn	e->1	i->1	
sägs	 ->5	
säke	r->321	
säkr	a->40	i->24	
säkt	 ->7	.->1	a->4	e->3	
sälj	a->5	n->3	
säll	a->2	s->10	
sämn	e->2	
sämr	a->10	e->5	
säms	t->5	
sänd	a->6	e->11	n->1	r->4	
sänk	a->5	n->2	t->1	
sär 	d->2	s->1	
sära	r->1	
särb	e->1	
säre	n->4	
särk	i->1	
särs	k->156	
säso	n->1	
säte	.->1	
sätt	 ->181	,->25	.->47	:->2	?->2	a->111	e->88	l->1	n->211	s->14	
så "	m->1	
så -	 ->2	
så 1	9->1	
så E	u->4	
så F	l->1	
så M	o->1	
så a	b->1	k->1	l->7	m->1	n->11	r->1	t->179	v->10	
så b	a->4	e->16	i->2	l->5	o->3	r->5	y->2	ä->2	ö->4	
så d	e->29	i->1	o->1	r->2	ä->2	
så e	f->3	k->1	n->26	r->1	t->10	
så f	a->5	i->7	o->4	r->10	u->2	å->9	ö->29	
så g	a->1	e->5	l->1	o->2	r->3	ä->3	å->3	ö->5	
så h	a->13	e->9	j->4	o->4	u->3	ä->6	å->1	ö->1	
så i	 ->23	a->1	l->1	m->1	n->29	
så j	a->2	
så k	a->23	l->3	o->26	r->5	u->2	ä->1	ö->1	
så l	i->5	y->1	ä->16	å->12	
så m	a->1	e->17	i->3	o->1	y->38	å->30	ö->2	
så n	o->3	y->1	ä->5	å->5	ö->4	
så o	a->2	c->1	f->4	g->1	m->8	r->1	
så p	a->4	e->1	l->1	o->1	å->16	
så r	a->1	e->4	i->2	ä->2	å->1	ö->2	
så s	a->7	e->8	i->1	j->1	k->21	l->1	m->6	n->28	o->22	p->1	t->20	v->4	ä->30	å->3	
så t	a->18	i->17	o->1	r->4	y->1	ä->1	
så u	n->4	p->12	t->7	
så v	a->16	e->4	i->42	ä->4	å->3	
så z	i->1	
så ä	g->1	n->2	r->33	
så å	t->3	
så ö	p->1	v->3	
så, 	a->2	e->1	f->2	h->2	i->2	m->1	n->1	o->4	s->2	t->1	
så. 	D->1	
så.D	e->2	
så.I	 ->1	n->1	
så.J	a->1	
så.N	i->1	
så.O	c->1	
så.P	å->1	
så: 	a->1	
såda	n->163	
såg 	a->7	d->2	e->1	i->1	n->1	o->1	s->2	u->2	Ö->1	
sågs	 ->2	.->2	
sågv	e->1	
såhä	r->1	
såld	e->2	
såle	d->40	
sålu	n->4	
sång	 ->1	e->2	
sårb	a->3	
såre	t->1	
såso	m->32	
såte	 ->1	r->1	
såtg	ä->11	å->1	
såti	l->1	
såvi	d->3	
såvä	l->40	
sí ä	r->1	
söda	n->1	
söde	 ->1	
södr	a->6	
sök 	a->4	i->5	o->1	s->1	
sök,	 ->2	
söka	 ->41	,->1	n->7	r->6	s->5	
söke	n->1	r->21	t->4	
sökn	i->24	
sökt	 ->14	e->6	
sönd	e->7	
söne	r->1	
sörj	a->9	d->1	e->2	n->4	
söve	r->15	
sövn	i->1	
t "E	U->1	
t "K	u->2	v->2	
t "O	l->1	
t "P	o->1	
t "e	g->1	k->1	n->1	u->1	
t "k	u->1	
t "o	b->1	
t "r	e->2	
t (5	7->1	
t (8	0->2	
t (9	6->1	
t (B	5->2	
t (C	E->1	
t (E	U->2	
t (F	P->1	
t (I	C->1	F->1	
t (S	P->1	
t (a	r->1	
t (d	e->1	
t (f	i->2	
t (h	ä->1	
t (i	 ->1	n->1	
t (k	o->1	
t (t	.->1	y->1	
t (Ö	V->1	
t , 	d->1	
t - 	a->7	d->7	e->5	f->6	g->2	h->2	i->5	j->4	k->4	m->3	n->3	o->12	p->1	s->11	t->1	u->1	v->9	ä->2	å->2	ö->2	
t -,	 ->2	
t -e	r->1	
t 1 	0->1	u->1	
t 1,	 ->1	
t 10	 ->2	
t 11	 ->1	
t 12	 ->1	
t 13	 ->1	
t 18	0->1	
t 19	4->1	9->18	
t 2 	i->2	
t 20	0->1	
t 21	:->1	
t 22	 ->1	
t 23	,->1	
t 25	 ->2	
t 26	 ->1	
t 27	 ->1	
t 3 	p->2	
t 39	 ->1	
t 4 	i->1	l->1	
t 40	 ->1	0->2	
t 48	 ->1	
t 5 	0->1	
t 5,	 ->1	5->1	
t 50	-->1	
t 6 	o->1	
t 7 	i->1	
t 70	 ->1	0->2	
t 8 	r->1	
t 80	 ->1	
t 88	/->2	
t 9 	f->1	
t 90	 ->1	
t 93	 ->1	
t 94	/->1	
t 95	 ->1	
t 98	 ->1	
t : 	P->1	
t AB	B->1	
t Ad	o->1	
t Ai	d->1	
t Ak	k->1	
t Al	e->1	t->3	
t Am	s->3	
t As	s->1	
t Au	s->1	
t BN	P->1	
t Ba	r->3	
t Be	r->2	
t Bo	u->1	
t Br	e->1	o->1	y->1	
t CE	N->1	
t Ca	m->1	s->1	
t Cl	i->1	
t D 	k->1	
t Da	l->2	n->4	
t De	 ->1	
t Du	b->1	i->1	
t EG	-->10	:->2	
t EI	F->1	
t EK	S->1	
t EL	D->1	
t EU	 ->8	-->4	.->3	:->7	
t El	l->1	
t Eq	u->8	
t Er	i->3	
t Eu	r->111	
t Ev	a->1	
t FE	O->1	
t FN	-->1	:->1	
t FP	Ö->3	
t Fl	o->4	
t Fr	a->3	
t Fö	r->5	
t Ga	r->1	
t Go	e->1	
t Gr	e->3	u->1	ö->1	
t Ha	d->1	i->3	
t He	b->1	
t I 	T->1	
t IC	E->1	
t IN	T->1	
t In	t->2	
t Ir	l->1	
t Is	r->4	
t It	a->3	
t Jo	n->3	
t Jö	r->3	
t Ka	r->1	
t Ki	r->1	
t Ko	s->2	u->2	
t Ku	l->3	
t Ky	o->2	
t La	n->1	
t Le	a->2	
t Ma	l->1	r->1	
t Mi	d->1	n->1	
t Mo	n->1	r->3	
t Mü	n->1	
t Na	t->1	
t OL	A->3	
t Pa	t->1	
t Pe	t->1	
t Po	r->6	
t RI	N->2	
t Ra	n->2	p->3	
t Ro	t->1	
t SE	M->1	
t Sa	n->1	v->1	
t Sc	h->1	
t Sj	u->1	ö->1	
t So	k->1	u->1	
t St	o->3	
t Su	d->1	
t Sv	e->1	
t TV	-->1	
t Th	e->3	
t Ti	b->1	
t To	d->1	t->2	
t Tu	r->14	
t UN	M->1	
t Va	t->1	
t Ve	r->1	
t Vo	d->1	
t Vä	r->1	
t Wa	f->1	l->1	
t Wu	l->1	
t ab	s->8	
t ac	c->12	
t ad	 ->1	d->1	e->3	m->2	
t ag	e->16	
t ai	d->1	
t ak	t->17	u->1	
t al	b->1	d->3	i->1	l->112	t->2	
t am	b->3	e->3	
t an	a->10	d->63	f->5	g->16	l->3	m->2	n->32	o->2	p->2	s->95	t->70	v->31	
t ar	a->1	b->102	g->1	r->3	t->15	v->1	
t as	y->3	
t at	t->816	
t av	 ->485	a->1	b->2	d->1	f->4	g->15	h->3	l->4	s->60	t->18	v->6	
t ba	d->1	k->23	l->1	n->2	r->20	s->1	x->1	
t be	 ->3	a->10	d->11	f->15	g->29	h->47	k->44	l->7	m->4	n->1	r->36	s->83	t->114	v->35	
t bi	b->3	d->24	f->1	g->1	l->22	n->7	o->1	s->9	t->1	
t bl	.->2	a->6	e->1	i->73	u->1	y->3	
t bo	 ->1	g->1	m->1	r->17	s->2	t->1	
t br	a->32	e->10	i->11	o->9	y->8	ä->2	å->4	
t bu	d->11	
t by	g->18	r->3	
t bä	r->1	s->7	t->22	
t bå	d->7	t->1	
t bö	r->60	
t ca	s->1	
t ce	m->2	n->5	
t ch	a->2	
t ci	r->1	t->1	v->6	
t d)	 ->1	
t da	g->10	n->8	t->9	
t de	 ->236	,->1	b->11	c->2	f->7	l->25	m->27	n->292	p->1	r->5	s->50	t->684	
t di	a->1	l->2	p->1	r->40	s->38	v->1	
t dj	u->3	ä->4	
t do	c->4	k->11	l->2	m->10	
t dr	a->30	i->9	å->1	ö->3	
t du	b->2	
t dy	k->1	n->2	r->3	
t dä	m->2	r->42	
t då	 ->13	l->5	
t dö	 ->1	d->2	l->3	m->6	r->1	
t e)	 ->1	
t e-	m->1	
t ed	e->1	
t ef	f->20	t->42	
t eg	e->31	n->4	
t ek	o->24	
t el	-->1	e->3	i->1	l->38	
t em	b->1	e->3	o->5	
t en	 ->215	a->13	b->5	d->28	e->3	g->8	h->16	i->2	k->30	l->8	o->6	s->4	t->2	v->1	
t ep	o->1	
t er	 ->9	,->1	a->4	b->4	f->4	h->2	i->3	k->13	s->6	t->7	
t et	a->5	t->118	
t eu	r->48	
t ev	e->5	
t ex	 ->2	a->7	c->2	e->30	i->1	p->9	t->7	
t f.	d->1	
t fa	i->1	k->65	l->34	n->12	r->11	s->28	t->13	
t fe	d->1	l->11	m->14	n->1	
t fi	c->4	n->221	s->4	
t fj	ä->4	
t fl	e->27	y->7	
t fo	d->1	g->1	k->2	l->7	n->1	r->56	t->1	
t fr	a->104	e->11	i->15	u->4	y->1	ä->42	å->121	
t fu	l->20	n->17	
t fy	l->1	r->2	s->1	
t fä	n->1	s->2	
t få	 ->100	.->2	g->3	r->26	t->3	
t fö	d->1	l->14	r->1226	
t ga	m->4	n->4	r->21	v->3	
t ge	 ->55	.->1	m->43	n->95	o->2	r->12	s->1	t->2	
t gi	c->2	l->1	v->5	
t gj	o->7	
t gl	a->6	o->3	ä->11	
t go	d->82	t->13	
t gr	a->24	e->2	i->4	u->15	ä->2	ö->2	
t gy	n->6	
t gä	l->223	r->1	
t gå	 ->30	.->1	r->14	t->3	
t gö	r->141	
t ha	 ->55	,->1	d->9	f->4	l->4	m->3	n->130	r->208	
t he	d->1	l->27	m->8	n->1	r->1	s->1	
t hi	n->11	s->4	t->10	
t hj	ä->20	
t ho	n->8	p->7	r->2	s->12	t->9	
t hu	g->3	m->2	n->2	r->18	s->3	v->3	
t hy	c->2	s->1	
t hä	l->1	n->32	r->68	v->2	
t hå	l->33	n->1	r->7	
t hö	g->23	j->3	l->2	r->24	
t i 	2->1	A->3	B->6	C->1	D->2	E->13	F->8	G->1	H->9	I->5	K->5	L->1	M->4	N->2	P->4	S->2	T->8	a->23	b->10	d->91	e->25	f->51	g->11	h->15	j->3	k->15	l->6	m->18	n->5	o->10	p->11	r->13	s->65	t->9	u->7	v->26	Ö->4	ä->2	å->3	ö->2	
t i.	D->1	
t ia	k->1	
t ib	l->6	
t ic	k->4	
t id	e->6	é->3	
t if	r->15	
t ig	e->9	å->1	
t il	l->2	s->2	
t im	m->3	p->3	
t in	 ->9	b->7	c->2	d->1	f->59	g->31	h->1	i->21	k->1	l->17	n->59	o->46	r->28	s->49	t->290	v->9	
t ir	l->3	o->1	r->4	
t is	o->4	
t it	a->4	
t ja	 ->3	g->105	p->1	
t jo	b->1	r->5	
t ju	 ->7	n->1	r->7	s->13	
t jä	m->8	r->1	
t ka	l->2	m->6	n->108	o->1	p->6	s->1	t->1	
t ke	m->1	
t kl	a->53	o->2	y->1	
t kn	a->1	u->1	y->4	ä->1	
t ko	a->2	l->9	m->337	n->92	p->1	r->37	s->14	
t kr	a->19	i->21	o->1	ä->52	
t ku	l->18	n->68	s->1	
t kv	a->15	i->4	ä->2	
t ky	l->1	
t kä	m->1	n->18	r->7	
t kö	l->3	n->1	p->1	t->2	
t la	b->1	d->2	g->17	n->55	p->3	s->1	w->1	
t le	d->27	g->3	k->1	v->9	
t li	b->1	d->2	g->15	k->11	l->4	n->3	s->1	t->17	v->11	
t lj	u->2	
t lo	b->1	c->1	g->4	j->2	k->1	t->3	v->1	
t lu	d->2	f->1	g->2	t->2	
t ly	c->12	d->1	f->2	s->8	
t lä	g->68	m->21	n->18	r->5	s->1	t->8	x->1	
t lå	g->3	n->13	t->13	
t lö	f->2	n->1	p->8	s->21	
t ma	j->4	k->2	n->218	r->23	s->2	t->8	x->2	
t me	d->350	k->1	l->39	n->16	r->36	s->7	t->1	
t mi	g->72	l->14	n->88	r->1	s->16	t->5	x->1	
t mo	b->2	d->12	g->1	n->3	r->1	t->71	
t mu	l->3	n->2	s->1	
t my	c->89	n->12	t->1	
t mä	n->11	r->6	t->1	
t må	h->1	l->27	n->20	s->106	t->1	
t mö	d->1	j->47	r->1	t->8	
t na	m->2	r->2	t->16	z->2	
t ne	d->10	g->5	k->1	r->3	
t ni	 ->51	,->2	o->2	v->3	
t no	g->20	m->1	r->6	t->3	
t nr	 ->1	
t nu	 ->36	,->3	.->2	m->1	v->10	
t ny	 ->1	a->23	b->1	d->1	k->2	l->5	n->1	s->1	t->27	v->1	
t nä	m->6	r->72	s->8	t->2	
t nå	 ->10	d->1	g->58	r->1	
t nö	d->29	j->4	t->2	
t oa	c->12	v->1	
t ob	e->8	s->1	
t oc	h->666	k->58	
t od	j->1	
t oe	f->1	g->1	n->1	r->2	
t of	f->16	t->7	ö->4	
t og	r->2	
t ok	l->2	r->1	u->1	
t ol	a->1	i->2	j->7	y->6	ä->1	
t om	 ->225	,->1	.->5	b->2	d->2	e->5	f->17	h->1	k->3	o->2	p->1	r->44	s->6	v->3	ö->5	
t on	d->2	t->1	ö->3	
t op	a->1	e->2	p->1	r->2	t->2	
t or	d->25	e->2	g->10	i->3	o->15	s->2	w->1	ä->2	
t os	a->1	s->50	v->2	y->1	ä->1	
t ot	i->5	y->2	ä->1	
t ov	ä->2	
t oä	n->1	
t oö	v->2	
t pa	k->1	l->1	p->1	r->99	s->5	t->1	
t pe	a->1	k->3	n->10	r->27	s->2	
t pi	l->1	
t pl	a->23	ö->1	
t po	l->39	p->2	r->61	s->29	t->1	ä->3	
t pr	a->11	e->14	i->26	o->89	ä->1	ö->2	
t pu	n->5	
t på	 ->276	,->3	.->2	:->1	?->1	b->3	d->1	g->5	m->5	p->8	s->8	t->3	v->10	
t ra	d->3	k->4	m->2	n->1	p->2	s->2	t->4	
t re	a->4	d->18	e->1	f->19	g->48	k->5	l->3	n->7	p->8	s->49	t->6	v->4	
t ri	d->1	k->33	m->7	n->3	s->6	
t ro	 ->1	p->1	
t ru	b->1	l->1	m->10	t->1	
t ry	k->4	
t rä	c->14	d->5	k->1	t->47	
t rå	d->52	k->1	
t rö	r->19	s->38	t->1	
t s.	k->1	
t sa	d->7	g->9	k->18	l->1	m->107	n->7	t->5	
t se	 ->58	d->11	g->7	k->3	m->2	n->18	r->16	s->1	t->27	x->5	
t si	d->2	f->1	g->66	k->5	n->22	s->7	t->15	
t sj	u->8	ä->21	ö->1	
t sk	a->181	e->25	i->12	j->6	o->2	r->12	u->97	y->39	ä->15	ö->3	
t sl	a->9	i->1	u->22	ä->5	å->7	ö->2	
t sm	i->1	ä->1	å->2	
t sn	a->20	ö->1	
t so	c->20	l->4	m->517	r->2	
t sp	a->8	e->28	o->2	r->4	å->2	ö->1	
t st	a->57	e->19	i->5	o->68	r->31	u->1	y->9	ä->47	å->36	ö->163	
t su	b->4	c->1	d->1	n->1	v->2	
t sv	a->35	e->2	å->19	
t sy	f->15	m->3	n->7	r->1	s->46	
t sä	g->43	k->40	l->1	m->2	n->7	r->14	t->176	
t så	 ->66	,->1	.->2	d->49	g->1	l->3	s->2	v->6	
t sö	d->1	k->4	r->2	
t t.	o->1	
t ta	 ->95	.->1	?->1	b->1	c->38	g->10	k->1	l->24	n->5	p->1	r->10	s->5	
t te	c->5	k->2	m->1	o->1	r->3	x->2	
t th	e->1	
t ti	b->1	d->32	l->368	o->1	t->5	
t tj	u->1	ä->4	
t to	g->1	l->6	m->2	n->1	p->1	r->1	t->5	
t tr	a->13	e->27	o->7	u->2	y->2	ä->11	
t tu	f->1	n->3	r->1	s->1	
t tv	e->5	i->11	å->11	
t ty	c->7	d->30	s->5	v->2	
t tä	c->1	m->2	n->18	p->2	
t tå	g->2	l->1	
t ul	t->1	
t un	d->128	i->12	
t up	p->181	
t ur	 ->8	a->6	h->1	s->7	v->4	
t ut	 ->11	,->9	.->7	a->37	b->7	e->8	f->18	g->15	h->1	i->3	j->3	k->2	l->3	m->17	n->17	o->3	p->3	r->4	s->30	t->55	v->53	ö->13	
t va	c->3	d->34	g->1	k->4	l->15	n->5	r->162	t->4	
t ve	d->3	m->1	r->48	t->18	
t vi	 ->429	,->6	a->3	d->80	k->119	l->110	n->6	s->71	t->4	
t vo	l->1	r->12	
t vr	a->1	
t vä	c->2	g->6	l->50	n->15	r->14	s->7	x->8	
t vå	g->1	l->2	r->45	
t wo	r->1	
t yp	p->1	
t yt	t->34	
t zo	n->1	
t Ös	t->6	
t äc	k->1	
t äg	a->17	e->1	n->6	
t äm	b->4	n->4	
t än	 ->25	,->1	d->61	n->8	t->2	
t är	 ->874	,->2	.->1	:->1	a->1	e->5	l->1	
t äv	e->39	
t å 	e->3	
t åk	l->1	
t ål	d->1	i->4	ä->2	
t år	 ->22	,->4	.->4	e->1	h->2	l->1	s->1	
t ås	i->1	t->6	
t åt	 ->13	a->9	e->50	f->3	g->10	m->3	n->1	
t åv	i->1	
t öd	e->3	
t ög	o->5	
t ök	a->29	n->1	
t öl	 ->1	
t öm	s->1	
t ön	s->8	
t öp	p->13	
t ös	t->15	
t öv	e->111	r->2	
t! D	e->2	
t! J	a->2	
t! N	ä->1	
t! S	o->1	
t! V	a->1	
t!"J	a->1	
t!(P	a->1	
t!. 	(->1	
t!.(	N->1	
t!De	t->1	
t!Dä	r->1	
t!He	r->3	
t!Ja	g->1	
t!Ku	l->1	
t!Le	d->1	
t!Me	n->1	
t!Nä	r->1	
t!Pr	e->1	
t!Tv	ä->1	
t" (	s->1	
t" g	ö->1	
t" m	e->1	
t" o	c->1	
t" ä	r->1	
t", 	b->1	d->1	e->1	s->1	
t".E	n->1	
t".J	a->1	
t) (	C->1	
t) C	5->1	
t) h	a->2	
t) p	å->1	
t) s	o->1	
t) t	ä->1	
t), 	d->1	s->1	t->1	
t).D	e->1	
t).H	e->2	
t).L	i->1	
t)Nä	s->1	
t, "	e->1	
t, C	o->1	
t, D	a->1	
t, E	G->1	f->1	
t, G	i->1	
t, H	a->1	
t, I	I->2	n->1	
t, J	o->1	
t, L	a->1	
t, O	b->1	
t, P	V->1	
t, S	c->1	o->1	
t, W	e->1	
t, Z	i->1	
t, a	l->1	n->4	r->2	t->30	v->6	
t, b	e->7	l->4	o->1	r->1	y->1	ö->6	
t, c	i->1	
t, d	e->42	i->1	j->1	v->5	ä->9	å->3	
t, e	f->27	l->6	n->19	t->6	x->1	
t, f	a->4	i->2	o->1	r->17	u->1	å->3	ö->39	
t, g	e->4	i->1	l->1	r->1	ä->1	å->5	ö->2	
t, h	a->21	e->21	j->1	o->2	u->1	ä->3	å->1	
t, i	 ->26	n->24	
t, j	a->4	u->3	ä->2	
t, k	a->11	l->1	o->15	r->3	u->3	ä->3	
t, l	a->1	e->1	i->5	ä->2	å->2	
t, m	e->76	i->2	o->2	y->3	ä->1	å->5	
t, n	a->4	ä->16	å->1	
t, o	a->2	b->1	c->110	l->1	m->23	
t, p	a->1	e->1	l->1	o->1	r->4	å->8	
t, r	a->3	e->2	ä->3	å->2	ö->1	
t, s	a->3	e->5	i->2	j->1	k->9	o->55	p->2	t->3	ä->35	å->25	
t, t	.->1	a->3	i->6	o->1	r->5	v->4	y->4	
t, u	n->3	p->2	r->1	t->33	
t, v	a->13	e->2	i->43	o->1	ä->3	å->1	
t, ä	n->2	r->18	v->13	
t, å	 ->1	r->1	t->2	
t, ö	k->1	p->1	
t- o	c->3	
t-Ex	u->1	
t-an	a->5	
t-be	n->5	
t-fr	å->1	
t-st	a->2	
t. (	P->1	
t. 7	 ->1	)->1	
t. A	v->1	
t. D	e->17	ä->1	
t. E	t->1	
t. F	r->1	
t. H	e->1	ä->1	
t. I	 ->1	n->2	
t. J	a->1	
t. K	o->1	
t. M	e->1	
t. O	f->1	
t. S	o->1	
t. V	i->2	å->1	
t. a	i->1	
t.(A	r->1	
t.(F	R->1	
t.(P	T->1	a->1	r->1	
t.)A	n->1	
t.)B	e->2	
t.)F	r->1	
t.)R	e->1	
t.- 	H->1	
t.. 	(->2	
t..(	D->1	
t...	(->1	F->1	
t..H	e->1	
t.19	9->1	
t.Ac	c->1	
t.Al	d->1	l->4	
t.An	s->1	v->1	
t.Ar	a->1	t->1	
t.At	t->2	
t.Av	 ->3	s->6	
t.Be	r->1	t->4	
t.Bi	l->1	
t.Bl	a->1	
t.Bo	r->1	
t.Br	i->1	
t.Bå	d->2	
t.Da	g->1	
t.De	 ->24	l->2	n->35	s->11	t->170	
t.Di	r->3	
t.Dä	r->17	
t.Då	 ->5	
t.EG	-->1	
t.Ef	f->1	t->6	
t.Ek	o->1	
t.En	 ->9	d->3	l->6	
t.Er	f->1	
t.Et	t->6	
t.Eu	r->10	
t.FP	Ö->1	
t.Fe	l->1	
t.Fi	n->1	
t.Fl	e->1	o->1	
t.Fr	a->6	u->10	å->6	
t.Fö	l->2	r->39	
t.Ge	n->4	
t.Gi	v->1	
t.Gr	e->1	u->1	
t.Ha	n->5	
t.He	l->1	r->48	
t.Hi	t->1	
t.Hu	r->4	v->1	
t.Hä	r->7	
t.I 	F->1	N->1	a->3	b->1	d->13	e->2	f->4	k->1	l->1	m->2	n->1	o->1	r->2	s->4	u->1	v->5	ä->1	
t.Ib	l->1	
t.In	g->1	n->1	s->1	t->2	
t.Ja	 ->1	,->2	g->144	
t.Ju	 ->1	s->1	
t.Ko	m->14	n->4	
t.Kr	a->1	
t.Ku	l->2	
t.Kä	r->2	
t.La	 ->1	
t.Li	k->1	t->1	
t.Lä	n->1	
t.Lå	n->1	t->10	
t.Ma	n->14	r->1	x->1	
t.Me	d->11	l->1	n->39	r->1	
t.Mi	l->1	n->12	
t.Mo	r->1	t->3	
t.Må	n->1	
t.Na	t->5	
t.Ni	 ->7	
t.Nu	 ->6	m->1	v->1	
t.Nä	r->10	s->1	
t.Nå	g->1	
t.Nö	d->1	
t.OK	,->1	
t.Ob	e->1	
t.Oc	h->12	
t.Of	f->1	
t.Om	 ->16	
t.Or	d->1	k->1	o->1	
t.PP	E->1	
t.Pa	r->8	
t.Pl	ä->1	
t.Po	r->1	
t.Pr	e->1	o->3	
t.Pu	n->1	
t.På	 ->7	
t.Ra	p->1	
t.Re	d->1	g->1	s->1	
t.Ri	k->1	
t.Rä	t->1	
t.Sa	m->2	n->1	
t.Se	d->1	
t.Sk	a->1	o->1	u->1	
t.Sl	u->6	
t.So	c->1	m->5	
t.St	a->4	o->1	ö->3	
t.Sy	f->1	
t.Så	 ->9	v->1	
t.Ta	c->6	n->1	
t.Th	e->1	
t.Ti	l->4	
t.Tr	e->1	o->2	
t.Tu	s->1	
t.Tv	å->1	
t.Ty	 ->2	v->1	
t.Un	d->3	g->1	i->1	
t.Ur	 ->1	
t.Ut	b->1	f->1	s->1	
t.Va	d->15	l->1	r->7	
t.Vi	 ->84	d->3	l->1	s->2	
t.Vä	s->1	
t.Vå	r->3	
t.ex	.->20	
t.o.	m->7	
t.Än	d->3	
t.Är	 ->1	
t.Äv	e->7	
t.Å 	a->2	e->1	
t.År	 ->1	e->1	
t.Åt	e->1	
t.Ök	a->1	
t.Ös	t->1	
t.Öv	r->1	
t: "	D->2	M->1	a->1	
t: E	f->1	
t: F	r->1	
t: H	o->1	
t: J	a->2	
t: U	n->1	t->1	
t: V	i->1	
t: a	t->1	
t: d	e->5	
t: e	n->1	t->1	
t: f	r->1	ö->1	
t: h	a->1	
t: j	a->2	
t: k	a->1	
t: m	i->1	
t: o	m->2	
t: s	y->1	
t: t	a->1	
t: u	t->1	
t: v	i->1	å->1	
t: ö	n->1	
t; D	a->1	
t; a	l->1	r->1	
t; d	e->5	
t; e	n->1	
t; f	o->1	r->1	
t; u	n->1	
t; å	 ->1	
t? M	e->1	
t? R	å->1	
t?. 	(->2	
t?.(	E->2	
t?An	s->1	
t?At	t->1	
t?Av	 ->1	
t?De	 ->1	t->3	
t?Et	t->1	
t?Eu	r->1	
t?He	r->1	
t?Hu	r->2	
t?I 	v->1	
t?Ja	g->4	
t?Jo	 ->1	
t?Ko	m->1	
t?Kä	r->1	
t?Ne	j->3	
t?Ni	 ->2	
t?Nä	r->1	
t?Oc	h->1	
t?Om	 ->1	
t?RI	N->1	
t?Sk	u->2	
t?Tä	n->1	
t?Ut	g->1	
t?Va	d->1	
t?Vi	 ->1	l->2	s->1	
t?Är	 ->1	
tBet	ä->1	
tJag	 ->1	
tNäs	t->1	
ta -	 ->7	,->1	
ta 1	0->1	
ta A	l->1	m->1	
ta E	G->5	U->1	u->4	
ta F	P->1	
ta J	ö->1	
ta M	a->1	
ta N	a->1	
ta S	h->1	t->1	
ta a	b->1	d->1	k->1	l->7	n->21	r->9	t->47	v->30	
ta b	a->2	e->95	i->11	l->7	o->4	r->2	u->3	ä->1	ö->6	
ta c	e->2	h->1	
ta d	a->4	e->120	i->39	j->1	o->6	r->2	ä->1	ö->1	
ta e	f->6	g->1	k->2	l->4	m->9	n->52	r->11	t->36	v->1	x->1	
ta f	a->22	e->1	i->2	l->2	o->26	r->37	u->3	å->7	ö->142	
ta g	a->2	e->12	i->2	l->1	o->3	r->11	ä->9	å->21	ö->2	
ta h	a->67	e->4	i->3	j->1	o->4	u->3	ä->32	å->2	
ta i	 ->54	d->1	g->3	h->1	n->55	s->1	t->14	
ta j	o->1	u->1	
ta k	a->18	l->4	o->34	r->10	u->1	v->3	ä->5	
ta l	a->8	e->2	i->9	j->1	ä->8	å->1	
ta m	a->8	e->78	i->14	o->11	y->10	ä->2	å->28	ö->21	
ta n	a->14	o->4	u->2	y->5	ä->10	å->4	
ta o	a->1	b->1	c->39	e->1	f->1	g->1	l->4	m->74	n->1	r->13	s->13	
ta p	a->42	l->3	o->6	r->48	u->38	å->49	
ta r	a->17	e->35	i->6	u->2	ä->1	å->3	ö->4	
ta s	a->47	e->10	i->44	j->2	k->37	l->13	m->3	n->1	o->23	p->6	t->59	v->2	y->11	ä->25	å->4	
ta t	a->11	e->6	i->32	j->1	o->6	r->2	u->1	v->4	y->4	å->1	
ta u	n->7	p->76	r->4	t->29	
ta v	a->23	e->6	i->32	o->1	ä->4	å->5	
ta y	t->2	
ta Ö	s->2	
ta ä	g->6	m->3	n->12	r->169	v->4	
ta å	r->5	s->1	t->18	
ta ö	k->4	v->12	
ta!D	e->1	
ta!F	r->1	
ta, 	a->5	b->1	d->3	e->4	f->9	h->6	i->4	j->1	k->2	l->1	m->9	o->18	r->2	s->6	t->3	u->6	v->2	
ta. 	D->1	F->1	V->1	
ta.(	P->1	
ta.)	F->1	
ta.-	 ->1	
ta..	 ->1	(->1	
ta.A	n->1	
ta.B	e->2	
ta.C	o->1	
ta.D	e->26	ä->1	å->1	
ta.E	f->3	m->1	n->2	
ta.F	r->1	ö->2	
ta.G	e->1	
ta.H	e->4	
ta.I	 ->5	n->2	
ta.J	a->12	
ta.K	o->1	
ta.M	e->7	
ta.N	u->1	ä->1	
ta.O	c->2	m->2	
ta.P	r->2	å->1	
ta.S	e->1	i->1	j->1	o->1	t->2	å->1	
ta.T	o->1	r->1	
ta.V	a->4	i->11	å->1	
ta.Ä	r->1	
ta: 	I->1	J->2	V->1	u->1	v->1	
ta; 	d->1	v->1	
ta?D	e->1	
ta?J	a->1	
ta?N	ä->1	
ta?V	i->1	
taNä	s->1	
taaf	f->1	
tab 	s->1	
taba	s->1	
tabe	h->1	l->37	
tabi	l->24	
tabl	a->13	e->13	
tabr	i->3	
tabu	 ->1	l->1	
tack	 ->29	,->1	.->2	a->105	e->1	l->1	o->1	s->9	
tad 	a->1	f->6	m->3	o->3	p->2	s->1	ö->1	
tad,	 ->2	
tad.	"->1	(->1	D->1	F->1	H->3	J->1	M->2	O->14	R->1	
tade	 ->64	,->3	.->3	l->2	s->14	
tadg	a->28	o->1	
tadi	e->4	u->4	
tadk	o->24	
tadm	i->2	
tads	b->1	c->1	o->1	p->1	
tadt	,->1	
tafr	å->10	
tag 	a->3	b->1	e->2	f->5	g->1	h->5	i->11	k->4	l->2	n->1	o->7	p->3	s->21	t->1	u->1	v->2	ä->3	
tag,	 ->20	
tag.	A->1	D->4	E->2	F->1	I->3	J->1	K->2	M->1	O->1	R->1	S->1	T->1	V->2	
tag?	F->1	
taga	n->102	r->70	
tagb	a->15	
tage	l->1	n->68	t->22	
tagi	t->100	
tagl	i->5	
tagn	a->10	e->9	i->4	
tags	 ->3	a->4	b->1	e->5	f->3	g->2	i->1	j->2	k->1	l->1	m->1	n->1	r->5	s->3	t->2	
tain	,->1	e->1	s->24	
tak 	f->1	
tak,	 ->2	
taka	 ->5	
take	l->2	t->1	
takl	a->1	
takt	 ->8	.->2	e->12	i->4	
taku	l->1	
tal 	-->1	a->4	b->5	d->1	e->1	f->9	h->2	i->13	k->4	l->2	m->21	n->1	o->13	p->4	r->5	s->22	t->4	u->2	v->1	ä->3	å->1	ö->3	
tal"	 ->1	
tal,	 ->6	
tal-	F->3	
tal.	D->1	E->1	F->1	H->2	I->1	J->1	K->2	S->1	V->1	
tal:	 ->1	
talF	i->1	
tala	 ->109	"->1	,->3	.->6	?->3	d->35	n->57	r->118	s->11	t->32	
talb	e->1	l->1	
tale	n->15	s->4	t->61	
talf	å->4	ö->1	
tali	e->36	g->2	n->2	s->2	t->3	
talj	 ->2	,->2	.->1	a->1	e->26	f->1	k->2	
tall	,->1	d->1	e->9	i->1	k->2	
talm	a->418	
taln	i->15	
talo	g->2	
talr	i->4	
tals	 ->20	.->1	f->1	k->4	l->1	p->7	r->1	s->1	u->1	
talt	 ->6	.->1	e->1	s->1	
talv	o->1	
taly	s->2	
tame	-->1	n->8	
tami	n->2	
tamp	 ->1	
tan 	1->3	I->1	a->67	b->7	d->33	e->17	f->11	g->3	h->9	i->10	j->1	k->12	m->10	n->10	o->48	p->18	r->5	s->17	t->37	u->4	v->7	ä->36	ö->6	
tan,	 ->10	
tan.	(->2	A->1	D->1	F->1	H->1	J->4	M->1	S->1	T->1	U->1	V->3	
tan;	 ->1	
tan?	Ä->1	
tana	 ->1	
tanb	u->1	
tand	a->25	e->158	
tane	n->3	r->5	
tanf	ö->32	
tank	-->1	a->16	e->69	f->8	r->7	
tann	a->10	i->14	
tano	 ->1	
tans	 ->13	,->6	.->1	?->1	e->8	k->6	l->1	r->22	v->13	
tant	 ->2	,->1	e->12	i->3	
tanv	ä->1	
tapo	l->1	
tapp	 ->1	a->3	e->4	
tar 	A->1	E->1	F->1	a->21	b->12	d->28	e->20	f->18	g->5	h->5	i->29	j->11	k->6	l->1	m->28	n->7	o->24	p->24	r->2	s->30	t->33	u->19	v->17	y->1	ä->2	ö->3	
tar,	 ->6	
tar.	D->3	F->1	J->1	M->1	V->2	Ä->1	
tarb	e->32	
tare	 ->31	,->6	.->3	n->8	r->21	
tarh	u->1	
tari	a->2	k->9	n->1	s->23	t->3	u->1	
tark	 ->11	,->1	a->25	e->1	l->1	t->23	
tarl	ø->2	
tarm	a->10	
tarn	a->19	
tart	a->11	e->4	p->1	
tarv	l->1	
tas 	a->24	b->5	c->1	d->8	e->9	f->9	g->3	h->1	i->28	j->1	k->2	l->3	m->13	n->6	o->7	p->9	r->1	s->12	t->2	u->20	v->9	ä->3	
tas,	 ->10	
tas.	 ->1	B->1	D->1	F->1	J->3	O->1	P->3	V->3	Ä->1	
tasi	e->1	f->1	n->1	
task	 ->1	
tasp	e->2	
tast	 ->1	e->1	i->9	r->90	
tasä	k->1	
tat 	-->2	a->16	b->4	d->9	e->11	f->19	g->2	h->9	i->12	k->2	l->3	m->12	n->1	o->18	p->6	r->1	s->27	t->3	u->6	v->6	ä->2	å->1	
tat,	 ->16	
tat.	 ->2	B->1	D->8	E->2	G->1	H->2	I->3	J->4	K->2	L->1	O->2	P->1	T->1	
tat:	 ->2	
tat?	.->1	J->1	
tate	 ->2	n->42	r->341	t->29	
tati	n->1	o->33	s->9	v->15	
tatl	i->101	
tato	r->1	
tats	 ->38	,->2	-->5	.->3	b->2	k->1	m->4	n->4	p->1	s->19	
tatt	a->8	
tatu	e->2	r->3	s->8	
tatö	v->6	
tatü	r->1	
taue	n->1	
taun	i->3	
taur	e->1	
tav 	o->1	ö->1	
tavl	a->7	i->1	
tax-	f->3	
taxe	r->1	
tbal	a->2	
tban	k->4	
tbar	h->1	t->2	
tbas	i->1	u->1	
tbef	o->2	
tbeh	o->1	
tbes	t->4	
tbet	a->7	
tbev	a->1	
tbil	d->65	
tblo	c->1	
tbok	 ->12	,->1	.->5	e->35	
tbol	l->1	
tbra	n->1	
tbre	d->4	
tbri	n->1	
tbud	 ->3	s->1	
tbur	e->1	
tbyg	g->3	
tbyt	a->1	e->16	
tc. 	o->1	Ä->2	
tc.D	e->1	
tc.E	n->1	
tc?A	t->1	
tcha	n->1	
tche	r->1	
tdel	a->1	n->2	
tdem	o->11	
tder	a->1	
tdik	t->1	
tdir	e->1	
te (	K->2	
te -	 ->8	,->1	
te 1	9->1	
te B	e->1	
te E	M->1	U->2	k->1	u->8	
te F	N->1	o->1	
te I	s->1	
te J	o->1	
te O	u->1	
te Q	u->1	
te a	b->1	c->11	g->1	k->1	l->42	n->29	r->5	s->2	t->76	u->4	v->25	
te b	a->91	e->55	i->2	l->29	o->3	r->2	y->1	ä->2	ö->10	
te c	e->1	h->2	o->2	
te d	a->5	e->93	i->3	o->5	r->3	ä->14	å->3	ö->2	
te e	f->2	k->1	l->3	m->1	n->44	p->1	r->8	t->12	u->2	v->1	x->5	
te f	a->18	e->2	i->24	o->10	r->14	u->7	y->1	ä->1	å->30	ö->86	
te g	a->6	e->30	i->1	j->3	l->10	o->9	r->4	ä->4	å->19	ö->30	
te h	a->110	e->50	i->3	j->2	o->4	u->3	ä->6	å->5	ö->6	
te i	 ->47	a->2	f->3	g->1	l->1	n->46	s->1	
te j	a->9	o->1	u->3	ä->1	
te k	a->59	l->3	n->1	o->49	r->9	u->18	v->2	ä->4	ö->1	
te l	a->3	e->10	i->4	u->1	y->7	ä->39	å->8	ö->7	
te m	a->24	e->63	i->22	o->6	y->5	å->15	ö->7	
te n	a->4	e->2	i->4	o->5	u->7	ä->5	å->28	ö->11	
te o	b->1	c->49	f->2	l->2	m->28	p->2	r->3	
te p	a->4	e->12	l->2	o->2	r->7	u->2	å->52	
te r	a->12	e->33	i->2	u->1	ä->14	å->11	ö->2	
te s	a->13	e->25	i->2	j->6	k->61	l->3	n->5	o->31	p->2	t->22	v->4	y->7	ä->25	å->13	ö->4	
te t	a->49	e->4	i->52	j->1	o->1	r->6	u->3	v->2	y->2	ä->8	
te u	n->12	p->39	r->1	t->40	
te v	a->61	e->13	i->82	o->2	ä->9	å->3	
te ä	g->3	n->17	r->76	v->5	
te å	l->1	r->16	s->1	t->11	
te ö	k->4	n->2	p->2	v->14	
te!D	e->1	
te!M	e->1	
te, 	a->4	d->2	e->2	f->2	g->1	h->2	i->1	k->2	l->1	m->2	n->1	o->6	p->1	r->1	s->2	v->5	ä->3	
te- 	o->1	
te-L	e->1	
te. 	D->1	
te..	 ->1	
te.A	k->1	n->1	
te.B	e->1	
te.D	e->9	ä->1	
te.F	r->1	ö->2	
te.H	e->3	
te.I	 ->1	
te.J	a->5	
te.K	o->1	
te.L	i->1	ä->1	å->1	
te.M	a->1	e->2	
te.N	i->1	
te.O	m->1	
te.P	å->1	
te.R	e->1	å->1	
te.S	o->1	å->1	
te.U	p->1	
te.V	a->1	i->4	å->1	
te.Å	 ->1	r->1	t->1	
te: 	V->1	v->1	
te?F	ö->1	
te?H	u->1	ä->1	
te?I	 ->1	
te?S	o->1	
teat	e->1	
teau	 ->1	,->2	
teba	s->1	
tebe	s->2	t->12	
tebo	r->1	
teck	e->15	n->32	
tede	l->3	
tedt	 ->2	,->2	
teen	d->3	h->5	
teer	i->1	
tefe	l->1	
tefr	i->1	å->2	
tefö	r->6	
teg 	a->1	b->1	f->11	g->1	h->2	i->13	j->1	l->2	m->4	n->2	o->2	p->3	s->7	t->3	u->1	v->1	
teg,	 ->3	
teg.	D->2	
tege	n->5	t->2	
tegi	 ->17	,->3	.->3	e->14	n->8	p->1	s->17	
tego	r->8	
tegr	a->16	e->23	i->3	
tegå	n->1	
tein	.->1	c->1	s->1	
teke	n->2	
tekn	i->49	o->3	
teko	n->1	
tekt	i->4	
tel 	2->1	4->1	i->3	o->1	
tela	 ->1	,->1	
tele	f->1	k->3	n->1	v->2	
teli	g->1	
tell	-->3	a->1	b->2	e->4	f->3	i->8	m->1	r->4	t->1	
teln	 ->1	
tels	e->31	
telt	.->1	
telä	m->3	t->1	
tem 	-->1	a->3	d->3	e->1	f->21	g->1	i->5	k->2	m->10	o->7	p->3	s->16	ä->1	ö->1	
tem,	 ->9	
tem.	 ->1	D->3	E->1	G->1	H->2	M->1	T->1	U->1	
tem:	 ->1	
tema	,->1	l->1	n->5	t->12	
temb	e->15	
teme	n->21	t->69	
temo	t->27	
temp	e->4	o->2	
temä	n->37	
ten 	(->1	-->10	1->2	A->3	B->2	I->3	L->1	P->1	R->1	S->1	a->133	b->10	d->11	e->12	f->89	g->22	h->30	i->88	j->1	k->21	l->3	m->42	n->9	o->111	p->35	r->4	s->63	t->27	u->15	v->30	ä->32	å->6	ö->9	
ten!	 ->4	
ten"	 ->1	.->3	
ten)	 ->3	
ten,	 ->112	
ten.	 ->2	"->1	A->4	D->45	E->8	F->9	H->9	I->4	J->16	K->6	L->1	M->11	N->4	O->11	P->1	R->1	S->9	T->3	U->1	V->17	Ä->1	Å->2	Ö->1	
ten:	 ->2	
ten;	 ->2	
ten?	J->1	K->1	
tenF	r->1	
tenH	e->1	
tenN	ä->1	
tena	 ->7	r->3	
tenb	e->4	
tend	a->1	e->14	r->1	ö->1	
tene	n->1	r->18	
tenf	ö->2	
tenh	e->3	
tenk	o->1	
tenl	ö->1	
tenp	r->1	
tenr	e->2	
tens	 ->72	,->4	.->2	b->1	e->1	i->12	k->72	
tent	 ->3	a->7	i->7	
tenv	ä->8	
teor	e->2	
tepo	l->1	
tepr	o->1	
ter 	(->1	-->14	1->1	A->2	B->2	C->1	E->6	F->1	G->6	H->1	J->1	K->1	L->1	M->2	O->2	S->2	T->2	a->109	b->16	d->62	e->38	f->68	g->13	h->28	i->80	j->9	k->23	l->9	m->49	n->8	o->133	p->34	r->9	s->145	t->40	u->18	v->32	Ö->1	ä->29	å->6	ö->12	
ter!	 ->12	J->1	M->1	V->1	
ter"	 ->1	,->1	
ter)	 ->2	
ter,	 ->114	
ter-	b->1	k->1	n->1	
ter.	 ->4	)->1	.->1	A->1	B->1	D->35	E->12	F->11	H->4	I->3	J->21	K->4	L->3	M->8	N->3	O->4	P->4	S->6	T->6	U->1	V->15	Ä->3	Å->2	
ter:	 ->3	
ter;	 ->2	
ter?	B->1	D->1	H->1	T->1	
terH	e->1	
tera	 ->191	,->5	.->16	d->48	l->8	n->43	r->111	s->64	t->51	
terb	e->3	i->1	
terd	a->41	ö->1	
tere	r->1	
terf	a->1	i->5	r->8	u->2	ö->11	
terg	a->2	e->4	i->8	r->1	å->1	
terh	a->5	ä->2	å->2	
teri	 ->1	a->23	e->28	g->19	l->1	m->8	n->96	s->2	
terk	o->7	r->1	
terl	e->3	i->56	y->2	ä->3	
term	e->3	i->9	ö->2	
tern	 ->26	,->2	.->9	/->2	a->652	e->11	f->1	i->1	s->5	t->4	
tero	m->1	
terp	a->1	o->2	r->1	
terr	a->2	e->5	i->147	o->10	å->14	
ters	 ->13	-->1	a->4	e->1	k->5	o->190	p->3	t->72	
tert	 ->2	a->12	r->2	ä->1	
teru	p->34	
terv	e->8	i->66	j->3	u->2	ä->4	
terå	t->1	
tes 	3->1	a->4	e->1	i->6	m->2	t->1	u->1	
tes,	 ->1	
tes-	 ->1	
tes.	F->1	K->1	O->1	V->1	
tesa	t->1	
tese	k->2	n->1	
tesg	å->3	
tesi	s->3	
tesl	u->17	ö->2	
tess	 ->4	b->5	e->2	h->1	
test	 ->3	,->1	a->2	e->6	ä->4	å->1	
tesy	s->1	
tet 	(->1	,->1	-->7	1->2	K->1	M->1	a->105	b->20	c->2	d->16	e->10	f->159	g->17	h->40	i->73	j->3	k->31	l->9	m->59	n->6	o->108	p->15	r->5	s->54	t->13	u->9	v->17	ä->27	å->1	
tet!	H->1	
tet"	,->1	.->1	
tet,	 ->91	
tet-	 ->1	
tet.	 ->1	)->3	.->1	B->1	D->27	E->4	F->7	H->7	I->3	J->15	K->3	L->1	M->4	N->1	P->1	R->1	S->3	T->1	V->9	Ä->1	
tet:	 ->4	
tet?	D->1	H->2	N->1	Ä->1	
tete	n->56	r->20	
teti	s->2	
tets	 ->116	-->1	a->2	b->3	f->2	g->1	h->2	k->3	n->1	o->1	p->19	r->3	s->2	
teur	o->9	
text	 ->12	,->5	.->1	e->27	
tfal	l->7	
tfar	a->89	t->1	
tfas	n->3	
tfat	t->2	
tfed	e->1	
tfla	g->1	
tfle	r->1	
tfli	r->1	
tfly	t->1	
tfor	m->41	s->1	
tfra	m->1	
tfrå	g->16	
tful	l->15	
tfäl	l->8	
tfär	d->20	
tfäs	t->2	
tfån	g->1	
tföl	j->12	
tför	 ->46	a->18	b->1	d->7	e->1	f->2	k->7	l->4	o->6	s->5	t->13	ä->4	
tgav	s->1	
tgic	k->1	
tgif	t->16	
tgil	t->8	
tgiv	i->1	n->1	
tgjo	r->4	
tgru	p->7	
tgär	d->245	
tgå 	e->1	f->2	t->1	
tgå.	D->1	N->1	
tgåe	n->14	
tgån	g->18	
tgår	 ->8	
tgåv	o->1	
tgör	 ->46	,->1	.->1	a->13	s->2	
th S	c->1	
th h	a->1	
th n	ä->1	
th o	c->1	
th, 	o->1	
th-B	e->7	
than	d->1	t->1	
thar	 ->2	"->1	
thav	a->1	
the 	R->1	c->1	i->1	
then	 ->3	,->1	s->2	
ther	"->1	a->1	
thet	 ->2	.->1	e->1	s->1	
thie	s->2	
thom	 ->3	
thu 	o->1	
thus	e->3	g->4	
thy 	o->1	
thäl	s->1	
thär	d->4	
thål	l->11	
thör	a->1	
ti -	 ->1	
ti a	n->1	
ti d	e->2	
ti f	r->1	ö->9	
ti g	j->1	
ti h	a->3	e->1	
ti i	 ->5	g->1	n->3	
ti k	o->2	r->1	
ti m	e->2	
ti o	c->11	m->1	
ti p	å->2	
ti s	n->1	o->7	å->1	
ti t	i->2	
ti u	p->1	
ti v	a->1	
ti å	t->1	
ti! 	J->2	U->1	
ti" 	s->1	
ti, 	M->1	b->1	d->2	e->1	k->1	l->1	m->1	o->1	p->1	s->2	ä->2	
ti-g	e->1	
ti-i	r->1	
ti-r	a->1	
ti..	.->1	
ti.D	e->3	
ti.E	f->1	n->1	
ti.F	o->1	
ti.H	a->1	e->1	ä->1	
ti.I	 ->1	
ti.J	a->1	
ti.K	a->1	u->1	
ti.M	i->1	
ti.V	i->1	
tial	 ->1	,->1	.->1	
tian	 ->1	
tiat	i->80	
tibe	d->1	t->10	
tica	l->1	
tice	 ->4	
tich	e->1	
tick	 ->1	e->1	p->3	
tid 	E->1	a->29	b->11	c->1	d->10	e->8	f->18	g->3	h->16	i->14	j->1	k->9	l->3	m->7	n->5	o->7	p->4	r->2	s->16	t->8	u->2	v->6	y->1	ä->11	å->3	
tid,	 ->16	
tid.	.->1	D->5	F->1	K->1	M->1	N->1	O->1	S->1	T->2	V->1	
tid:	 ->1	
tida	 ->23	
tide	m->1	n->118	r->5	
tidi	g->152	
tidl	i->4	
tidn	i->6	
tidp	u->10	
tids	a->4	b->2	d->4	f->11	g->1	i->2	m->2	o->1	p->15	r->7	s->2	å->3	ö->1	
tidt	a->6	
tie-	 ->1	
tieb	ö->1	
tied	e->2	
tiel	f->1	l->10	
tiem	i->3	
tien	t->4	
tier	 ->17	,->2	a->3	i->4	n->12	
tiet	 ->6	)->4	,->4	n->3	s->16	
tieu	r->1	
tieä	g->2	
tifa	s->3	
tifi	c->15	e->16	k->4	q->1	
tifo	l->1	n->2	
tifr	å->18	
tift	a->15	n->113	
tig 	-->2	b->3	d->7	e->1	f->20	g->3	h->3	i->4	j->1	k->5	l->3	m->5	o->11	p->10	r->12	s->4	t->5	u->5	å->3	ö->2	
tig,	 ->8	
tig.	D->4	I->1	J->3	M->2	N->1	
tig?	J->1	
tiga	 ->131	,->6	.->3	d->10	n->2	r->17	s->48	t->10	
tigd	o->12	
tige	r->4	
tigg	e->1	
tigh	e->182	
tigi	t->2	
tigl	i->4	
tigm	a->1	
tigt	 ->167	,->17	.->13	
tiho	p->1	
tiin	t->1	
tik 	-->2	J->1	a->5	e->3	f->19	h->4	i->7	k->3	m->11	n->1	o->28	p->2	r->2	s->28	t->1	u->2	v->3	ä->4	ö->1	
tik!	O->1	
tik"	 ->1	
tik,	 ->31	
tik.	.->1	D->8	E->2	F->2	H->3	I->1	J->1	M->1	R->2	T->1	V->2	Ä->1	
tik?	H->1	V->1	
tika	 ->3	b->1	f->1	l->3	n->1	p->1	s->1	
tike	l->95	n->144	r->16	
tikl	a->15	
tiko	l->1	m->6	
tikr	a->1	y->2	
tiks	 ->1	
til 	-->1	m->1	n->1	
tila	t->1	
tile	d->1	r->1	
tili	s->1	
till	 ->1737	!->1	,->17	.->14	:->1	?->3	a->1	b->56	d->13	e->3	f->143	g->49	h->53	k->15	m->5	n->6	r->77	s->127	t->11	v->114	ä->194	å->45	
tima	 ->5	,->1	.->1	l->3	t->1	
time	r->5	t->1	
timi	s->4	t->6	
timm	a->6	e->5	
timt	 ->3	,->1	
timu	l->11	
timö	g->1	
tin 	a->2	b->1	f->2	h->1	i->1	m->1	o->3	s->3	v->1	
tin,	 ->2	
tin.	A->1	F->2	H->1	O->1	
tina	 ->6	-->1	f->2	s->1	t->5	
tind	u->2	
tine	n->6	r->6	z->1	
ting	 ->62	,->4	.->4	a->12	e->13	f->1	
tini	e->4	
tink	t->3	
tinm	ä->1	
tinn	e->1	o->1	
tino	s->4	t->1	
tinr	i->2	
tins	 ->5	k->8	
tinu	e->2	
tinv	e->1	
tio 	f->1	g->3	m->2	s->1	ä->1	å->7	
tioe	l->1	
tiof	e->1	
tion	 ->245	"->1	,->36	.->57	:->3	;->1	?->3	a->46	d->1	e->760	i->5	s->96	
tiop	i->3	
tios	j->1	
tiot	a->6	u->1	
tipe	n->1	
tipr	o->2	
tiqu	e->2	
tire	f->1	
tis 	d->1	e->1	i->1	r->1	t->1	u->1	å->1	
tis,	 ->1	
tis.	D->1	
tisd	a->2	
tise	k->2	m->3	r->17	
tish	 ->1	
tisk	 ->101	,->2	-->1	.->7	a->316	t->161	
tism	 ->2	,->2	.->3	
tisp	l->1	
tist	i->9	
tisy	s->1	
tit 	a->2	e->1	f->1	m->1	s->2	
tita	t->4	
tite	l->1	t->8	
titi	e->6	o->1	
titr	u->1	
tits	 ->8	
titt	 ->2	a->20	
titu	e->1	t->158	
tity	d->5	
tiv 	(->1	-->3	9->8	E->1	a->6	b->2	d->4	e->7	f->16	g->1	h->8	i->13	k->10	l->7	m->5	o->30	p->8	r->3	s->45	t->15	u->3	v->6	ä->6	å->2	ö->1	
tiv,	 ->23	
tiv.	 ->1	.->1	A->1	B->1	D->5	E->1	F->4	I->2	L->1	M->1	O->1	R->1	S->1	V->1	Y->1	
tiv:	 ->2	
tiv;	 ->1	
tiv?	F->1	N->1	
tiva	 ->105	,->4	.->3	n->1	r->11	s->1	t->1	v->7	
tivb	e->1	
tive	 ->15	n->12	r->17	t->100	
tivf	ö->4	
tivi	s->4	t->38	
tivl	i->2	
tivr	i->1	ä->4	
tivt	 ->100	,->7	.->7	
tiös	 ->2	,->1	a->8	t->1	
tja 	a->5	c->1	d->5	i->1	o->1	s->5	
tjad	e->4	
tjan	d->9	
tjar	 ->3	
tjas	 ->6	
tjat	 ->1	a->1	
tjoc	k->2	
tjug	o->4	
tjus	t->1	
tjäm	n->5	t->3	
tjän	a->21	s->123	t->29	
tjär	a->1	n->2	
tkan	t->1	
tkas	t->15	
tkat	e->1	
tkla	s->1	
tkom	.->1	m->18	p->1	s->1	
tkon	c->1	k->1	t->16	
tkos	t->2	
tkra	v->1	
tkri	g->1	
tkrä	v->3	
tkub	i->1	
tkus	t->2	
tkvä	l->1	
tkäl	l->1	
tköt	t->3	
tlag	t->1	
tlan	d->15	t->6	
tle 	o->2	ä->1	
tle.	V->1	
tlek	t->1	
tler	 ->3	,->1	-->1	s->1	
tlev	n->1	
tlig	 ->64	,->1	.->4	?->1	a->188	e->137	g->17	h->37	t->81	
tlin	j->76	
tlis	t->2	
tlov	a->3	
tläg	g->4	
tläm	n->2	
tlän	d->15	n->1	
tlåt	a->2	
tlös	.->1	a->1	h->2	t->1	
tmak	t->1	
tman	a->1	i->21	
tmar	g->1	k->1	
tmat	c->1	
tmed	e->1	l->1	
tmer	 ->1	
tmin	s->27	
tmis	s->1	
tmon	n->1	
tmyn	d->3	n->1	
tmän	g->2	
tmär	k->32	
tmäs	s->1	
tmät	i->1	
tmål	s->1	
tna 	a->1	b->2	d->2	e->1	f->1	h->1	i->1	m->1	o->18	p->1	s->1	t->4	v->1	
tna,	 ->3	
tna.	 ->2	D->1	E->1	S->1	U->1	
tnad	 ->10	.->1	;->1	e->75	s->22	
tnar	 ->8	
tnas	 ->2	.->1	
tne 	o->1	t->1	
tnen	 ->1	,->1	.->1	
tner	 ->7	.->1	?->1	n->1	s->18	
tnes	s->1	
tnet	 ->4	.->2	
tnin	g->648	
tnis	k->14	
tnju	t->1	
tnyt	t->42	
tnäm	n->8	
tnät	 ->1	
to -	 ->1	
to a	c->1	
to f	ö->3	
to h	a->1	å->1	
to i	 ->1	
to k	a->1	
to o	c->1	m->1	
to s	a->1	å->1	
to t	i->1	
to v	i->1	
to ö	p->1	
to-a	n->1	
to-p	r->1	
to.J	a->1	
to.V	i->1	
to/O	i->1	
toak	t->1	
toan	a->1	
toba	k->2	s->1	
tobe	r->8	t->1	
tock	h->3	
tod 	a->4	b->1	d->2	e->2	f->3	i->1	j->1	m->3	n->1	p->2	s->6	ä->1	å->1	
tode	n->4	r->12	
todo	n->1	
tog 	1->1	b->1	d->3	e->4	h->2	i->3	k->3	l->5	m->2	n->1	o->2	p->1	r->4	s->1	u->9	
toga	m->2	
toge	n->2	
togs	 ->20	,->2	
toko	l->26	
tol 	b->1	d->1	i->1	o->1	s->2	v->1	
tol.	D->1	E->1	
tola	r->25	
tole	n->46	r->18	
toli	k->4	
tolk	a->12	n->14	
tolp	e->1	
tols	a->1	b->1	f->2	k->4	p->1	s->1	t->1	u->1	v->1	
tolt	 ->6	a->3	h->2	
tolv	 ->1	
tom 	P->1	a->15	b->9	d->4	e->2	f->7	g->3	h->4	i->5	k->8	m->7	n->2	o->5	p->3	r->4	s->6	t->4	v->5	ä->5	
tom!	T->1	
tom)	 ->1	
tom,	 ->5	
tom.	V->1	
toma	t->8	
tome	n->3	u->3	
tomf	o->1	
tomm	a->1	
tomo	r->7	
tomr	u->2	å->6	
toms	t->2	
ton 	5->1	a->3	f->3	i->3	k->1	m->9	o->5	p->1	s->3	t->1	v->1	å->2	
ton,	 ->1	
ton-	H->1	
ton.	 ->1	H->1	V->1	
ton/	å->2	
ton?	 ->1	
tona	 ->26	d->6	r->7	s->1	t->6	
tond	e->3	
tone	 ->27	n->1	r->2	
tong	i->1	
tonh	u->1	
toni	n->1	
tons	 ->4	
tonv	i->4	
tonå	r->1	
top-	s->1	
topi	l->1	
topp	 ->8	a->10	e->3	m->10	
topr	o->2	
tor 	a->5	b->16	c->1	d->14	e->4	f->9	g->2	h->6	i->4	j->2	k->3	l->1	m->12	o->7	p->3	r->6	s->7	t->3	u->16	v->4	ä->1	ö->1	
tor,	 ->10	
tor.	A->1	D->1	J->3	O->1	R->1	T->1	
tora	 ->153	,->2	.->3	?->1	t->18	
torb	r->15	
torc	y->4	
tord	e->1	r->2	
tore	 ->1	n->1	r->42	t->1	
torf	ö->2	
torg	a->1	
torh	a->1	e->1	
tori	a->10	e->20	k->4	n->10	s->33	t->5	u->10	
tork	a->2	n->1	
torl	ä->1	
torm	 ->1	,->1	a->20	e->6	f->1	
torn	 ->22	)->1	,->12	.->10	?->1	a->4	e->1	s->4	
torp	e->2	o->1	
tors	 ->1	a->1	d->8	i->1	k->3	l->2	ö->1	
tort	 ->41	a->1	e->1	y->1	
torv	e->4	
tos 	b->9	e->1	f->1	k->1	o->1	v->1	
tota	l->34	
town	 ->2	,->1	
toxi	s->1	
tpar	t->9	
tpek	a->1	
tpen	s->1	
tper	i->10	
tpla	n->3	t->1	
tplå	n->2	
tpol	i->3	
tpos	t->10	
tpra	t->1	
tpre	s->1	
tpri	o->1	
tpro	b->1	g->1	j->1	t->1	
tprä	g->1	
tpun	k->3	
tra 	A->1	E->3	F->1	J->1	T->1	a->1	b->2	c->1	d->13	f->4	g->3	h->1	i->2	k->7	l->2	m->5	o->4	p->1	r->1	s->13	t->3	u->1	v->1	ö->1	
tra,	 ->1	
trad	 ->5	e->2	i->19	
traf	f->41	i->9	
trag	e->4	i->6	
trak	a->1	o->5	t->30	
tral	 ->7	-->6	.->2	a->20	b->8	e->2	f->1	i->26	t->7	
tram	 ->1	n->2	p->2	
tran	 ->1	d->37	s->113	
trao	r->1	
trap	e->1	p->1	r->1	
trar	 ->21	,->3	.->1	:->1	n->6	s->1	
tras	 ->8	.->2	a->1	b->5	m->1	s->1	t->2	
trat	 ->3	e->63	i->44	s->2	
trau	m->1	
trav	a->1	e->1	
trax	 ->3	
tre 	a->10	b->3	d->2	e->1	f->13	g->6	h->1	i->2	k->10	l->1	m->20	o->11	p->3	r->5	s->22	t->6	u->1	v->6	ä->6	å->3	ö->1	
tre,	 ->5	
tre.	E->1	I->1	J->2	P->1	T->1	
tre:	 ->1	
trea	 ->1	l->2	m->8	
trec	k->1	
tred	a->3	d->1	j->72	n->4	
treg	e->1	i->1	
trek	l->1	
trel	a->1	
trem	a->2	h->14	i->10	t->4	å->1	
tren	d->1	
trep	r->5	
trer	a->28	i->3	
tres	 ->3	s->120	u->3	
tret	 ->2	a->1	t->5	
trev	l->3	
tri 	b->1	d->1	i->1	o->2	s->6	
tri,	 ->3	
tri-	 ->1	
trib	u->1	
tric	h->6	i->1	
trid	 ->9	a->2	d->2	e->8	i->1	l->1	
trie	l->6	r->2	
trif	r->4	
trik	e->19	t->25	
tril	i->1	j->1	o->1	
trin	 ->39	!->1	,->15	.->14	:->1	?->1	g->24	s->9	
trio	 ->1	t->1	
trip	o->2	
tris	 ->3	
tro 	a->4	d->1	m->1	n->2	p->2	t->1	ä->1	
tro.	V->1	
troa	k->12	
trod	d->3	u->6	
troe	n->58	
trof	 ->24	,->4	.->4	a->1	d->1	e->51	h->1	s->4	
trog	e->2	
troj	k->1	
trol	,->1	.->1	e->1	i->11	l->178	
tron	 ->1	i->9	o->4	
trop	a->2	
tror	 ->150	,->1	
tros	 ->2	
trot	a->2	n->2	s->46	t->4	
trou	x->1	
trov	e->4	i->1	ä->14	
true	r->5	
truk	i->1	t->186	
trum	 ->6	!->1	,->2	e->54	
trun	t->4	
trup	p->3	
trus	t->9	
trut	t->1	
tryc	k->101	
tryg	g->8	
tryk	.->1	a->29	e->2	s->2	
trym	m->11	
tryp	s->1	
trä 	u->1	ö->1	
träc	k->32	
träd	 ->4	,->1	.->1	a->78	d->10	e->65	s->2	
träf	f->117	
trän	d->2	g->66	i->1	
träp	r->1	
träs	k->1	
trät	o->1	t->14	
träv	a->31	i->1	
tråd	a->3	e->1	
tråe	t->1	
tråk	i->3	
trål	k->1	n->3	s->1	
trån	g->2	
trög	h->1	
tröj	o->1	
trök	 ->1	,->1	s->1	
tröm	 ->4	,->1	:->1	m->7	n->6	
trös	k->3	t->1	
tröt	t->2	
ts "	B->1	g->1	
ts (	u->1	
ts -	 ->9	
ts 8	0->1	
ts B	a->1	
ts E	u->1	
ts L	e->1	
ts S	p->2	
ts a	b->1	l->15	m->2	n->9	r->6	t->23	u->1	v->69	
ts b	e->28	i->2	o->1	u->2	ä->1	
ts c	e->1	o->1	
ts d	e->31	i->14	o->2	ä->3	
ts e	f->3	g->2	l->3	n->6	r->1	t->1	x->1	
ts f	a->3	e->1	i->1	j->1	l->1	o->2	r->30	u->2	å->3	ö->57	
ts g	e->17	i->3	o->1	r->15	å->1	ö->2	
ts h	a->3	i->4	j->1	o->2	u->1	ä->10	å->2	
ts i	 ->48	k->1	n->15	
ts k	a->1	l->3	o->4	r->3	u->1	ä->1	
ts l	a->2	e->7	i->2	o->2	ö->1	
ts m	a->1	e->23	i->4	o->5	y->1	å->3	ö->5	
ts n	e->4	u->2	y->2	ä->1	å->3	
ts o	c->39	h->1	i->1	l->1	m->6	r->18	t->1	
ts p	a->1	e->2	l->1	o->4	r->6	u->2	å->18	
ts r	e->15	i->2	ä->6	å->1	
ts s	a->1	e->5	i->5	k->3	l->5	o->7	p->1	t->15	u->2	v->1	y->4	ä->1	å->1	
ts t	a->3	e->1	i->38	j->1	r->3	
ts u	n->9	p->20	t->16	
ts v	a->5	e->3	i->6	ä->2	
ts y	t->3	
ts ä	n->5	r->4	
ts å	l->1	s->1	t->3	
ts ö	n->1	v->3	
ts!F	ö->1	
ts, 	S->1	a->3	b->2	d->2	e->4	f->1	h->1	i->3	m->5	n->4	o->5	p->1	s->4	t->2	u->2	v->5	ä->1	å->2	
ts- 	o->12	
ts-b	e->1	
ts.A	n->1	
ts.B	e->1	
ts.D	e->16	ä->2	å->2	
ts.E	f->1	n->4	r->1	
ts.F	a->1	
ts.H	e->1	o->1	
ts.I	 ->1	
ts.J	a->5	
ts.K	o->3	
ts.M	e->1	i->1	
ts.N	ä->1	
ts.R	a->1	e->1	
ts.S	l->2	o->1	å->1	
ts.T	a->1	
ts.V	i->3	
ts.Ä	n->1	
ts: 	v->1	
ts?F	r->1	
ts?K	o->1	
tsa 	a->1	m->1	p->4	s->1	
tsak	t->5	
tsam	 ->3	,->1	h->6	m->9	t->6	
tsan	a->3	d->5	l->4	
tsar	 ->6	.->1	b->1	g->1	
tsas	 ->4	p->3	
tsat	 ->1	s->59	t->27	
tsav	b->1	t->1	
tsba	n->2	s->2	
tsbe	h->2	k->3	s->6	t->1	
tsbu	d->1	
tsbö	r->5	
tsce	n->1	r->1	
tsch	e->4	
tsde	b->1	
tsdo	k->4	
tse 	d->1	e->2	f->4	m->1	o->2	v->1	
tse.	E->1	
tsed	a->3	d->1	
tsee	n->1	
tsek	t->2	
tsel	 ->4	.->1	
tsen	 ->22	!->1	,->1	.->3	;->1	h->3	
tser	 ->46	,->7	.->8	n->20	
tses	 ->2	.->1	
tset	t->4	
tsfa	t->11	
tsfi	e->1	
tsfl	a->15	
tsfo	r->3	
tsfr	å->10	
tsfå	n->1	
tsfö	r->12	
tsga	r->3	
tsgi	v->8	
tsgr	e->2	u->5	ä->1	
tsha	n->2	
tshj	ä->2	
tsif	f->2	
tsig	a->1	
tsik	t->5	
tsin	s->5	
tsit	u->2	
tska	 ->1	f->1	l->1	m->1	n->1	p->2	
tski	l->3	p->7	
tskl	a->1	i->1	
tsko	e->1	l->1	n->2	t->163	
tskr	a->5	i->4	
tsku	l->1	
tsky	d->8	
tsla	g->20	
tsle	d->28	
tsli	g->134	n->2	v->2	
tslo	g->2	p->2	
tslä	g->3	m->2	n->1	p->9	
tslå	 ->5	r->4	s->8	
tslö	s->43	
tsma	k->2	n->1	r->12	
tsme	d->1	t->3	
tsmi	n->2	
tsmy	n->10	
tsmä	n->2	
tsmå	l->2	
tsni	n->4	v->6	
tsno	r->6	
tsnä	t->1	
tsof	f->2	
tsol	y->1	
tsom	r->6	
tsor	d->13	g->3	
tsos	 ->2	,->1	ä->2	
tspa	k->4	r->1	
tspe	r->2	
tspl	a->11	
tspo	l->7	
tspr	a->1	i->73	o->13	
tspå	r->2	
tsra	m->1	p->2	
tsre	a->1	g->5	
tsri	s->1	
tsru	b->1	m->1	t->1	
tsrä	t->4	
tsrå	d->18	
tssa	n->1	
tsse	k->5	
tssi	f->2	
tssk	i->3	ä->2	
tssp	r->1	
tsst	a->10	y->5	ö->19	
tssy	n->1	s->22	
tssä	k->21	
tsta	g->40	k->1	t->11	
tsti	d->10	l->40	
tstj	ä->1	
tstr	a->3	u->1	ä->30	
tsty	c->3	
tstä	l->53	n->2	
tstå	n->10	r->2	t->1	
tstö	d->2	t->1	
tsug	a->1	
tsut	b->5	s->2	
tsva	g->1	n->1	r->17	
tsve	n->1	r->1	
tsvi	l->5	
tsvä	s->4	
tsyn	p->1	
tsys	t->1	
tsäg	a->2	e->8	
tsäk	e->8	
tsät	t->152	
tså 	E->1	a->5	b->2	d->2	e->4	f->5	g->1	i->11	k->1	l->1	m->2	p->2	r->3	s->11	t->5	v->5	
tså,	 ->2	
tsåg	s->3	
tsåt	g->2	
tt "	P->1	o->1	
tt (	5->1	9->1	
tt -	 ->11	
tt 1	9->3	
tt 2	3->1	5->1	
tt 4	0->1	
tt 5	0->1	
tt 7	0->1	
tt 8	 ->1	0->1	
tt 9	8->1	
tt A	l->1	m->3	
tt B	a->3	e->1	o->1	r->1	
tt C	E->1	
tt D	a->3	
tt E	G->10	I->1	K->1	L->1	U->13	r->1	u->79	v->1	
tt F	E->1	N->2	P->1	l->2	ö->1	
tt G	r->1	
tt H	a->1	
tt I	C->1	N->1	r->1	s->3	t->1	
tt J	ö->3	
tt K	o->2	y->1	
tt M	a->2	
tt N	a->1	
tt O	L->3	
tt P	a->1	o->2	
tt R	I->1	a->1	o->1	
tt S	a->1	o->1	t->1	
tt T	h->2	o->1	u->13	
tt V	ä->1	
tt a	b->1	c->5	d->4	g->14	k->7	l->55	m->3	n->145	r->58	s->1	t->72	v->78	
tt b	a->7	e->217	i->37	l->49	o->8	r->49	u->3	y->16	ä->12	å->4	ö->24	
tt c	e->3	i->2	
tt d	a->9	e->1002	i->59	j->4	o->14	r->25	u->2	y->2	ä->8	å->1	ö->10	
tt e	-->1	f->26	g->14	k->5	l->8	m->1	n->127	p->1	r->20	t->37	u->11	v->3	x->26	
tt f	a->33	e->5	i->19	l->19	o->41	r->79	u->23	y->2	å->90	ö->341	
tt g	a->22	e->135	i->2	l->2	o->26	r->24	y->4	ä->5	å->25	ö->107	
tt h	a->103	e->14	i->11	j->17	o->13	u->12	y->2	ä->12	å->28	ö->19	
tt i	 ->70	.->1	a->1	b->3	c->1	d->6	f->6	g->4	m->3	n->202	r->5	s->2	t->1	
tt j	a->86	o->4	u->7	ä->4	
tt k	a->22	l->20	n->4	o->241	r->32	u->61	v->9	ä->6	ö->4	
tt l	a->48	e->26	i->23	j->1	o->3	u->5	y->15	ä->59	å->14	ö->21	
tt m	a->229	e->77	i->60	o->25	u->3	y->57	ä->11	å->24	ö->12	
tt n	a->6	e->4	i->47	o->6	u->3	y->30	ä->24	å->29	ö->4	
tt o	a->1	b->3	c->53	d->1	e->2	f->10	g->1	k->2	l->7	m->83	n->2	p->4	r->26	s->6	t->1	ä->1	ö->1	
tt p	a->69	e->20	i->1	l->8	o->28	r->69	u->1	å->69	
tt r	a->8	e->92	i->23	o->2	u->2	y->1	ä->21	å->25	ö->33	
tt s	.->1	a->57	e->68	i->17	j->12	k->140	l->24	m->1	n->7	o->58	p->18	t->176	u->3	v->14	y->31	ä->91	å->63	ö->3	
tt t	.->1	a->122	e->4	h->1	i->152	j->3	o->9	r->17	u->3	v->8	y->14	ä->13	å->2	
tt u	l->1	n->75	p->83	r->10	t->164	
tt v	a->76	e->28	i->483	r->1	ä->38	å->22	
tt w	o->1	
tt y	p->1	t->18	
tt z	o->1	
tt ä	g->21	m->2	n->38	r->22	v->20	
tt å	 ->3	k->1	l->1	r->22	s->6	t->50	
tt ö	d->1	g->1	k->22	m->1	n->3	p->9	s->1	v->53	
tt, 	E->1	a->3	b->2	d->2	e->7	f->9	g->3	h->4	i->4	k->4	l->1	m->4	n->1	o->11	p->1	r->1	s->9	t->8	u->2	v->4	ä->3	å->1	
tt. 	D->2	I->1	
tt..	(->1	.->1	
tt.A	l->2	
tt.B	e->1	
tt.D	e->28	ä->2	
tt.E	n->2	r->1	
tt.F	ö->7	
tt.H	e->9	
tt.I	 ->4	
tt.J	a->13	
tt.K	o->3	
tt.L	å->4	
tt.M	a->1	e->7	i->2	o->2	
tt.N	a->1	i->1	ä->1	
tt.O	b->1	m->1	r->1	
tt.P	P->1	a->3	
tt.S	l->1	o->1	t->1	y->1	
tt.T	a->1	
tt.U	t->1	
tt.V	i->7	
tt.Ä	v->3	
tt: 	"->2	H->1	j->1	o->1	s->1	
tt?A	n->1	
tt?D	e->1	
tt?O	m->1	
tt?S	k->1	
tt?V	i->1	
ttBe	t->1	
tta 	-->6	A->1	E->8	F->1	a->55	b->77	c->2	d->75	e->55	f->93	g->14	h->32	i->58	k->39	l->15	m->76	n->14	o->76	p->99	r->14	s->145	t->26	u->26	v->34	y->2	ä->160	å->9	ö->6	
tta!	D->1	F->1	
tta,	 ->47	
tta.	 ->1	(->1	.->1	A->1	B->2	C->1	D->20	E->5	F->2	G->1	H->3	I->6	J->8	K->1	M->6	N->2	O->3	P->3	S->5	T->1	V->11	Ä->1	
tta:	 ->1	
tta?	J->1	
ttac	k->3	
ttad	 ->2	e->22	
ttag	.->1	a->11	e->1	i->3	n->2	
ttal	a->98	
ttan	 ->2	.->1	d->66	t->1	
ttar	 ->62	.->1	e->18	h->1	n->5	
ttas	 ->51	,->4	.->4	
ttat	 ->20	.->1	s->14	
ttav	l->7	
tte 	O->1	d->2	i->2	j->1	m->1	o->2	p->10	r->6	ö->2	
tte,	 ->1	
tte-	 ->1	L->1	
tteb	a->1	e->14	
tted	e->1	
ttef	r->2	ö->1	
tteg	å->1	
ttei	n->2	
ttel	i->1	s->3	ä->1	
tten	 ->124	!->2	)->1	,->27	.->37	;->2	?->1	F->1	H->1	d->2	f->2	l->1	p->1	r->2	s->10	t->5	v->8	
ttep	o->1	
tter	 ->88	,->3	.->2	a->35	d->3	i->8	l->55	n->4	o->1	r->2	s->34	v->1	
ttes	 ->6	.->2	a->1	y->1	
ttet	 ->135	,->9	.->11	:->1	s->7	
ttfr	a->1	
ttfu	l->1	
ttfä	r->7	
ttfö	r->1	
ttgö	r->1	
tthå	l->9	
tti 	g->1	
ttic	h->1	
ttid	e->1	
ttig	 ->7	a->43	d->12	h->103	t->4	
ttil	l->47	
ttin	,->1	n->1	
ttio	f->1	t->1	
ttis	k->16	
ttit	 ->1	y->5	
ttja	 ->18	d->4	n->9	r->3	s->6	t->1	
ttjä	n->25	
ttkr	i->1	
ttkv	ä->1	
ttla	n->5	
ttle	 ->3	.->1	
ttli	g->2	
ttmä	t->1	
ttmå	l->1	
ttna	 ->3	.->1	d->1	r->7	s->3	
ttne	 ->2	n->3	t->6	
ttni	n->287	
tto 	a->1	f->1	
tto-	a->1	
ttoa	n->1	
ttol	k->1	
tton	 ->4	a->1	d->2	e->1	s->1	
ttor	 ->1	k->1	n->1	
ttra	 ->47	d->6	f->1	k->1	n->33	r->6	s->7	t->4	
ttre	 ->69	,->3	.->6	t->1	
ttri	n->21	
ttry	c->72	
tträ	d->5	
tts 	a->8	b->1	f->9	g->1	h->1	i->4	k->1	m->2	n->1	o->1	p->1	u->5	v->1	ö->1	
tts,	 ->3	
tts-	 ->1	
tts.	D->3	E->1	I->1	N->1	R->1	
ttsa	k->4	
ttsb	e->6	
ttsd	e->1	
ttsf	r->1	ö->1	
ttsh	j->2	
ttsi	n->2	
ttsk	a->1	i->7	u->1	
ttsl	i->132	ä->3	
ttsm	y->1	å->1	
ttso	f->2	m->1	r->3	s->2	
ttsp	a->1	r->3	
ttsr	e->2	u->1	
ttss	e->1	k->3	t->9	y->20	ä->20	
ttst	i->2	j->1	r->1	
ttsv	ä->4	
ttvi	k->2	l->1	s->72	
ttys	k->2	
ttän	k->1	
tté 	-->2	e->1	f->3	h->1	m->1	s->2	
ttée	r->4	
ttéf	ö->2	
ttén	 ->23	,->4	.->2	?->1	s->11	
ttés	y->2	
ttöm	d->1	m->3	t->1	
tu m	e->21	
tual	i->1	
tuat	i->129	
tud 	7->1	
tude	n->2	r->3	
tudi	e->9	
tuel	l->55	
tuer	a->3	
tuff	 ->1	a->1	
tuga	l->26	
tugi	s->70	
tugo	r->1	
tugu	e->1	
tula	t->6	
tule	r->33	
tull	a->2	f->1	g->1	
tum 	a->56	d->1	f->3	i->1	m->1	o->3	s->5	ä->4	å->1	
tum,	 ->3	
tum.	D->1	I->1	V->2	
tume	t->3	
tumm	a->3	
tunc	 ->1	
tund	 ->8	a->2	e->7	
tung	 ->6	a->3	m->6	r->1	t->2	
tuni	s->2	
tunn	e->3	l->2	
tur 	-->2	2->20	b->3	d->3	e->1	f->7	g->1	h->1	i->4	k->1	o->7	p->1	s->8	u->2	v->2	ä->4	
tur,	 ->19	
tur-	 ->2	
tur.	D->3	F->1	N->1	O->1	T->1	V->3	
tur?	M->1	
tura	.->1	k->1	n->1	r->6	
turb	e->1	
ture	l->40	n->54	r->42	
turf	o->59	ö->2	
turh	i->1	
turi	e->1	s->24	
turk	-->1	a->15	i->6	
turl	i->102	
turm	ä->1	
turn	ä->1	ö->1	
turo	m->2	
turp	o->16	r->4	
turr	e->1	
turs	e->5	t->3	
turu	t->3	
turv	e->1	
turå	t->1	
tus 	a->1	e->1	q->2	
tus.	D->1	
tus?	O->1	
tuse	n->17	
tusf	ö->1	
tusi	a->3	
tuti	o->158	
tuts	k->12	
tutv	i->2	
tvak	t->1	
tval	d->1	
tvap	e->1	
tvar	a->2	o->1	
tvec	k->238	
tvek	a->23	l->1	s->5	
tver	k->29	s->1	
tvet	y->7	
tvid	g->107	
tvik	t->6	
tvil	l->2	
tvin	 ->1	g->32	
tvis	 ->132	,->6	.->4	a->51	o->3	t->19	
tviv	e->33	l->10	
tvun	g->11	
tvän	l->1	
tvär	d->33	l->1	p->2	s->1	t->14	
tvät	t->5	
två 	a->10	b->3	d->2	e->7	f->23	g->2	h->2	i->3	j->1	k->4	l->2	m->8	n->2	o->2	p->12	r->2	s->12	t->8	u->3	v->5	y->1	å->8	
två.	B->1	
två:	 ->2	
tvåh	u->1	
tvån	g->6	
ty E	u->1	
ty d	e->4	
ty i	 ->1	
ty n	a->1	ä->1	
ty p	å->2	
ty v	i->2	
ty ä	r->1	
ty-p	r->1	
tyck	a->3	e->71	l->5	s->8	t->7	
tyd 	g->1	i->1	s->1	t->1	
tyd.	S->1	
tyda	 ->1	n->16	
tydd	e->3	
tyde	l->73	r->24	
tydi	g->11	
tydl	i->124	
tyg 	d->1	f->5	i->4	m->3	n->1	o->3	s->15	u->3	
tyg)	,->1	
tyg,	 ->3	
tyg.	E->1	F->1	V->2	
tyg;	 ->1	
tyg?	D->1	
tyga	 ->10	d->21	n->5	r->1	
tyge	l->5	n->13	t->7	
tygs	b->1	i->1	s->9	t->1	ä->1	
tymp	a->1	n->2	
tyna	n->1	
tyng	a->1	d->6	e->1	s->2	
typ 	C->1	a->18	f->1	
typ,	 ->2	
typ.	D->1	E->1	
type	n->12	r->4	
typf	a->1	
typg	o->1	
tyr 	a->1	
tyr.	E->1	
tyra	 ->9	n->4	r->5	s->2	
tyre	 ->1	,->1	k->3	l->7	n->1	t->3	
tyrk	a->13	e->2	o->2	
tyrn	i->7	
tyrs	 ->2	
tysk	a->21	l->2	t->2	
tyst	 ->3	
tyvä	r->30	
tz i	 ->1	
tz o	c->1	
tz s	o->1	
tz, 	p->1	
tz. 	E->1	
tzid	a->2	
täck	a->9	e->10	n->1	s->6	t->5	
täda	 ->1	t->1	
täde	r->17	s->2	
täkt	s->5	
täll	a->136	b->1	d->67	e->104	i->6	n->70	s->20	t->22	
tämd	 ->5	a->8	e->5	h->1	
täml	i->3	
tämm	a->24	e->159	i->4	
tämn	i->2	
tämp	e->1	l->1	
täms	 ->1	
tämt	 ->13	,->3	
tän 	e->1	
tänd	a->6	i->107	l->1	
täng	a->2	d->1	e->1	n->6	t->1	
tänk	 ->1	a->318	b->3	e->36	l->5	s->2	t->12	
täpp	a->3	e->1	
tär 	a->2	f->1	o->2	v->1	
tär,	 ->1	
tär.	R->1	
tära	 ->11	
täre	n->2	r->2	
tärk	a->28	e->3	n->6	s->5	t->9	
tärt	 ->2	
täta	,->1	r->1	
täte	n->2	
täth	e->1	
täv 	m->1	
tävj	a->1	
tävl	a->2	i->1	
tå a	l->1	t->11	v->4	
tå d	e->3	
tå e	n->1	
tå f	o->1	r->8	ö->12	
tå h	u->2	
tå i	 ->4	n->1	
tå k	l->3	v->1	
tå n	y->1	ä->1	
tå o	c->2	m->1	
tå s	o->1	
tå t	i->1	
tå u	t->2	
tå v	a->4	
tå, 	a->1	f->1	s->1	
tå.F	P->1	
tå.J	u->1	
tå: 	å->1	
tådd	 ->1	a->1	
tåel	i->6	s->8	
tåen	d->32	
tåg 	e->1	
tåg,	 ->1	
tåge	t->1	
tågk	r->1	
tågo	l->1	
tål 	a->1	
tåla	m->2	
tålf	ö->5	
tålg	e->1	
tåli	g->2	n->25	
tåls	e->5	t->1	
tålv	e->5	
tånd	 ->54	,->8	.->10	?->2	a->5	e->30	i->1	p->97	s->19	
tår 	a->25	d->13	e->6	f->20	g->1	h->9	i->44	j->3	k->10	l->2	m->7	n->2	o->2	p->14	s->2	t->4	u->1	v->8	ä->1	å->1	ö->2	
tår,	 ->3	
tår.	D->2	H->1	
tåre	t->10	
tås 	d->1	f->1	k->1	s->1	u->1	v->1	
tåt"	,->1	
tåtg	ä->3	
tått	 ->27	,->1	.->1	s->1	
té -	 ->2	
té e	l->1	
té f	ö->3	
té h	a->1	
té m	e->1	
té s	o->2	
téer	.->1	n->3	
téfö	r->2	
tén 	(->2	f->3	i->1	k->1	l->1	o->11	s->2	v->1	ä->1	
tén,	 ->4	
tén.	H->1	M->1	
tén?	V->1	
téns	 ->11	
tésy	s->2	
tête	 ->3	
tóni	o->1	
töd 	-->2	a->5	b->1	d->3	e->3	f->26	g->1	h->2	i->11	k->5	l->1	m->5	o->16	p->7	s->20	t->43	v->4	ä->2	å->2	ö->1	
töd,	 ->14	
töd.	"->1	.->1	A->1	D->10	E->1	F->2	H->5	I->2	J->2	M->1	N->1	O->1	R->1	S->1	T->1	U->1	V->2	Ä->2	Å->2	
töd;	 ->1	
töd?	-->1	
tödd	e->2	
töde	n->32	r->58	t->32	
tödj	a->71	e->1	
tödm	e->1	o->1	
tödn	i->1	
tödp	o->1	
tödr	a->2	
töds	 ->8	p->1	y->4	
tödå	t->5	
töka	 ->6	d->1	n->1	s->2	t->1	
tökn	i->1	
töld	,->1	
tömd	,->1	
tömm	a->3	e->1	
tömt	 ->1	
tör 	b->1	i->1	k->1	m->1	s->1	
tör,	 ->1	
töra	 ->2	s->3	
törd	a->1	e->2	
töre	l->5	n->3	r->23	
töri	n->2	
törn	i->5	
törr	e->75	
törs	 ->1	,->1	k->1	o->1	t->37	
tört	n->1	s->2	
töta	 ->1	n->1	r->1	
töte	r->1	s->1	
tötf	å->1	
tött	 ->10	a->2	s->1	
töva	 ->7	n->1	r->3	s->4	
töve	r->21	
tövn	i->1	
türk	d->1	
u - 	a->1	
u 34	 ->1	
u Ah	e->2	
u An	g->1	
u Be	r->1	
u Eg	y->1	
u Er	i->1	
u Fr	a->1	
u Ly	n->1	
u Mc	N->1	
u Mo	r->1	
u Pe	i->1	
u Pl	o->1	
u Re	d->3	
u Sc	h->3	
u Su	d->1	
u Th	e->1	
u Wa	l->1	
u ab	s->1	
u al	l->6	
u an	g->1	m->1	s->1	v->1	
u at	t->8	
u av	 ->2	
u ba	i->1	r->2	
u be	f->1	h->3	r->1	t->1	
u bl	i->3	o->1	
u co	m->1	
u de	 ->1	f->1	s->1	t->3	
u di	r->1	s->2	
u du	 ->1	
u dä	r->1	
u då	 ->1	
u dö	p->1	
u ef	t->1	
u eg	e->1	
u em	e->1	
u en	 ->13	
u et	t->8	
u eu	r->1	
u fa	k->1	t->1	
u fi	n->4	
u fl	e->1	
u fr	a->1	å->2	
u få	r->2	t->2	
u fö	g->1	r->16	
u ge	m->1	n->1	r->2	t->1	
u gä	l->3	
u gå	 ->3	n->1	
u gö	r->3	
u ha	r->19	
u ho	t->1	
u hä	r->1	
u hå	l->1	r->2	
u hö	g->4	r->1	
u i 	T->1	p->1	s->1	v->1	
u ig	e->1	
u in	b->1	d->1	g->2	l->1	n->3	o->1	s->1	t->40	
u is	o->1	
u ka	n->7	
u ko	m->51	n->1	
u le	d->2	
u li	g->1	
u ly	s->1	
u lä	g->1	n->1	s->1	t->1	
u me	d->23	n->1	r->11	
u mi	g->1	n->2	
u mo	r->1	
u mä	r->1	
u må	s->10	
u nu	m->1	
u nä	r->8	
u nå	t->1	
u oc	h->6	k->8	
u of	f->1	t->2	
u om	s->1	
u pa	r->1	
u pl	a->1	
u po	r->1	
u pr	i->1	ö->1	
u pu	n->1	
u på	 ->2	.->1	g->2	
u re	d->2	s->1	
u ru	l->1	
u rå	d->2	
u rö	s->1	
u sa	 ->1	d->2	m->3	
u se	r->1	s->1	
u si	f->1	n->1	
u sk	a->4	e->1	u->1	ö->1	
u sl	å->1	
u sm	i->1	
u so	m->2	
u sp	e->1	
u st	a->1	r->1	ä->3	å->3	ö->6	
u sv	å->1	
u sä	g->1	t->1	
u så	 ->2	
u ta	g->2	l->84	r->2	
u ti	l->5	
u ty	d->2	v->1	
u un	d->1	
u up	p->3	
u ut	t->1	
u va	d->1	
u ve	m->1	r->2	
u vi	d->2	k->2	l->2	s->1	
u vä	n->1	
u äl	d->1	
u än	 ->1	d->2	t->5	
u är	 ->23	,->1	
u åt	e->2	
u", 	d->1	
u, L	a->1	
u, a	n->1	
u, e	f->2	n->1	
u, h	a->1	
u, i	 ->1	
u, m	e->2	
u, o	c->2	
u, p	r->1	
u, s	i->1	o->2	
u, u	n->1	
u, å	t->1	
u, ö	v->1	
u-lä	n->1	
u..T	a->1	
u.De	t->1	
u.Et	t->1	
u.Ja	g->1	
u.Ko	m->1	n->1	
u.Lå	t->1	
u.Vi	 ->2	
u: g	ö->1	
u; i	 ->1	
u?Ja	g->1	
uMed	 ->1	
ua n	o->2	
uade	s->1	
ual 	D->1	h->1	s->2	v->1	ä->1	
ual"	 ->1	
ual,	 ->1	
uali	s->2	t->1	
uanz	e->1	
uari	 ->19	!->1	,->10	.->2	
uate	m->1	
uati	o->129	
ubba	 ->1	r->1	s->1	
ubbe	l->6	
ubbl	a->11	
ubet	ä->1	
ubik	m->2	
ubje	k->1	
ubla	n->1	
ubli	c->6	k->20	n->7	
ubri	k->2	
ubsi	d->23	
ubst	a->4	
ubve	n->12	
uc s	e->1	
ucce	s->5	
ucen	t->22	
ucer	a->12	i->1	
uchn	e->12	
ucka	 ->1	"->1	,->1	
ucki	t->1	
uckn	e->1	
ucko	r->2	
ucto	r->1	
ud 7	 ->1	
ud B	a->2	
ud e	l->1	
ud f	a->1	ö->4	
ud m	e->2	o->7	
ud o	c->4	
ud r	e->1	
ud t	a->9	
ud v	i->1	
ud ä	r->1	
ud, 	a->1	e->1	h->1	s->1	
ud.D	e->2	
ud.V	a->1	
uda 	a->1	b->3	d->1	e->3	i->1	k->1	m->1	n->1	o->1	p->1	u->1	
udak	t->2	
udan	 ->1	d->4	g->1	s->4	
udap	e->1	
udar	s->1	
udas	,->1	.->1	
udda	 ->2	
udde	l->3	
uddh	i->1	
uddi	g->2	
ude 	M->1	
uden	 ->1	t->2	
uder	 ->11	,->1	a->7	
udet	 ->11	,->1	.->1	?->1	
udeu	t->1	
udfr	å->4	
udfö	r->1	
udge	t->107	
udic	e->1	
udie	 ->1	b->1	p->1	r->6	
udik	a->3	
udis	k->1	
udit	 ->1	
udli	g->1	n->2	
udmå	l->2	
udna	 ->2	
udni	n->1	
udor	d->1	
udre	 ->1	,->1	k->1	
udro	l->2	n->1	
uds 	s->2	
udsa	k->16	
udsf	ö->3	
udsi	n->3	
udsk	a->10	
udsm	a->10	
udsp	r->1	
udst	a->2	ä->2	
udsy	f->1	
udup	p->1	
ue k	a->1	
ue, 	s->1	v->1	
uece	d->1	
ueir	a->1	
uela	 ->1	
uell	 ->9	.->4	a->38	t->16	
uen,	 ->1	
uer 	h->1	s->1	t->1	
uer,	 ->1	
uera	 ->5	d->1	r->1	t->1	
uerl	i->2	
uern	t->1	
ues 	D->3	e->1	
ues"	.->1	
uesa	 ->1	
uff 	n->1	
uffa	r->1	
ufma	n->1	
uft 	g->1	
uft.	V->1	
uftb	u->1	
ufte	t->1	
ufti	g->11	
ufto	m->1	
uför	a->1	
uga,	 ->1	
ugal	 ->15	,->4	s->7	
ugar	e->1	
ugen	 ->1	.->1	
uger	 ->1	
ugg 	p->3	
ugga	 ->1	n->1	
uggb	o->1	
ugge	n->1	
uggl	i->1	
ugis	i->70	
ugli	g->6	
ugn 	o->1	
ugna	 ->2	d->1	n->1	s->1	
ugo 	g->1	å->1	
ugof	e->1	
ugon	d->1	
ugor	,->1	
ugos	l->1	
ugue	s->1	
uham	e->1	
uhe 	o->1	
uhe,	 ->1	
uhne	,->1	
uier	d->1	
uigo	u->1	
uine	r->1	
uins	 ->1	
uiol	a->1	
uise	n->3	
uisi	t->1	
uita	 ->1	
uiz 	s->1	
uk a	l->1	v->1	
uk m	e->1	
uk o	c->5	
uk p	å->1	
uk s	o->1	
uk!A	n->1	
uk, 	d->3	e->1	i->1	m->1	t->2	v->1	
uk.J	a->1	
uka 	P->1	
uka,	 ->1	
ukad	e->2	
ukar	 ->3	:->1	e->8	n->5	
ukas	 ->1	.->1	u->3	
ukdo	m->1	
uken	.->1	
uket	 ->13	,->2	.->1	;->2	s->1	
ukfö	r->1	
ukhu	s->7	
ukit	s->1	
ukni	n->3	
ukse	k->1	
uksf	o->1	r->1	
uksl	o->1	
ukso	m->2	
uksp	o->6	r->3	
uksr	e->2	
ukss	e->5	y->1	
ukt 	a->2	h->1	p->1	s->3	
ukt,	 ->1	
ukt.	H->1	
ukta	n->7	r->4	t->1	
uktb	a->2	
ukte	n->7	r->10	
ukti	g->1	n->1	o->39	v->21	
ukto	r->6	
ukts	 ->2	
uktu	r->153	
uktö	r->3	
ukvå	r->3	
ul f	ö->1	
ul o	c->1	m->1	
ul s	o->1	
ul.V	i->1	
ula 	o->1	ö->1	
ula.	J->1	
ulad	a->1	
ulan	s->5	
ular	i->1	y->1	
ulat	i->12	o->2	
ulda	 ->1	n->1	
uldb	e->1	
ulde	n->2	r->1	
ulen	 ->1	
uler	 ->3	a->55	i->6	
ulf-	M->2	
ulfe	r->1	
ulfk	r->1	
ulga	r->1	
uli 	1->4	2->2	f->1	u->1	
uli,	 ->2	
ulis	m->1	s->1	t->3	
ulkl	a->1	
ull 	a->2	b->3	e->1	f->2	g->4	h->3	i->2	n->1	o->1	p->1	r->2	s->3	v->1	ä->1	ö->1	
ull,	 ->3	
ull.	D->3	K->1	O->1	V->1	
ulla	 ->19	,->1	.->2	r->6	s->1	
ullb	o->3	
ulle	 ->484	,->2	
ullf	ö->4	
ullg	j->1	å->1	ö->1	
ullh	e->1	
ulli	t->1	
ullk	a->1	o->5	
ullo	 ->5	
ulls	t->44	
ullt	 ->40	,->1	.->2	
ullv	ä->2	
ullä	n->2	
ulor	 ->1	
ulos	 ->5	
uls 	f->1	t->1	
ulse	r->4	
ulsk	a->1	
ult 	d->1	k->1	
ulta	t->111	
ultb	a->1	
ulte	n->20	r->9	
ulth	e->6	
ulti	e->3	l->1	m->1	n->5	
ultr	a->2	
ultu	r->146	
ulz 	e->1	s->2	
uläg	e->1	
ulär	a->2	t->1	
um -	 ->1	
um a	t->56	v->3	
um b	l->1	
um d	å->1	
um e	g->1	n->1	
um f	i->1	r->1	ö->9	
um h	a->2	ä->1	
um i	 ->17	n->5	
um m	e->2	i->1	å->1	
um o	c->9	m->3	
um p	å->4	
um s	k->2	o->6	
um u	n->1	t->1	
um v	ä->1	
um y	t->1	
um ä	n->1	r->4	
um å	s->1	t->1	
um!D	e->1	
um!M	e->1	
um, 	b->1	d->2	k->2	m->1	o->3	p->1	u->1	v->1	
um. 	D->1	
um.A	t->1	v->1	
um.D	e->4	
um.H	e->1	
um.I	 ->1	
um.L	å->1	
um.M	e->1	
um.O	M->1	
um.P	r->1	
um.R	å->1	
um.S	o->1	
um.V	i->2	
um.Ä	n->1	
uman	 ->1	i->5	
umar	 ->1	
umat	i->1	
umba	r->1	
umbä	r->4	
umen	t->176	
umer	a->6	
umet	 ->5	.->1	
umgä	n->1	
umhe	t->3	
umle	n->1	
umma	 ->5	d->1	n->2	t->1	
umme	l->6	r->2	
ummi	p->1	
ummo	r->8	
ump 	a->2	s->1	
ump.	D->1	
umpa	n->1	s->2	
umpe	r->2	
umpn	i->3	
umra	 ->1	
umt 	a->1	
umta	n->1	
umti	o->2	
umul	a->1	e->1	
umän	i->1	
umör	 ->2	
un s	a->1	
un.D	e->1	
una 	p->1	ä->1	
unal	a->2	p->1	
unan	s->1	
unc 	d->1	
unch	t->1	
unci	l->1	
und 	(->2	L->1	a->81	e->1	f->17	i->3	o->1	s->7	t->1	u->1	v->2	ä->2	
und,	 ->2	
und.	D->1	N->1	P->1	
und?	 ->1	
unda	 ->19	,->1	.->2	d->8	m->1	n->58	r->4	s->6	t->5	
undb	u->1	
unde	 ->31	n->42	r->498	t->14	
undf	ö->4	
undg	ä->2	å->1	
undi	 ->2	:->1	t->3	
undk	u->1	
undl	i->16	ä->74	
undn	a->4	
undo	r->1	
undp	e->1	r->1	
undr	a->33	e->2	i->1	
unds	a->1	j->1	k->1	l->2	r->5	t->1	
undt	e->1	
undv	a->26	i->39	
undä	r->1	
uner	 ->7	a->1	n->2	s->1	
ung 	a->1	b->1	m->1	o->3	p->2	u->1	
ung.	 ->1	I->1	O->1	
unga	 ->6	,->2	n->1	r->15	
ungd	o->14	
unge	f->8	l->2	n->5	r->54	t->2	
ungf	r->1	
ungl	i->13	
ungm	e->6	
ungn	a->6	
ungr	o->1	
ungs	l->1	
ungt	 ->1	,->1	
unha	s->1	
uni 	1->6	2->2	f->2	i->1	v->1	
unic	e->2	
unik	a->17	t->1	
unil	a->2	
unio	n->437	
unis	m->2	t->1	
unit	e->1	
univ	e->4	
unka	 ->3	.->1	
unke	r->3	
unki	t->2	
unkl	a->1	
unkn	a->4	
unkt	 ->133	,->14	.->19	:->2	?->1	e->173	i->32	s->2	u->1	
unna	 ->211	.->1	n->2	r->2	t->43	
unne	l->3	n->2	t->1	
unni	g->6	t->16	
unnl	a->2	
unno	r->1	
uno 	L->1	
unsk	a->17	
unt 	o->3	t->1	
unt.	D->1	
unta	 ->2	r->5	
untl	i->8	
unto	m->1	r->1	
untp	r->1	
untr	a->21	
uo s	o->1	
uo, 	d->1	
up ,	 ->1	
up d	e->1	
up ö	n->1	
upa 	f->1	m->1	o->1	s->1	u->1	
upa,	 ->1	
upad	 ->1	
upan	t->1	
upar	e->1	
upas	 ->1	t->2	
upat	 ->2	i->1	
uper	a->3	
upet	 ->3	,->2	
upgå	e->7	
upni	n->5	
upp 	(->2	-->1	E->1	T->1	a->20	b->4	d->41	e->21	f->17	g->3	h->9	i->24	k->6	l->5	m->9	n->5	o->9	p->12	r->6	s->16	t->16	u->8	v->7	ä->9	
upp,	 ->20	
upp.	A->1	D->4	F->1	J->7	M->1	P->1	V->2	Ä->2	
upp?	H->1	
uppb	a->1	r->3	y->20	ä->1	å->1	
uppd	a->2	e->3	r->22	
uppe	h->13	n->98	r->57	
uppf	a->52	y->54	ö->23	
uppg	i->77	r->1	å->8	ö->2	
upph	e->1	o->13	ä->5	ö->10	
uppk	o->7	
uppl	e->17	i->1	y->4	ö->3	
uppm	a->58	j->2	u->21	ä->55	
uppn	å->93	
uppo	r->1	
uppr	e->54	i->6	o->5	u->1	y->1	ä->38	ö->5	
upps	 ->4	a->7	k->29	p->2	t->39	ä->3	
uppt	a->10	i->1	o->2	r->10	ä->11	
uppu	n->1	
uppv	i->6	ä->2	
upra	n->1	
upsi	n->1	
upsk	h->1	
upt 	b->2	d->1	o->1	s->1	v->1	ö->1	
upti	o->7	
upér	y->1	
uqal	 ->2	
ur -	 ->2	
ur 2	0->20	
ur E	G->1	U->1	u->2	
ur U	C->1	
ur a	l->1	n->2	r->1	v->1	
ur b	a->1	e->5	i->2	r->4	u->2	y->1	
ur d	e->46	i->1	r->1	ä->1	
ur e	k->2	n->8	r->1	t->5	
ur f	a->1	o->2	r->1	ö->11	
ur g	e->1	o->1	å->1	ö->1	
ur h	a->3	o->2	ö->1	
ur i	 ->2	n->4	
ur j	o->1	
ur k	a->2	l->3	o->10	u->1	ä->1	
ur l	e->1	i->2	ä->3	å->5	
ur m	a->19	e->1	i->6	y->2	ä->1	å->7	
ur n	i->3	u->2	
ur o	c->9	f->1	
ur p	a->3	e->2	o->1	r->2	å->1	
ur r	i->1	
ur s	a->1	e->3	i->1	k->11	m->1	n->1	o->19	t->12	v->5	ä->1	ö->1	
ur t	e->1	i->1	r->1	u->1	ä->1	
ur u	n->3	p->1	r->1	t->4	
ur v	e->1	i->30	ä->2	å->1	
ur ä	r->6	
ur, 	(->1	G->1	a->3	f->1	h->1	l->1	m->3	o->3	s->1	t->2	u->3	å->1	
ur- 	o->4	
ur.D	e->3	ä->1	
ur.F	o->1	
ur.H	e->1	
ur.K	o->1	
ur.N	i->1	
ur.O	m->1	
ur.R	å->1	
ur.T	y->1	
ur.V	i->3	
ur?M	e->1	
ura 	f->3	o->1	s->2	
ura,	 ->2	
ura.	D->1	
urak	t->1	
ural	i->1	
uran	 ->3	.->1	?->1	i->2	s->1	v->4	
urar	 ->1	b->1	n->1	t->1	v->5	
uras	 ->1	
urat	 ->1	o->4	
urba	n->1	
urbe	s->1	
urd 	i->1	
urel	l->40	
uren	 ->37	,->5	.->4	?->1	s->8	
urer	 ->12	,->4	.->4	a->6	i->10	n->6	s->1	
ures	 ->1	
uret	 ->2	
urfo	d->4	n->58	r->1	
urfö	r->2	
urg 	f->1	i->1	m->2	u->1	ö->1	
urg,	 ->4	
urg.	D->1	J->1	L->1	V->1	
urga	r->1	
urgh	.->1	
urhi	s->1	
urho	l->4	
uri.	B->1	
urid	i->30	
urie	-->1	n->1	
uris	 ->4	.->1	d->5	m->20	t->11	
urit	 ->1	a->1	
urk-	d->1	
urka	r->2	t->13	
urki	e->35	s->6	
urkm	e->2	
urla	n->6	
urli	g->102	v->2	
urmi	n->1	
urmä	s->1	
urna	.->1	l->2	
urne	r->1	
urnä	t->1	
urnö	d->1	
uro 	1->1	b->1	f->6	h->1	i->1	o->1	p->3	t->1	u->1	
uro!	A->1	
uro,	 ->8	
uro-	r->1	
uro.	D->3	H->1	K->1	N->1	S->1	V->1	
urod	a->5	
urof	e->1	
uroj	u->6	
urom	r->2	
uron	 ->3	,->1	s->3	
uroo	m->1	
urop	a->468	e->712	o->16	r->1	é->10	
uros	k->3	t->1	
urpo	l->16	
urpr	o->4	
urre	f->1	g->1	n->280	r->5	
urs 	d->1	i->1	m->2	o->1	
urs,	 ->1	
urs.	D->1	
ursb	r->1	
urse	k->5	n->4	r->52	
ursf	ö->1	
ursk	i->3	u->1	
ursp	r->19	å->1	
urss	l->1	
urst	i->1	ö->3	
ursä	k->14	n->1	
urt 	a->1	m->1	
urtz	 ->2	,->1	
urut	g->1	s->1	v->1	
uruv	i->15	
urva	l->5	t->8	
urve	t->1	
urvi	s->1	
uråt	g->1	
us 1	9->1	
us 2	0->1	
us a	n->1	v->1	
us b	e->3	
us e	n->2	
us f	y->1	ö->1	
us h	a->1	
us j	u->5	
us k	a->1	r->1	
us o	c->3	
us p	å->1	
us q	u->2	
us s	o->1	t->1	
us t	j->1	r->1	
us u	n->1	
us ä	r->1	
us, 	e->1	f->1	h->1	m->2	
us-b	e->1	
us.D	e->2	
us.E	u->1	
us.G	e->1	
us.H	e->1	
us.I	n->1	
us?O	c->1	
usa 	v->1	
usal	e->2	
usar	 ->2	
usch	w->1	
usdi	m->1	
use"	,->1	
usef	f->3	
usen	 ->5	,->1	d->3	t->10	
user	a->3	
uset	 ->10	.->1	
usew	i->1	
usfö	r->1	
usga	s->4	
usgr	a->2	
ush 	P->1	
ush,	 ->1	
ushå	l->1	
usia	s->3	
usik	 ->2	e->2	
usio	n->8	
usiv	 ->1	a->1	e->17	t->1	
usk.	H->1	
usko	u->1	
uslä	k->1	
usp"	,->1	
uspe	n->1	
usqu	i->1	
ussa	 ->1	g->1	r->2	s->1	
usse	l->2	n->1	
ussi	n->1	o->61	
ussl	a->2	
ust 	a->3	b->3	d->18	e->2	f->12	g->3	h->15	i->6	l->2	m->3	n->14	o->1	p->6	r->1	s->8	v->3	ö->1	
ust,	 ->1	
ust.	D->1	K->1	V->1	
ust:	 ->1	
usta	 ->1	a->1	d->2	
ustb	e->2	r->1	
uste	n->18	r->21	
usti	c->4	t->6	
ustl	i->2	
ustm	y->3	
ustn	i->5	
usto	m->2	
ustr	a->1	e->2	i->114	
ustv	a->1	
usul	 ->2	.->1	e->3	
usí 	ä->1	
usöv	e->1	
ut -	 ->1	
ut 1	0->1	
ut 8	8->2	
ut 9	4->1	
ut T	o->1	
ut a	c->1	m->1	n->2	t->8	v->3	
ut b	e->4	o->1	ö->2	
ut d	e->7	i->1	
ut e	n->5	t->2	x->1	
ut f	a->1	o->1	r->9	ö->9	
ut g	e->1	o->1	
ut h	a->6	ö->1	
ut i	 ->10	n->10	
ut k	a->2	o->2	u->1	
ut l	a->1	y->1	ä->1	å->1	
ut m	e->4	i->2	o->2	y->2	ö->1	
ut n	a->1	r->1	ä->1	å->1	ö->10	
ut o	c->11	m->20	s->1	
ut p	e->2	l->1	o->1	r->2	å->24	
ut r	e->3	
ut s	e->1	i->2	k->1	o->14	t->2	y->1	ä->1	å->2	
ut t	a->1	i->4	
ut u	n->2	p->1	t->3	
ut v	a->1	i->2	
ut ä	n->1	r->3	
ut å	s->1	
ut ö	v->5	
ut, 	a->4	b->1	e->1	f->2	h->4	i->2	m->4	n->1	o->5	s->4	t->2	u->2	v->1	å->1	
ut. 	D->2	
ut.(	P->1	
ut.)	F->1	
ut.D	e->7	å->2	
ut.F	i->1	r->1	ö->2	
ut.G	r->1	
ut.I	n->1	
ut.J	a->5	
ut.K	r->1	
ut.N	a->2	
ut.O	c->1	
ut.S	k->1	t->1	
ut.T	v->1	
ut.V	a->1	i->1	
ut.Ä	v->1	
ut: 	f->1	
ut; 	d->1	
ut?.	 ->1	
ut?E	t->1	
uta 	a->2	d->4	e->2	f->2	g->2	i->2	k->1	l->1	m->7	o->12	p->1	r->2	s->7	u->6	v->2	Ö->2	
uta,	 ->5	
utab	e->2	l->1	
utad	,->1	.->18	e->11	
utaf	r->10	
utal	.->1	a->1	
utan	 ->292	,->4	.->1	d->27	f->32	v->1	
utap	o->1	
utar	 ->8	.->1	b->31	m->10	
utas	 ->11	p->2	
utat	 ->11	s->3	
utau	n->3	
utba	s->1	
utbe	s->1	t->7	
utbi	l->60	
utbr	e->4	
utbu	d->4	
utby	g->3	t->17	
utde	l->1	
ute 	e->1	p->1	t->1	u->1	
utea	u->3	
utel	ä->3	
uten	 ->15	,->2	.->3	s->1	
uter	 ->17	,->1	.->6	a->78	r->2	
utes	l->19	t->4	
utet	 ->52	,->2	.->1	?->1	s->1	
utfa	l->1	s->3	
utfl	a->1	y->1	
utfo	r->40	
utfr	å->7	
utfä	r->12	s->1	
utfö	r->46	
utga	v->1	
utgi	c->1	f->14	l->8	v->2	
utgj	o->4	
utgå	 ->4	n->16	r->8	v->1	
utgö	r->59	
utha	n->1	
uthe	r->1	
uthä	r->4	
utie	r->1	
utif	r->16	
utik	 ->1	
utin	e->7	m->1	
utio	n->260	
utiq	u->1	
utit	 ->4	s->7	
utjä	m->5	
utka	n->1	s->15	
utko	m->3	n->1	
utkr	ä->3	
utla	n->5	
utli	g->72	
utlo	v->3	
utlä	g->1	m->2	n->4	
utlå	t->2	
utlö	s->2	
utma	n->20	
utmy	n->1	
utmä	r->32	
utna	 ->10	,->3	.->4	
utni	n->41	
utny	t->41	
utnä	m->4	
uto/	O->1	
utom	 ->78	,->2	a->8	e->3	o->7	s->2	
utop	i->1	
utor	 ->1	
utpe	k->1	r->1	
utpl	å->2	
utpr	e->1	ä->1	
utpu	n->1	
utra	l->2	
utre	 ->1	d->8	s->4	
utri	k->19	
utro	p->2	t->4	u->1	
utru	s->4	
utry	m->11	
uträ	t->2	
uts 	k->1	s->1	u->4	
uts-	b->1	
utsa	m->14	r->1	t->50	
utsc	e->1	h->1	
utse	 ->7	.->1	d->1	e->1	r->1	s->3	t->3	
utsf	a->11	ö->1	
utsi	g->1	k->1	
utsk	o->157	
utsl	a->15	ä->9	
utsp	r->4	
utsr	ä->1	
utst	a->11	r->28	ä->2	å->1	ö->1	
utsu	g->1	
utsä	g->2	t->61	
utså	g->3	
utta	 ->2	l->98	
utte	 ->1	n->1	
utti	g->1	t->1	
uttj	ä->24	
uttn	a->2	
utto	l->1	n->3	r->1	
uttr	y->72	ä->1	
uttö	m->5	
utva	l->1	p->1	r->2	
utve	c->237	r->4	
utvi	d->106	s->1	
utvä	r->32	
utyp	,->1	
utän	d->5	
utåt	"->1	
utök	a->11	n->1	
utöv	a->15	e->14	n->1	
uum 	o->1	
uumt	a->1	
uva 	i->1	
uvar	a->46	
uvel	e->2	
uver	g->1	n->1	ä->17	
uvid	a->15	
uvri	è->1	
uvud	 ->9	a->7	d->3	e->1	f->5	l->2	m->2	r->3	s->21	u->1	
ux, 	n->2	
ux-a	f->1	
uxem	b->6	
uxha	v->1	
uxit	 ->1	
uxna	 ->1	.->1	
uyu 	i->1	s->1	
v "p	a->1	
v "r	e->1	i->1	
v (K	O->1	
v - 	d->1	i->1	o->3	p->1	s->2	u->1	
v 14	 ->1	
v 19	 ->1	9->2	
v 20	0->1	
v 40	 ->1	
v 41	0->1	
v 5 	0->1	
v 54	0->1	
v 8 	4->1	
v 93	/->1	
v 94	/->2	
v 96	/->5	
v Ah	e->2	
v Am	e->1	s->1	
v Ar	a->1	
v BN	I->1	P->5	
v BS	E->1	
v Ba	r->2	
v Be	r->8	
v Bo	u->1	
v Br	o->2	
v Ca	n->1	
v Da	 ->1	v->1	
v De	m->1	
v Di	m->2	
v Du	b->1	
v Dü	h->1	
v EG	-->1	
v EU	 ->3	,->1	-->4	.->2	:->7	
v En	l->1	
v Er	i->1	
v Eu	r->70	
v Ex	x->2	
v FN	:->1	
v FP	Ö->2	
v Fl	o->1	
v Fö	r->8	
v Ga	z->1	
v Ge	n->2	
v Gr	a->2	o->1	
v Ha	i->1	
v He	n->1	
v Hi	t->1	
v Is	r->2	
v Ja	c->1	
v Je	r->1	
v Jo	n->2	
v Ki	n->3	
v Ko	c->3	s->7	
v Ku	l->1	
v La	n->3	
v Li	b->1	
v Lö	ö->1	
v Ma	r->2	
v Mc	N->1	
v Mo	r->1	
v OL	A->3	
v Os	m->1	
v Oz	 ->1	
v Pa	l->1	t->1	
v Po	r->1	
v Pé	t->1	
v Ra	p->1	
v Ri	i->1	
v Sa	m->1	
v Sc	h->6	
v Ta	c->1	
v Te	r->1	
v Th	e->3	y->1	
v Ti	b->1	
v To	t->1	
v UN	M->1	
v Va	n->1	r->1	
v Vä	s->1	
v Wa	l->1	
v Wi	e->1	
v Wy	e->1	
v ac	c->1	
v ad	m->1	v->1	
v ag	e->1	
v al	b->1	d->1	k->1	l->33	
v an	b->1	d->5	l->2	m->1	o->1	s->16	t->3	v->2	
v ap	r->2	
v ar	b->20	t->20	
v as	y->1	
v at	t->70	
v av	 ->15	,->1	.->1	f->1	g->4	p->1	s->2	t->2	v->2	
v ba	r->2	s->1	
v be	d->1	f->6	g->1	h->6	k->1	s->16	t->9	v->2	
v bi	d->3	l->11	o->1	
v bl	a->2	y->1	å->1	
v bo	l->1	m->2	
v br	e->1	i->4	o->4	u->1	
v bu	d->8	
v by	g->2	
v bå	d->2	
v bö	c->1	r->2	
v ce	n->2	
v ci	r->2	v->4	
v co	m->1	
v da	g->5	t->1	
v de	 ->165	b->3	f->1	l->3	m->27	n->183	r->6	s->45	t->128	
v di	p->1	r->21	s->6	v->1	
v dj	u->2	
v do	k->1	m->11	
v dr	i->1	
v dä	r->2	
v ef	f->2	t->3	
v eg	e->2	
v ek	o->12	
v en	 ->99	b->1	e->9	h->1	i->1	o->1	t->2	
v er	 ->9	,->2	:->1	a->3	f->1	t->2	
v et	n->1	t->51	
v eu	r->7	
v ev	e->1	
v ex	a->6	p->1	t->1	
v fa	k->3	l->3	r->39	t->4	
v fi	n->3	s->3	
v fj	o->2	
v fl	e->9	o->1	y->6	
v fo	l->1	n->1	r->6	
v fr	a->1	e->1	i->11	ä->5	å->18	
v fu	l->2	n->1	s->2	
v fy	s->1	
v fä	d->1	
v få	 ->1	n->1	r->3	
v fö	l->2	r->123	
v ga	m->3	
v ge	m->28	n->3	o->1	
v gi	f->1	g->1	v->1	
v gl	o->1	
v go	d->2	
v gr	a->2	o->1	u->3	ä->4	ö->1	
v gö	r->1	
v ha	 ->1	n->5	r->8	t->2	v->4	
v he	l->6	m->1	
v hi	e->1	g->1	s->3	
v hj	ä->1	
v ho	n->1	
v hu	n->1	r->7	
v hä	n->1	r->1	
v hö	g->2	r->1	
v i 	K->1	d->8	e->1	s->4	v->1	
v ib	e->1	
v ic	k->3	
v id	e->1	é->1	
v im	p->5	
v in	 ->1	d->1	e->1	f->4	i->2	n->3	o->2	r->2	s->5	t->13	v->3	
v jo	r->5	
v ju	r->1	s->3	
v jä	m->2	
v ka	m->2	n->4	p->1	r->3	t->3	
v kl	a->4	
v kn	u->1	
v ko	a->2	l->4	m->61	n->43	r->2	s->7	
v kr	i->4	ä->1	
v ku	l->4	s->1	
v kv	a->2	i->4	o->1	
v kä	r->8	
v la	g->12	n->8	s->1	
v le	d->10	g->1	j->1	
v li	b->2	c->1	k->2	s->3	v->8	
v lo	j->2	k->3	
v lä	g->1	m->1	n->2	t->1	
v lå	n->1	
v lö	s->1	v->1	
v ma	k->2	n->2	r->10	t->4	
v me	d->27	n->1	r->3	
v mi	g->2	l->14	n->18	s->3	t->3	
v mo	d->2	n->1	t->3	
v my	c->3	
v mä	n->7	
v må	l->3	n->4	s->1	
v mö	j->1	
v na	t->13	z->1	
v ni	 ->1	
v no	r->1	
v ny	 ->2	a->6	b->1	h->1	l->1	n->1	s->1	
v nä	r->1	s->1	
v nå	g->6	
v nö	d->2	
v oa	c->1	n->1	v->1	
v ob	e->3	l->1	
v oc	h->25	k->4	
v of	f->4	r->1	
v ok	l->1	
v ol	i->8	j->3	y->3	
v om	 ->25	b->1	e->1	f->1	k->1	r->2	s->2	
v on	d->1	
v op	i->1	
v or	d->7	i->1	k->1	s->2	
v os	s->12	
v ot	r->1	v->1	
v ou	n->1	
v ov	a->1	
v pa	k->1	l->1	r->20	
v pe	n->7	r->5	
v pi	o->1	
v po	l->9	
v pr	e->1	i->8	o->28	
v på	 ->31	v->2	
v ra	m->2	p->3	s->1	
v re	f->3	g->17	k->1	n->1	p->1	s->8	t->1	v->1	
v ri	k->5	s->3	
v ro	l->2	
v ry	s->1	
v rä	d->1	k->5	t->6	
v rå	d->12	
v rö	s->1	
v sa	k->1	m->15	
v sc	e->1	
v se	 ->1	d->1	g->1	k->2	n->1	r->1	s->2	x->1	
v si	d->1	g->3	n->13	s->1	t->7	
v sj	u->1	ä->1	ö->1	
v sk	a->10	e->1	o->4	r->3	u->1	ä->3	ö->1	
v sl	u->2	
v sm	å->2	
v sn	a->1	
v so	c->7	l->1	m->38	
v sp	e->1	l->1	
v st	a->24	i->2	o->14	r->16	y->1	ä->1	å->3	ö->20	
v su	b->3	c->1	
v sv	a->1	ä->1	
v sy	f->2	n->1	s->21	
v sä	g->1	k->9	r->5	
v så	 ->6	d->8	s->1	
v ta	 ->1	l->3	
v te	k->4	l->1	r->3	
v ti	d->2	l->36	m->2	
v tj	ä->28	
v to	t->2	
v tr	a->7	e->3	y->1	ä->2	
v tu	n->5	r->1	
v tv	u->1	å->1	
v ty	d->1	p->1	
v tä	n->1	
v un	d->8	g->2	i->20	
v up	p->6	
v ut	a->6	b->2	f->2	g->3	n->1	r->2	s->7	t->3	v->11	
v va	d->12	n->3	p->1	r->6	t->1	
v ve	d->1	r->3	t->6	
v vi	 ->1	c->4	d->1	k->3	l->7	s->9	t->1	
v vo	n->4	
v vä	g->1	l->3	n->2	r->8	x->6	
v vå	r->24	
v yt	t->5	
v Ös	t->2	
v äl	d->1	
v äm	n->1	
v än	 ->1	d->4	n->1	
v är	 ->9	
v ål	d->1	
v år	 ->6	e->1	h->1	
v ås	i->1	
v åt	e->4	g->12	
v öb	o->1	
v öd	e->1	
v ök	a->4	
v öp	p->4	
v ös	t->2	
v öv	e->4	
v", 	d->1	
v, 9	5->1	
v, a	n->1	t->2	
v, b	a->1	
v, d	e->3	v->1	ä->1	
v, e	f->1	n->2	
v, f	r->1	
v, h	a->1	e->2	y->1	
v, i	n->1	
v, j	a->1	
v, l	i->1	
v, m	e->4	i->1	
v, n	ä->1	å->1	
v, o	c->7	m->1	
v, s	o->4	t->1	ä->1	å->2	
v, t	i->1	r->1	
v, u	n->1	
v, ä	r->2	
v. D	e->1	
v. M	e->1	
v. V	a->1	i->1	
v. m	e->1	
v."D	e->1	
v.(S	a->1	
v., 	ä->1	
v.. 	(->2	
v..H	e->1	
v.?A	n->1	
v.At	t->1	
v.Av	 ->1	s->1	
v.Ba	r->1	
v.Bl	a->1	
v.De	 ->3	n->1	t->7	
v.Dä	r->1	
v.Då	 ->1	
v.Ef	f->1	
v.En	 ->2	
v.Er	i->1	
v.Fr	u->1	
v.Fö	r->4	
v.He	r->1	
v.I 	d->1	v->1	
v.In	g->1	
v.Ja	g->2	
v.Ko	m->1	
v.Lå	t->1	
v.Me	n->3	
v.OL	A->1	
v.Om	 ->1	
v.Ri	k->1	
v.Rå	d->1	
v.Sv	e->1	
v.Så	s->1	
v.Up	p->1	
v.Vi	 ->2	s->1	
v.Yt	t->1	
v: F	ö->1	
v: v	å->1	
v; a	n->1	
v?Fö	r->1	
v?Ne	j->1	
v?Vi	l->1	
va 4	0->1	
va E	u->2	
va a	n->5	r->1	t->7	v->5	
va b	a->1	e->5	i->3	j->1	o->2	r->1	ä->1	
va c	e->1	
va d	a->1	e->18	r->1	u->2	ä->1	
va e	f->7	n->17	t->2	u->1	x->1	
va f	a->3	i->1	l->1	u->1	ö->10	
va g	a->1	ä->1	ö->3	
va h	a->3	u->2	ö->1	
va i	 ->9	d->1	g->1	m->1	n->3	
va j	u->1	
va k	a->4	l->2	o->7	r->3	u->1	ä->4	
va l	a->1	e->1	i->2	ö->1	
va m	e->4	i->1	o->1	å->2	
va n	i->1	å->4	
va o	c->13	f->1	m->1	r->3	
va p	a->2	o->4	r->2	u->1	å->6	
va r	a->1	e->6	i->1	o->1	u->1	ä->1	å->1	
va s	a->3	e->1	i->3	j->1	k->2	l->1	o->2	t->3	v->1	y->3	
va t	e->2	i->14	r->1	v->1	
va u	n->1	p->2	r->1	t->3	
va v	e->29	ä->2	å->2	
va ä	r->2	
va å	r->2	s->1	t->5	
va ö	k->2	v->1	
va, 	d->1	f->1	i->1	s->3	u->2	ä->1	
va.A	l->1	
va.D	e->1	
va.H	e->1	
va.L	å->1	
va.N	ä->1	
va.O	m->1	
va.V	a->1	å->1	
va?N	e->1	
vack	e->2	l->1	r->6	
vad 	B->1	E->1	G->1	K->2	S->1	a->1	b->14	d->30	e->3	f->3	g->47	h->4	i->1	j->7	k->8	m->9	n->5	o->3	p->1	r->2	s->60	t->1	v->27	ä->6	
vad?	D->1	
vade	 ->9	.->1	s->2	
vag 	i->1	p->1	s->1	
vaga	 ->10	,->2	d->3	r->6	s->7	t->2	
vagh	e->12	
vagn	e->2	i->1	
vagt	.->1	
vaka	 ->10	.->1	r->5	s->2	t->1	
vaki	e->1	
vakn	i->14	
vaks	a->9	
vakt	 ->1	a->6	e->1	
vaku	u->2	
val 	a->22	d->1	e->1	f->1	g->1	i->2	l->1	m->1	s->2	u->1	ä->1	å->1	
val,	 ->3	
val.	D->1	I->1	M->1	S->1	V->1	
val;	 ->1	
vala	r->3	
valb	a->1	
vald	 ->8	.->1	a->16	e->8	i->1	
vale	n->6	s->1	t->6	
valf	r->5	
vali	f->15	t->36	
valk	r->4	
vall	f->1	p->1	
valr	e->1	
vals	k->1	
valt	 ->5	,->1	a->3	i->1	n->47	s->4	
valu	t->23	
van 	D->2	G->1	H->20	V->1	a->3	d->9	e->3	m->1	o->1	
van,	 ->1	
van.	D->1	T->1	
vana	 ->2	
vanc	e->1	
vand	a->1	e->36	l->9	r->18	
vanh	e->2	
vani	f->1	
vanl	i->12	
vann	ä->2	
vano	r->1	s->2	
vanp	å->1	
vans	 ->4	,->4	e->1	i->1	k->3	t->1	v->1	
vant	 ->4	a->6	i->8	
vape	n->26	
vapn	e->2	
var 	-->2	1->5	9->1	K->1	W->1	a->25	b->14	d->37	e->36	f->40	g->5	h->8	i->26	j->4	k->6	l->6	m->18	n->11	o->15	p->25	r->5	s->27	t->8	u->3	v->11	ä->7	ö->4	
var,	 ->30	
var.	 ->1	D->14	E->1	F->1	G->3	I->2	J->5	M->4	N->1	O->1	P->1	R->1	S->3	V->5	
var;	 ->1	
var?	I->1	
vara	 ->388	"->1	,->2	.->4	:->1	d->11	k->4	n->122	r->35	s->2	t->6	v->4	
vard	a->4	e->1	
vare	 ->48	"->2	,->5	.->7	f->1	n->11	s->1	t->72	
varf	ö->39	
varg	a->1	
varh	ä->1	å->2	
vari	 ->1	e->2	g->62	t->71	
varj	e->84	
vark	e->14	o->1	
varl	i->62	ä->1	
varm	a->3	t->12	
varn	a->23	i->7	
varo	 ->4	,->1	n->3	r->2	
varp	a->1	
varr	 ->1	
vars	 ->28	.->1	a->2	b->3	f->55	k->4	l->1	m->3	o->7	p->5	t->10	
vart	 ->4	a->5	e->1	
varv	,->1	e->1	i->3	s->3	
vas 	a->8	e->3	f->1	h->1	i->3	m->2	o->4	s->1	
vas,	 ->2	
vas.	C->1	G->1	H->1	I->1	M->1	V->1	
vast	e->1	
vat 	-->1	E->1	a->2	b->1	d->2	e->1	f->1	o->1	r->1	t->1	u->1	
vat.	J->1	Å->1	
vata	 ->18	
vate	k->1	
vati	o->8	s->2	v->9	
vats	 ->4	,->1	.->1	
vatt	e->33	n->16	
vatö	r->1	
vavt	a->7	
vbes	t->3	
vbet	ä->1	
vbio	g->1	
vbor	d->1	
vbri	n->1	
vbro	t->4	
vbru	t->2	
vbry	t->3	
vbrö	t->6	
vbär	a->1	
vda 	a->6	d->1	
vdad	e->3	
vdar	 ->10	,->1	.->1	
vdat	 ->4	.->1	
vde 	d->1	e->1	f->1	g->2	
vde,	 ->1	
vdel	n->8	
vdes	 ->2	
vdvu	n->1	
ve (	C->2	
ve 1	9->1	
ve E	u->1	
ve a	l->1	n->1	
ve b	e->3	u->1	
ve d	e->4	
ve e	n->1	t->2	
ve f	o->1	
ve k	a->1	o->3	
ve l	a->2	
ve m	y->2	å->1	
ve p	a->3	
ve r	e->1	u->1	ä->1	
ve s	j->1	
ve t	i->1	r->1	
ve ä	r->1	
ve, 	a->1	å->1	
ve- 	p->1	
ve-p	r->2	
veNä	s->1	
vebr	ö->1	
vec 	l->1	
veck	a->24	l->248	o->17	
vede	r->13	
vek 	h->1	o->1	
veka	 ->3	d->1	n->15	r->3	t->2	
vekh	e->4	
vekl	ö->1	
veko	n->1	
veks	a->5	
vel 	a->7	g->3	l->1	n->1	o->6	p->1	s->1	t->2	u->1	v->1	ä->2	
vel,	 ->2	
vela	k->3	t->7	
vele	n->1	r->1	
vels	e->6	u->3	
vem 	b->1	f->1	i->1	s->13	ä->1	
vemb	e->11	
vems	 ->1	
ven 	-->1	7->1	E->4	G->1	R->2	a->17	b->4	d->22	e->12	f->29	g->2	h->7	i->51	j->13	k->11	l->4	m->19	n->9	o->88	p->17	r->3	s->12	t->12	u->7	v->6	y->1	ä->5	ö->3	
ven,	 ->4	
ven.	D->2	K->1	N->1	S->2	T->2	V->1	
ven:	 ->1	
vene	m->1	r->2	
venh	e->4	
vens	 ->5	.->1	e->41	k->3	
vent	 ->10	,->2	a->5	e->1	i->42	u->21	y->9	
vep 	a->1	
vepe	s->1	
veps	k->1	
vept	e->1	
ver 	-->2	1->1	2->1	3->2	4->1	5->1	7->1	8->2	9->1	B->1	E->5	H->1	O->1	a->58	b->3	d->48	e->40	f->14	g->14	h->38	i->11	j->5	k->10	l->4	m->15	n->9	o->12	p->7	r->9	s->22	t->7	u->11	v->32	y->1	Ö->1	ä->4	å->1	
ver,	 ->8	
ver.	 ->1	D->2	H->1	J->1	K->2	M->1	O->1	S->2	T->1	V->2	
vera	 ->6	d->10	l->9	n->7	r->7	s->2	t->2	
verb	a->1	e->4	l->1	r->4	
verc	e->1	
verd	r->14	
vere	n->71	r->5	t->1	
verf	a->3	i->1	l->3	ö->16	
verg	e->15	i->2	n->1	r->14	å->15	
verh	a->1	e->1	ä->1	ö->2	
veri	 ->5	,->1	e->2	f->1	g->7	n->7	
verk	 ->27	,->3	.->4	?->1	a->203	e->46	l->211	n->15	s->70	t->8	
verl	a->1	e->5	ä->21	å->8	
verm	o->2	
vern	a->3	i->1	ö->1	
vero	r->1	
verp	r->1	
verr	a->1	e->2	ö->1	
vers	,->1	a->2	e->7	i->35	k->23	t->9	v->7	y->1	ä->11	
vert	a->6	i->3	o->2	r->7	y->38	ä->1	
verv	a->25	i->8	u->1	ä->38	
very	,->1	
verä	n->17	
ves 	h->1	o->1	
vest	e->15	o->3	
vet 	"->1	-->2	E->8	L->1	S->1	a->77	b->3	f->12	g->5	h->11	i->19	j->3	k->4	m->6	n->5	o->21	p->11	r->2	s->13	t->2	u->7	v->10	ä->12	
vet"	 ->1	
vet,	 ->28	
vet.	 ->1	D->7	E->2	F->3	H->1	I->1	J->4	M->2	N->1	R->1	S->1	T->1	V->1	
veta	 ->27	,->1	n->4	
vete	n->85	r->12	t->8	
vetn	a->17	
vets	 ->12	s->1	
vett	e->1	i->3	v->1	
vetv	i->27	
vety	d->7	
veur	o->1	
vfal	l->25	
vfol	k->1	
vför	d->1	m->1	s->4	t->2	
vgas	e->1	
vgav	 ->1	
vge 	e->3	
vger	 ->5	
vges	 ->1	
vget	t->1	
vgic	k->4	
vgif	t->4	
vgiv	i->1	
vgjo	r->4	
vgrä	n->4	
vgå.	S->1	
vgåe	n->1	
vgån	g->3	
vgår	 ->1	
vgåt	t->1	
vgör	 ->1	a->57	s->3	
vhet	 ->1	
vhjä	l->3	r->1	
vhän	d->1	g->1	
vhål	l->1	
vi -	 ->3	
vi 1	9->1	
vi 5	5->1	
vi E	u->2	
vi I	n->1	
vi L	i->1	
vi P	r->1	
vi a	)->1	b->3	c->1	g->2	l->37	n->30	r->6	t->41	v->7	
vi b	a->5	e->54	i->3	l->6	o->10	r->2	y->1	ö->27	
vi d	a->1	e->26	i->15	o->1	r->1	ä->6	å->6	
vi e	f->5	g->3	k->1	m->5	n->14	r->3	t->9	u->2	v->1	x->1	
vi f	a->14	i->2	o->13	r->6	u->3	å->18	ö->41	
vi g	a->1	e->15	i->1	j->4	l->4	o->4	r->2	ä->2	ö->19	
vi h	a->135	e->7	i->5	j->1	o->4	ä->14	å->7	ö->2	
vi i	 ->56	a->1	b->2	g->1	n->134	
vi j	u->11	
vi k	a->65	l->2	n->1	o->41	r->4	u->7	v->1	ä->2	
vi l	a->3	i->7	o->1	y->5	ä->9	å->2	
vi m	e->20	i->3	o->3	y->1	å->63	
vi n	a->4	u->21	y->2	ä->6	å->2	
vi o	b->1	c->31	f->2	m->1	s->9	
vi p	l->2	r->1	å->12	
vi r	e->13	i->2	o->1	u->2	ä->2	å->1	ö->7	
vi s	a->6	e->17	j->4	k->68	l->3	n->8	o->16	p->2	t->24	v->1	y->2	ä->6	å->4	
vi t	.->1	a->24	e->1	i->15	o->1	r->8	v->1	y->7	ä->4	
vi u	n->7	p->17	r->1	t->13	
vi v	a->9	e->22	i->34	ä->6	å->3	
vi y	t->1	
vi ä	g->4	n->10	r->28	v->5	
vi å	l->1	r->1	s->1	t->4	
vi ö	n->5	v->3	
vi, 	g->1	j->3	k->1	l->1	m->1	n->1	s->5	t->1	ä->2	
vi.V	i->1	
vi?.	H->1	
via 	B->1	E->1	R->1	a->1	b->1	d->1	e->1	k->1	o->1	s->1	t->1	u->1	
vian	o->1	
vic 	i->1	
vice	 ->13	.->4	k->2	n->1	
vick	s->3	
vid 	1->1	7->1	B->3	E->6	G->1	H->1	K->1	L->1	M->1	P->1	a->14	b->7	d->35	e->15	f->21	g->3	h->6	i->1	j->2	k->8	l->1	m->5	n->5	o->8	p->9	r->5	s->17	t->12	u->14	v->8	å->2	ö->2	
vid,	 ->2	
vid.	H->1	J->1	
vida	 ->21	r->37	
vidd	 ->3	.->1	e->1	
vide	r->22	
vidg	a->38	n->71	
vidh	å->4	ö->1	
vidl	a->1	
vidm	a->1	
vids	t->1	
vidt	a->62	o->2	
vidu	a->1	e->7	
vien	n->1	s->1	
vier	 ->1	
vift	a->1	
vig 	v->1	
vigl	a->1	
vigt	 ->1	,->1	.->1	
vigv	a->1	
vigö	r->1	
vika	 ->27	n->4	s->4	
vike	l->5	n->2	r->6	t->1	
viki	t->1	
vikl	i->4	
vikn	a->1	
vikt	 ->15	,->2	.->2	;->1	e->12	i->328	n->3	s->2	
vil 	e->2	s->3	
vil-	 ->1	
vila	 ->3	r->3	
vilb	e->2	
vild	a->1	
vile	g->6	
vilf	ö->2	
vili	g->1	s->2	
vilj	a->227	e->2	
vilk	a->90	e->227	
vill	 ->529	,->8	.->2	e->10	i->20	k->63	o->1	
vilr	ä->1	
vils	e->3	k->2	
vilt	 ->1	,->1	
vin 	E->1	o->1	
vind	 ->1	f->4	
ving	a->32	
vini	s->1	
vink	e->11	l->1	
vinn	a->29	e->18	i->49	l->2	o->61	s->2	
vins	 ->2	e->1	t->12	
virk	e->3	
virr	a->4	i->8	v->1	
vis 	-->3	A->1	G->1	a->23	b->9	d->9	e->7	f->14	g->9	h->12	i->22	k->6	l->3	m->11	n->1	o->24	p->11	r->3	s->27	t->3	u->5	v->10	ä->18	å->2	ö->3	
vis)	 ->1	
vis,	 ->17	
vis.	 ->1	D->2	E->1	H->1	J->1	M->1	S->1	Ä->1	
visa	 ->65	,->8	.->14	?->1	d->19	n->8	r->71	s->10	t->38	v->1	
visb	a->1	e->9	ö->7	
visd	o->1	
vise	n->3	r->9	t->8	
visf	i->3	
vish	e->3	
visi	o->24	
visk	 ->1	a->1	v->2	
vism	 ->1	
visn	i->14	
viso	r->5	
viss	 ->35	a->130	e->11	h->4	o->6	t->10	
vist	 ->15	,->1	a->4	e->7	
visu	a->1	e->1	m->1	
vit 	a->2	b->2	d->1	e->8	f->2	g->1	h->1	i->1	l->3	m->1	o->1	s->7	t->2	u->6	v->1	
vit.	F->1	
vitb	o->50	
vite	t->39	
vits	 ->9	,->1	
vitt	 ->2	n->5	
vive	l->33	
vivl	a->10	
vjas	 ->1	
vjet	t->1	
vju 	m->1	s->1	
vjua	d->1	
vkar	t->1	
vkla	r->21	
vkon	s->1	
vkos	t->1	
vkra	f->3	
vkrä	v->1	
vkun	n->1	
vla 	d->1	f->1	s->1	v->1	ä->1	
vla"	 ->2	
vla.	V->1	
vlad	e->4	
vlag	t->1	
vlan	"->1	
vlar	 ->6	
vlat	 ->2	
vled	d->2	
vlig	 ->2	.->1	a->3	e->1	h->1	t->2	
vlin	g->1	
vlis	t->2	
vliv	a->1	
vlop	p->1	
vläg	g->1	s->9	
vlåd	e->1	
vmat	t->1	
vmil	j->1	
vna 	a->1	b->3	c->1	f->2	i->1	ä->1	
vnad	 ->4	,->2	.->1	?->1	e->2	s->6	
vnin	g->36	
vo (	K->2	
vo T	r->1	
vo a	t->1	
vo b	ä->1	
vo f	r->1	ö->2	
vo h	a->1	
vo i	n->1	
vo k	a->1	ä->1	
vo m	e->1	
vo o	c->7	
vo t	i->1	
vo u	t->1	
vo v	a->1	
vo ä	r->3	
vo, 	e->2	h->1	i->1	m->2	o->3	s->1	v->1	
vo.-	 ->1	
vo.A	v->1	
vo.D	e->2	
vo.E	u->1	
vo.F	ö->1	
vo.H	e->1	
vo.K	o->1	
vo.L	å->1	
vo.M	e->1	
vo.O	c->1	
vo.V	i->1	
vo? 	D->1	
vo?H	u->1	
voNä	s->1	
voff	e->1	
voka	t->5	
voko	n->1	
vokr	i->1	
volu	n->4	t->1	
volv	e->9	
voly	m->4	
von 	B->1	E->1	W->16	
vor 	t->1	
vor.	L->1	
vord	a->2	
vore	 ->29	
vori	t->1	
vos 	a->1	d->1	e->1	l->1	m->1	s->1	y->1	
vot 	p->1	s->1	v->1	ä->1	
vot!	D->1	
vot,	 ->1	
vote	n->3	r->10	
votu	m->1	
voår	 ->1	
vplå	g->1	
vpri	c->1	
vrad	e->1	
vrak	 ->4	,->1	.->2	?->1	e->2	
vran	d->1	
vrap	p->1	
vrar	,->1	
vras	,->1	
vred	g->1	
vreg	l->2	
vrid	a->1	e->6	n->7	
vrig	 ->1	a->33	t->32	
vrik	 ->1	
vriè	r->1	
vrun	d->1	
vräk	t->1	
vrän	g->2	
vrät	t->5	
vs a	v->6	
vs b	e->1	
vs d	e->13	r->1	
vs e	f->1	g->1	n->16	t->2	
vs f	r->1	ö->9	
vs g	e->1	
vs h	a->3	
vs i	 ->10	n->3	
vs k	r->1	
vs m	e->3	y->1	
vs n	å->1	
vs o	c->3	m->1	
vs p	r->1	å->1	
vs r	a->1	
vs s	k->1	o->4	p->1	t->1	ä->1	å->2	
vs u	p->1	t->2	
vs v	e->2	i->2	
vs ä	r->1	
vs ö	v->1	
vs, 	f->2	m->4	o->2	s->2	
vs. 	1->2	E->1	W->1	a->11	d->4	e->3	f->3	g->1	h->2	i->5	j->1	m->4	n->1	o->2	p->1	s->1	v->2	
vs.A	l->1	
vs.D	e->3	
vs.E	t->2	
vs.F	r->1	
vs.I	 ->1	
vs.R	e->1	
vs.S	a->1	l->1	
vs.V	i->1	
vs?T	i->1	
vsak	n->4	
vsar	b->3	
vsat	t->4	
vscy	k->3	
vsdu	g->2	
vse 	f->1	
vsed	d->3	
vsee	n->47	
vser	 ->15	
vses	 ->1	
vset	t->14	
vsev	ä->14	
vsfo	r->1	
vsfö	r->1	
vsid	a->1	e->1	
vsik	t->38	
vsin	d->1	
vska	f->19	
vske	d->5	
vski	l->1	
vsko	g->1	n->2	
vskr	a->1	ä->2	
vskv	a->5	
vsky	 ->1	v->1	
vsla	g->2	
vslo	g->2	
vslu	t->74	
vslä	n->2	
vslå	 ->2	r->1	
vslö	j->6	
vsma	n->2	
vsme	d->88	
vsmi	l->5	
vsmä	n->3	
vsni	t->4	
vsom	r->1	
vspe	g->5	
vsst	ö->2	
vsta	 ->1	m->1	
vste	s->1	
vsto	d->2	
vsty	m->1	r->6	
vstä	n->11	
vstå	 ->7	e->1	n->11	r->5	t->2	
vsup	p->1	
vsva	t->1	
vsvi	l->1	
vsäg	a->1	
vsäk	e->1	
vsät	t->4	
vt -	 ->1	
vt a	n->1	r->3	t->7	
vt b	e->3	l->1	
vt d	e->3	i->1	
vt e	l->1	n->2	t->1	
vt f	r->1	u->1	ö->6	
vt h	a->2	ö->1	
vt i	 ->4	n->5	
vt k	a->3	o->1	
vt m	e->2	o->1	y->1	
vt n	å->1	
vt o	c->12	m->4	t->1	
vt p	r->2	å->4	
vt r	e->2	ä->2	
vt s	a->2	e->2	i->1	k->2	n->1	o->2	p->1	t->5	v->2	ä->15	
vt t	a->1	i->6	
vt u	t->2	
vt v	e->1	
vt y	t->1	
vt ä	r->1	
vt å	l->2	r->2	
vt ö	k->1	
vt, 	d->2	i->1	m->1	o->1	p->1	r->1	
vt. 	D->1	
vt.D	e->2	
vt.E	n->1	
vt.I	n->1	
vt.P	a->1	
vt.Ä	v->1	
vtal	 ->51	"->1	,->2	.->5	:->1	e->28	s->1	
vtar	.->1	
vtid	s->1	
vtim	m->2	
vtru	p->1	
vts 	d->1	ä->1	
vts.	E->1	
vtvi	n->1	
vud 	t->9	
vuda	k->2	n->5	
vudd	e->3	
vude	t->1	
vudf	r->4	ö->1	
vudl	i->2	
vudm	å->2	
vudr	e->1	o->2	
vuds	a->16	t->4	y->1	
vudu	p->1	
vule	n->1	
vuls	k->1	
vund	s->1	
vung	e->5	n->6	
vunn	a->2	e->2	i->7	
vuxi	t->1	
vuxn	a->2	
vvak	t->6	
vvec	k->8	
vver	k->2	
vvik	a->4	e->4	
vvis	a->13	n->2	
vväg	d->2	n->1	s->2	
vvär	d->2	
vytt	r->1	
väck	a->10	e->5	s->1	t->7	
väde	r->2	
vädj	a->9	
vädr	e->1	
väg 	[->1	a->8	b->1	e->6	f->2	g->2	h->2	i->2	k->1	m->2	o->2	s->1	t->1	ä->1	å->1	
väg,	 ->16	
väg.	A->1	B->1	D->1	E->1	J->1	M->2	O->1	V->1	
vägN	ä->1	
väga	 ->19	,->1	.->1	g->6	n->8	r->20	
vägb	y->1	
vägd	 ->2	a->1	
väge	n->17	r->10	
vägg	i->3	
vägl	e->5	
vägm	ä->1	
vägn	a->16	i->1	
vägr	a->22	ö->1	
vägs	 ->2	k->2	n->2	o->1	
vägt	 ->2	
väka	r->1	
väkt	a->2	
väl 	S->1	a->9	b->3	d->5	e->3	f->7	g->2	h->4	i->11	k->5	l->1	m->9	o->2	p->3	r->3	s->10	t->3	u->10	v->4	ä->3	å->1	ö->1	
väl,	 ->2	
väl.	J->1	M->1	S->1	
välb	e->1	
väld	i->23	
välf	u->1	ä->8	
välg	r->2	ö->1	
välj	a->17	e->5	
välk	l->1	o->50	ä->3	
väll	 ->2	,->2	.->2	?->1	a->1	e->3	
välm	e->2	å->2	
väls	i->1	t->7	
vält	 ->1	a->2	s->1	
välu	t->3	
välv	a->1	n->3	
väml	i->15	
vämm	a->3	
vämn	i->4	
vämt	 ->1	
vän 	o->1	
vänd	 ->4	a->74	b->9	e->41	i->125	n->63	p->5	s->20	
vänl	i->15	
vänn	e->3	
väns	k->1	t->15	
vänt	 ->8	a->68	n->7	s->5	
väpn	a->2	
värd	 ->12	.->1	a->20	e->108	i->27	
väre	t->1	
värl	d->55	i->6	
värn	a->3	
värp	o->2	
värr	 ->36	,->2	.->1	a->4	e->6	
värs	 ->1	t->8	
värt	 ->18	,->3	.->3	o->17	
värv	a->4	s->3	
väse	n->36	
väst	k->1	r->2	v->1	
väts	k->1	
vätt	 ->1	,->2	.->1	a->1	
väva	 ->2	
vävn	a->4	
vävt	 ->1	
växa	 ->1	.->2	n->6	
växe	l->3	r->7	
växl	a->2	i->2	
växt	 ->7	,->2	.->2	b->1	e->10	h->7	s->3	
vå -	 ->1	
vå a	k->1	l->1	s->2	v->9	
vå b	e->2	o->1	
vå d	a->1	e->1	ä->1	
vå e	l->2	t->1	u->2	x->2	
vå f	a->3	i->1	l->1	o->1	r->4	ö->18	
vå g	e->2	r->1	å->1	
vå h	a->2	u->1	
vå i	 ->3	n->3	r->1	
vå j	o->1	
vå k	o->2	r->1	ä->1	
vå l	a->1	i->1	
vå m	e->3	i->4	y->1	å->3	ö->1	
vå n	e->1	y->1	ä->1	
vå o	c->5	f->1	l->1	m->1	r->1	
vå p	e->1	r->3	u->8	å->2	
vå r	e->1	ö->1	
vå s	a->3	e->2	k->2	m->1	o->8	t->3	ä->1	å->1	
vå t	i->5	r->2	y->1	
vå u	n->1	p->2	t->3	
vå v	e->1	i->6	
vå y	t->1	
vå ä	n->2	r->1	
vå å	r->7	s->1	
vå, 	a->1	b->2	d->1	f->2	g->1	m->1	o->2	r->2	v->1	
vå.A	t->1	
vå.B	i->1	r->1	
vå.D	e->6	ä->1	
vå.F	ö->1	
vå.G	e->1	
vå.H	e->2	
vå.J	a->3	ä->1	
vå.M	e->1	
vå.N	ä->1	
vå.P	å->1	
vå.V	i->1	
vå: 	d->2	
vå; 	d->1	
vå?S	e->1	
vådl	i->1	
våer	 ->6	,->2	.->4	:->1	n->1	
våg 	a->2	
våga	r->5	t->1	
våge	n->1	r->1	
vågl	ä->1	
vågr	u->3	
våhu	n->1	
våld	 ->2	e->2	s->6	t->2	
våll	a->1	
vån 	-->1	f->1	i->2	m->1	p->3	
vån.	D->3	H->1	
våna	 ->1	d->3	n->1	r->11	s->1	
vång	 ->1	r->1	s->5	
våni	n->2	
vår 	a->2	b->9	d->12	e->3	f->13	g->15	i->4	k->8	l->6	m->10	n->1	o->2	p->9	r->10	s->18	t->4	u->9	v->5	å->4	ö->1	
vår,	 ->1	
våra	 ->169	,->1	r->5	
vårb	e->2	
vård	 ->2	)->1	,->1	s->4	
våre	t->2	
våri	g->31	
vårl	ö->2	
vårs	s->2	
vårt	 ->132	,->2	
vårö	v->1	
vö, 	f->1	
vö.D	e->1	
vön 	s->1	
vörd	n->1	
w Yo	r->1	
w fö	r->1	
w ti	l->1	
w, s	o->1	
w-ho	w->1	
w.Me	d->1	
wage	n->1	
wald	,->1	
wale	s->1	
wan 	i->1	
warz	w->1	
we.E	u->1	
we.V	i->1	
webb	p->1	
weiz	,->1	
well	s->1	
wer 	k->1	
wer,	 ->2	
wies	 ->1	
will	 ->1	
wis 	h->1	n->1	
witt	s->1	
witz	.->1	
wn a	v->1	
wn ä	r->1	
wn, 	m->1	
wobo	d->3	
wood	 ->1	f->1	s->1	
wors	t->1	
x al	l->1	
x an	t->4	
x av	 ->1	s->1	
x ef	t->1	
x eu	r->1	
x fl	e->1	
x in	n->1	
x mi	n->1	
x må	n->10	
x oc	h->1	
x pl	a->1	
x po	s->1	
x sa	d->1	
x ti	l->1	
x tu	n->1	
x öv	e->1	
x!Ja	g->1	
x, j	a->1	
x, n	o->1	ä->1	
x, s	j->1	o->1	
x-af	f->1	
x-fr	e->3	
x. E	u->1	
x. F	r->1	
x. N	e->1	
x. U	S->1	
x. a	t->1	v->1	
x. d	e->2	
x. e	t->1	
x. i	n->1	
x. k	u->1	ä->1	
x. m	i->2	
x. n	ä->2	
x. o	l->1	
x. p	å->1	
x. u	t->1	
x. v	a->1	
x.De	 ->1	
x.Ja	g->1	
xa e	t->1	
xa u	t->2	
xa, 	t->1	
xa.H	ä->1	
xa.M	e->1	
xakt	 ->10	,->1	a->6	h->1	
xal 	s->2	
xala	 ->1	
xalt	 ->2	
xame	n->6	
xami	n->10	
xan?	V->1	
xand	e->8	
xas 	d->5	g->1	i->1	
xat 	u->1	
xbel	o->1	
xcep	t->6	
xelk	u->1	
xelr	y->1	
xelv	e->2	
xemb	u->6	
xemp	e->110	l->8	
xen 	s->1	
xer 	d->1	f->1	o->2	s->2	
xer,	 ->1	
xeri	n->1	
xfic	k->1	
xhav	e->1	
xibe	l->11	
xibi	l->10	
xibl	a->6	
xid 	i->1	o->3	
xidu	t->1	
xiko	,->1	
xilr	e->1	
xilt	i->1	
xima	l->6	
xime	r->2	
ximi	å->1	
xin 	o->1	
xink	r->1	
xis 	a->1	i->1	s->2	ä->1	
xis.	D->1	F->1	
xise	n->1	
xisk	a->1	
xism	e->1	
xist	e->19	
xit 	u->1	
xklu	s->3	
xlan	d->1	
xlar	 ->1	.->1	
xlin	g->2	
xmån	a->1	
xna 	e->1	
xna.	H->1	
xnin	g->1	
xon 	V->3	
xor.	D->1	
xpan	d->5	s->1	
xped	i->1	
xper	t->46	
xpli	c->1	
xplo	s->2	
xpon	e->2	
xpor	t->4	
xt a	v->2	
xt f	å->1	
xt i	 ->1	
xt k	o->1	
xt l	i->1	
xt o	c->6	m->1	
xt s	k->1	o->5	
xt ä	r->1	
xt, 	i->1	o->1	s->4	ä->1	
xt.K	o->1	
xt.M	e->1	
xt.O	c->1	
xtbr	a->1	
xten	 ->17	"->2	,->4	.->2	
xter	 ->3	,->2	.->3	n->11	
xthu	s->7	
xton	.->1	
xtra	 ->5	n->1	o->1	
xtre	m->30	
xtsk	y->3	
xuel	l->3	
xupé	r->1	
xvär	t->1	
xxon	 ->3	
y - 	s->1	
y Ca	n->3	
y Eu	r->1	
y Fo	r->1	
y bi	l->1	
y de	n->1	t->3	
y en	d->1	l->1	
y eu	r->1	
y fa	s->1	
y fo	r->1	
y fö	r->6	
y gr	a->1	
y ha	n->1	r->1	
y hä	r->1	
y i 	h->1	
y in	f->1	g->1	s->1	
y ke	m->1	
y ko	m->3	
y ku	l->3	
y kv	a->1	
y la	g->1	
y le	d->1	
y li	v->1	
y my	n->1	
y na	t->1	
y nä	r->1	
y oc	h->3	
y ol	j->1	
y pe	r->2	
y på	 ->2	
y rö	s->2	
y se	k->1	
y si	t->1	
y so	m->1	
y sp	e->1	
y st	o->1	
y sy	n->1	s->1	
y ty	p->1	
y un	d->1	
y up	p->1	
y va	r->1	
y ve	t->1	
y vi	 ->4	g->1	t->1	
y är	 ->1	
y åt	e->1	
y! G	e->1	
y, H	a->1	
y, J	o->1	
y, a	t->1	
y, d	e->1	
y, h	a->1	
y, k	a->1	v->1	
y, s	o->1	t->1	
y-pr	o->1	
y.An	d->1	
y.De	 ->1	
y.Vi	 ->2	
yDe 	f->1	
ya "	l->1	
ya 8	1->1	
ya E	U->1	u->2	
ya Z	e->2	
ya a	r->9	t->1	v->2	
ya b	e->6	i->6	u->1	y->1	
ya d	e->2	i->2	o->1	
ya e	u->1	x->1	
ya f	e->1	r->3	ö->6	
ya g	e->2	r->1	
ya i	m->1	n->3	
ya j	o->1	
ya k	l->1	o->16	
ya l	a->1	e->1	i->1	ä->4	
ya m	a->1	e->8	i->1	o->1	y->2	å->1	ö->3	
ya n	o->1	ä->1	
ya o	b->1	c->2	m->2	r->1	
ya p	a->1	e->3	r->9	
ya r	a->1	e->11	i->2	u->1	ä->2	
ya s	i->1	p->1	y->4	ä->1	
ya t	e->4	i->1	j->2	y->1	
ya u	p->1	t->2	
ya v	e->2	i->1	å->1	
ya ä	n->2	
ya å	r->1	t->5	
ya, 	u->1	
ya; 	k->1	
yabe	r->1	
yabu	k->2	
yago	l->4	
yal 	U->1	
yand	e->1	
yann	a->2	
yans	e->1	t->2	
yar 	l->1	
yarb	e->1	
yas 	o->1	
yast	e->1	
yavt	a->1	
ybar	 ->4	,->1	a->34	
ybet	ä->2	
ybil	a->1	s->2	
yck 	a->7	e->1	f->10	i->2	k->1	m->1	p->1	s->1	
yck,	 ->2	
yck.	D->1	
ycka	 ->35	,->2	.->1	?->1	d->13	n->14	s->26	t->20	
yckb	ä->1	
ycke	 ->7	.->3	l->8	n->3	r->67	t->464	
yckl	a->2	e->4	i->28	
yckn	i->5	
ycko	r->16	s->1	
ycks	 ->11	b->1	d->3	f->2	r->2	ö->1	
yckt	 ->4	e->16	s->1	
yckö	n->5	
ycli	n->1	
yd g	e->1	
yd i	 ->1	
yd s	o->1	
yd t	i->1	
yd.S	a->1	
yda 	m->1	u->2	
ydaf	r->2	
ydan	a->1	d->17	
ydd 	a->4	b->1	e->1	f->13	i->2	m->3	o->3	s->4	v->2	ö->1	
ydd)	,->1	
ydd,	 ->3	
ydd.	D->2	J->1	N->1	R->1	V->1	
ydda	 ->25	d->2	n->1	r->2	s->2	
ydde	 ->2	s->1	t->18	
ydds	m->4	n->6	o->2	p->1	s->2	t->1	
ydel	 ->1	s->75	
yder	 ->25	,->1	:->1	
ydeu	r->1	
ydig	 ->1	a->3	h->4	t->3	
ydko	r->1	
ydku	s->1	
ydli	g->125	
ydos	t->2	
yds 	i->1	
ydvä	s->1	
ydös	t->1	
ye P	l->1	
ye o	r->1	
ye-a	v->2	
yed 	i->2	
yels	e->6	
yens	 ->1	
yer 	h->1	n->1	
yer.	O->1	
yern	,->1	
yeta	b->1	
yfal	l->1	
yfas	c->1	
yft 	f->2	
yfta	 ->5	d->3	n->2	r->30	s->3	
yfte	 ->15	.->1	n->6	r->2	t->22	
yfto	r->3	
yför	s->1	v->1	
yg d	e->1	
yg f	r->1	å->1	ö->3	
yg i	 ->4	
yg m	e->3	
yg n	ä->1	
yg o	b->1	c->1	m->1	
yg s	o->14	å->1	
yg u	n->2	t->1	
yg),	 ->1	
yg, 	d->1	h->1	s->1	u->1	
yg.E	n->1	
yg.F	ö->1	
yg.V	a->1	i->1	
yg; 	m->1	
yg?D	ä->1	
yga 	a->2	d->1	g->1	i->1	m->1	o->1	s->2	v->1	y->1	
ygad	 ->16	e->5	
ygan	d->6	
ygar	 ->1	
ygbl	a->1	
ygd 	i->1	o->1	
ygd.	D->2	
ygde	n->31	
ygds	b->1	k->1	o->4	r->2	t->1	u->1	
ygel	l->1	s->4	
ygen	 ->3	,->3	s->7	
yger	 ->1	
yget	 ->7	s->1	
ygga	 ->36	d->1	n->23	s->3	
yggd	 ->2	e->2	
ygge	 ->1	l->1	n->3	r->7	t->4	
yggh	e->6	
yggn	a->19	
yggo	r->1	
yggr	a->1	
yggs	 ->2	t->1	
yggt	 ->4	s->1	
ygie	n->2	
ygkr	a->1	
ygni	n->1	
ygpl	a->4	
ygru	p->2	
ygsa	m->4	
ygsb	e->1	
ygsi	n->1	
ygss	k->7	t->1	ä->1	
ygst	a->1	
ygsä	g->1	
ygt 	4->1	e->1	t->1	
ygtr	a->2	
yhet	 ->1	.->2	e->9	s->1	
yhun	 ->1	
yhög	a->1	
yist	e->2	
yk.H	e->1	
yka 	-->1	P->1	a->11	d->5	e->1	f->1	m->1	s->1	u->2	v->1	
yka,	 ->2	
ykas	 ->4	
ykel	 ->1	,->1	.->1	
yker	 ->7	
ykla	r->4	
ykol	o->1	
yks 	o->1	v->1	
ykta	 ->1	d->1	
yktb	a->1	
ykte	 ->4	,->1	.->1	n->3	r->3	
ykti	n->13	
yktr	a->1	
yl g	e->1	
yl o	c->3	
yl, 	f->1	r->1	
yl- 	o->1	
yl.D	e->1	
yl.J	a->1	
yl.V	i->1	
yla.	H->1	
ylan	 ->1	
ylbe	s->1	
yldi	g->29	
ylfö	r->2	
ylib	e->1	
ylig	a->1	e->30	
ylik	a->2	t->1	
ylla	 ->25	.->1	n->3	s->10	
ylld	e->1	
ylle	r->21	
ylln	i->1	
yllr	a->1	
ylls	 ->3	.->1	
yllt	 ->1	,->2	s->1	
ylrä	t->2	
ylsö	k->6	
ym a	t->1	
ym m	e->1	
ym o	m->1	
ym s	o->1	
ym.D	e->1	
yma 	B->1	
ymas	k->1	
ymbo	l->9	
ymd 	t->1	
ymde	n->1	
ymen	 ->1	
ymer	 ->1	
ymit	e->1	
ymma	 ->1	
ymme	 ->10	,->1	r->6	
ympa	d->1	t->8	
ympi	c->1	s->1	
ympn	i->2	
ympt	o->1	
ymra	d->7	r->2	t->1	
yms 	i->1	
ymt 	a->1	
ymts	 ->1	
yn -	 ->1	
yn a	t->1	v->1	
yn g	e->1	
yn h	a->1	
yn i	 ->2	
yn l	y->1	
yn o	c->5	
yn p	å->4	
yn t	i->65	
yn v	a->1	
yn ä	n->1	v->1	
yn å	l->1	
yn, 	m->1	o->1	
yn.A	t->1	
yn.E	t->1	
yn.S	i->1	l->1	
yn; 	d->1	
yna 	h->1	
ynam	i->5	
ynan	d->1	
ynas	 ->1	.->2	
ynaz	i->6	
ynd 	a->1	f->1	g->1	ä->1	
ynda	 ->5	b->2	n->1	r->3	s->3	
ynde	r->1	
yndi	g->164	
yndr	o->1	
ynds	a->4	
ynen	 ->5	.->1	
yner	g->2	
ynes	 ->1	
ynga	n->1	
yngd	 ->2	p->4	
ynge	r->1	
yngr	e->1	
yngs	t->3	
ynli	g->8	
ynn,	 ->1	
ynna	 ->7	d->6	r->5	
ynne	 ->1	!->1	r->52	s->2	
ynns	a->3	
ynon	y->1	
ynpu	n->29	
yns 	s->1	
ynst	a->2	
ynsä	t->4	
ynt 	n->1	v->1	
ynt,	 ->1	
ynte	s->1	
ynvi	n->12	
yo s	k->1	
yola	 ->2	
yon 	1->1	s->1	
yon,	 ->1	
yost	a->1	
yoto	 ->2	-->1	.->1	p->2	s->1	
yp C	a->1	
yp a	v->18	
yp f	å->1	
yp, 	d->1	l->1	
yp.D	e->1	
yp.E	f->1	
ypen	 ->12	
yper	 ->3	n->2	
ypfa	l->1	
ypgo	d->1	
yphå	l->3	
ypla	n->1	
ypot	e->2	
yppa	s->1	
yppe	r->1	
yps.	M->1	
ypte	n->2	
ypto	g->2	
yr a	l->1	
yr e	r->1	
yr f	r->1	
yr h	i->1	
yr j	a->1	
yr.E	f->1	
yra 	a->1	d->3	e->1	f->3	g->1	h->1	i->1	k->2	l->1	m->4	n->1	o->2	p->6	r->1	s->3	u->1	ä->3	å->2	
yra,	 ->1	
yra:	 ->1	
yram	i->1	
yran	d->4	
yrar	 ->5	e->2	
yras	 ->1	.->1	
yrd 	a->1	
yre 	s->1	
yre,	 ->1	
yreg	i->1	
yrek	o->3	
yrel	s->7	
yren	,->1	
yret	 ->1	s->2	
yrie	n->22	r->6	
yrig	h->1	
yris	k->4	
yrka	 ->8	,->1	.->1	n->5	r->1	
yrke	f->1	n->3	p->1	s->15	
yrko	g->1	r->2	
yrne	 ->1	,->1	
yrni	n->7	
yrs 	a->2	
yrt 	o->1	
yrt.	 ->1	
yrti	o->4	
yrå 	s->1	ä->1	
yråe	r->1	
yråk	r->30	
yrån	 ->3	
ys -	 ->1	
ys a	v->16	
ys b	e->3	
ys d	e->1	
ys f	a->1	l->1	ö->1	
ys g	e->1	
ys i	 ->1	
ys j	a->1	
ys o	c->2	r->1	
ys s	o->1	
ys v	i->1	
ys, 	a->1	d->1	u->1	v->1	
ys-d	e->1	
ys.D	e->2	
ys.F	r->1	
ys.G	e->1	
ys.H	ä->1	
ys?D	e->1	
ys?I	 ->1	
ysa 	f->1	m->1	o->2	s->1	u->3	v->1	ä->1	
ysan	d->4	
ysat	o->2	
ysen	 ->5	
yser	 ->7	.->1	a->15	
ysis	k->9	
ysk 	e->1	
yska	 ->21	,->1	p->1	
yskl	a->22	
yskt	 ->2	
ysni	n->5	
yss 	a->1	b->1	e->1	g->1	n->1	o->3	s->2	
yss,	 ->2	
yss.	S->1	
yssa	 ->1	r->1	
ysse	l->122	n->5	
yssl	a->10	
yssn	a->28	i->1	
yst 	f->1	m->4	
yste	m->190	r->2	
ystr	a->1	
yta 	a->1	b->1	d->3	e->1	h->1	k->1	m->4	s->1	
yta.	I->1	
ytan	d->13	
ytas	 ->1	
yte 	a->3	f->2	k->1	m->3	s->1	
yte,	 ->1	
ytel	s->3	
yter	 ->8	i->1	
ytet	 ->6	
ytis	k->1	
ytli	g->2	
ytni	n->3	
yts 	t->1	
ytt 	I->1	a->1	b->2	e->1	f->3	g->1	i->3	k->2	l->1	m->2	o->2	p->5	s->11	t->1	u->1	v->1	å->2	ö->2	
ytt,	 ->3	
ytt.	D->2	J->2	
ytta	 ->20	,->1	.->4	n->1	r->3	s->1	t->1	
ytte	r->91	
ytti	g->13	
yttj	a->41	
yttn	i->4	
ytto	-->1	a->1	
yttr	a->39	e->3	i->1	
ytts	 ->1	
yu i	 ->1	
yu s	a->1	
yval	d->1	
yver	i->1	k->1	
yvär	d->1	r->39	
ywoo	d->1	
yxfi	c->1	
yårs	a->1	
z Fi	s->3	
z Fl	o->2	
z Go	n->1	
z an	g->1	
z be	t->1	
z dy	k->1	
z el	l->1	
z en	 ->1	
z et	t->1	
z fr	å->1	
z få	r->1	
z fö	r->2	
z ha	d->1	
z i 	B->1	
z oc	h->7	k->1	
z om	 ->1	
z sa	d->2	
z so	m->2	
z to	g->2	
z)(T	a->1	
z).H	e->1	
z, G	i->1	
z, L	a->3	
z, b	e->1	
z, i	n->1	
z, p	å->1	
z, t	a->1	
z, u	t->1	
z-ka	t->3	
z. E	u->1	
zFru	 ->1	
za o	c->1	
za, 	d->1	
za.D	e->1	
za.S	i->1	
zaks	t->1	
zare	m->2	
zbek	i->2	
zbet	ä->1	
zen.	J->1	
zes-	C->1	
zida	k->2	
zige	n->4	
zio-	P->4	
zism	 ->2	.->1	e->5	
zist	 ->1	!->1	a->5	e->2	f->1	i->3	
zjik	i->5	
zman	n->2	
zon 	3->1	V->2	o->1	
zone	n->1	r->2	
zoni	n->1	
zore	r->2	
zqui	e->1	
zuel	a->1	
zwal	d->1	
zále	z->1	
º C.	 ->1	
Ämna	r->1	
Än e	n->3	
Ända	 ->1	
Ändr	a->1	i->13	
Ändå	 ->5	
Ännu	 ->3	
Äntl	i->1	
Är I	s->1	
Är d	e->19	
Är h	y->1	
Är i	n->1	
Är k	o->2	
Är r	å->1	
Är s	t->1	
Är v	i->1	
Ärad	e->6	
Även	 ->46	
Å ED	D->1	
Å PS	E->1	
Å an	d->10	
Å en	a->2	
Å ko	m->1	
Å so	c->1	
ÅDSK	A->1	
ÅGOR	N->1	
År 1	9->4	
År 2	0->1	
Året	 ->1	
Årli	g->1	
Åtag	a->1	
Åter	i->1	u->2	v->1	
Åtgä	r->5	
Île-	d->1	
Ö (Ö	s->2	
Ö fö	r->1	
Ö hä	v->1	
Ö in	o->1	
Ö mi	n->1	
Ö oc	h->3	
Ö om	 ->1	
Ö so	m->1	
Ö vi	d->1	
Ö är	 ->1	
Ö) s	i->1	
Ö).J	a->1	
Ö-le	d->1	
Ö-me	d->1	
Ö:s 	a->1	d->1	f->1	s->1	
ÖSTN	I->2	
ÖVP 	(->2	a->2	m->1	
ÖVP)	 ->1	
Ögon	b->2	
Ökad	 ->1	
Öppe	n->1	
Öste	r->81	u->5	
Östt	y->2	
Över	 ->1	v->1	
Övri	g->1	
ález	 ->1	
án, 	a->1	
ánch	e->1	
ão T	o->2	
ä ut	g->1	
ä öv	e->1	
äck 	m->1	o->1	s->1	
äcka	 ->22	,->1	d->1	n->12	s->1	
äcke	n->1	r->37	
äckh	e->1	
äckl	a->1	i->77	
äckn	i->32	
äcko	r->1	
äcks	 ->6	.->1	;->1	c->1	
äckt	 ->9	e->6	s->3	
äckv	i->3	
äd b	e->1	
äd f	ä->1	
äd h	a->2	
äd u	p->1	
äd, 	o->1	
äd.D	e->1	
äda 	E->1	e->1	i->6	s->1	u->2	
äda,	 ->1	
ädan	d->10	
ädar	e->47	n->10	
ädat	 ->1	
ädd 	a->2	f->3	
ädd,	 ->1	
ädda	 ->9	d->3	r->1	t->1	
ädde	 ->7	
äddn	i->4	
äde 	-->1	a->1	e->1	f->1	h->1	i->1	k->1	m->1	o->3	t->4	
äde.	H->1	J->2	
ädeH	e->1	
ädeP	r->1	
ädel	s->6	
äden	 ->3	a->1	
äder	 ->41	,->3	.->1	a->1	i->3	n->8	s->1	
ädes	 ->1	,->1	p->7	v->2	
ädet	 ->10	,->1	.->1	
ädja	 ->6	n->4	r->6	s->1	
ädje	 ->7	
ädre	t->1	
äds 	a->1	d->1	i->1	m->1	r->1	å->2	ö->1	
ädsl	a->9	
äer;	 ->1	
äffa	 ->5	,->2	.->1	d->6	n->41	r->49	s->2	t->9	
äffl	i->2	
äfta	 ->11	,->1	d->3	r->3	s->5	t->7	
äfte	l->1	
äfti	g->1	
äg [	K->1	
äg a	n->1	t->6	v->1	
äg b	o->1	
äg e	l->6	
äg f	ä->1	ö->1	
äg g	e->2	
äg h	i->1	ä->1	
äg i	 ->1	n->1	
äg k	u->1	
äg m	e->1	i->1	o->1	
äg o	c->2	
äg s	i->1	
äg t	r->1	
äg ä	r->1	
äg å	s->1	
äg, 	e->1	f->1	g->1	j->6	o->1	p->1	s->4	v->1	
äg.A	l->1	
äg.B	i->1	
äg.D	e->1	
äg.E	f->1	
äg.J	a->1	
äg.M	e->1	i->1	
äg.O	a->1	
äg.V	a->1	
äg: 	D->1	
ägNä	s->1	
äga 	"->1	-->1	F->1	S->2	a->80	b->2	d->13	e->6	f->5	g->1	h->6	i->5	j->1	k->2	l->3	m->1	n->11	o->9	r->19	s->3	t->8	v->2	ä->2	å->1	
äga,	 ->16	
äga.	D->1	J->1	M->1	
äga:	 ->4	
ägag	å->6	
ägan	d->13	
ägar	 ->7	,->6	.->5	a->1	e->18	n->6	
ägas	 ->4	,->1	
ägby	g->1	
ägd 	g->1	l->1	
ägda	 ->1	
ägde	 ->1	
äge 	d->2	g->1	m->2	s->3	ä->1	
äge,	 ->1	
äge.	H->1	V->1	
ägel	s->8	
ägen	 ->15	,->3	.->1	:->1	h->12	
äger	 ->78	,->4	.->2	:->5	i->36	
äges	b->1	r->2	
äget	 ->16	,->1	.->2	
ägg 	d->1	f->1	g->1	h->2	i->4	k->1	l->1	m->1	s->1	t->4	u->4	v->1	
ägg"	 ->1	
ägg,	 ->1	
ägg.	F->1	
ägga	 ->92	,->1	n->76	s->11	
ägge	n->2	r->39	t->2	
äggi	g->3	
äggn	i->27	
äggs	 ->17	,->1	b->1	f->1	k->1	
ägla	d->4	s->1	
ägle	d->5	
ägli	g->2	
ägmä	r->1	
ägna	 ->16	,->2	r->29	s->2	t->4	
ägne	r->1	
ägni	n->2	
ägra	 ->4	d->4	n->5	r->4	s->1	t->4	
ägre	 ->8	.->2	n->1	
ägrö	j->1	
ägs 	d->2	e->1	g->1	h->1	i->2	
ägse	n->2	t->4	
ägsk	ä->2	
ägsn	a->5	ä->2	
ägso	m->1	
ägst	a->1	
ägt 	d->1	f->1	r->9	
äkar	e->4	k->2	
äkem	e->1	
äken	s->9	
äker	 ->20	,->1	.->1	h->235	l->15	s->24	t->28	
äkna	 ->9	d->1	r->21	s->4	t->5	
äkne	e->1	l->1	
äkni	n->14	
äkra	 ->31	r->4	s->5	
äkri	n->24	
äkt 	f->7	
äkt.	O->1	
äkta	 ->6	d->1	r->5	
äkte	n->3	r->1	t->1	
äkti	g->2	n->1	
äkts	 ->1	a->3	b->1	f->1	
äl -	 ->2	
äl 6	,->1	
äl S	h->1	
äl a	l->1	t->6	v->4	
äl b	e->3	i->1	
äl d	e->6	å->1	
äl e	f->1	k->1	n->2	
äl f	r->1	u->1	ö->9	
äl g	e->2	ä->1	
äl h	a->5	u->1	ä->1	
äl i	 ->6	n->10	
äl k	a->2	u->1	v->1	ä->1	
äl l	ä->1	
äl m	a->1	e->6	o->1	y->1	
äl n	i->1	
äl o	c->3	f->1	
äl p	å->3	
äl r	e->3	
äl s	i->1	k->1	o->12	t->2	
äl t	i->8	
äl u	n->1	p->1	r->3	t->5	
äl v	a->1	e->1	i->1	å->1	
äl ä	n->2	r->3	
äl å	t->1	
äl ö	v->1	
äl, 	i->1	k->1	m->2	o->1	
äl.A	l->1	
äl.D	e->1	
äl.F	r->1	ö->2	
äl.J	a->2	
äl.M	i->1	
äl.S	a->1	
äla 	d->1	v->1	
älan	 ->1	
älbe	s->1	
äld 	å->1	
älda	 ->1	
äldi	g->23	
äldr	e->7	
älen	 ->3	"->1	.->1	
äler	.->1	i->1	
älet	 ->8	,->1	
älft	e->3	
älfu	n->1	
älfä	r->8	
älgr	u->2	
älgö	r->1	
älha	v->1	
älig	 ->1	
älja	 ->8	r->13	s->1	
älje	r->5	
äljn	i->3	
älkl	i->1	
älko	m->50	
älkä	n->3	
äll 	u->1	ä->1	
äll,	 ->2	
äll.	J->1	O->1	
äll?	K->1	
älla	 ->94	,->1	.->2	:->1	n->54	r->6	s->20	
ällb	a->1	
älld	 ->5	a->23	e->29	h->23	
älle	 ->36	,->1	.->1	l->7	n->64	r->405	s->2	t->88	
älli	g->56	
älln	i->71	
ällo	r->39	
älls	 ->18	.->2	e->3	k->8	m->1	o->1	s->1	v->1	y->2	
ällt	 ->15	,->1	.->1	s->9	
älme	n->2	
älmå	e->2	
älni	n->12	
älp 	a->27	d->1	f->6	n->1	o->2	p->1	s->2	t->5	v->2	ö->1	
älp,	 ->2	
älp.	D->1	H->1	I->1	J->1	V->1	
älpa	 ->37	n->3	r->1	
älpe	n->4	r->1	
älpl	i->1	
älps	.->1	
älpt	 ->1	a->1	e->1	
älpv	i->1	
äls 	m->1	t->1	
älsa	 ->15	,->3	.->1	n->4	r->1	
älsi	g->1	
älsk	a->2	
älsn	i->2	
älso	-->1	e->1	r->2	s->1	v->3	
älst	r->1	å->6	
ält 	a->1	e->1	i->1	o->1	p->1	s->1	
älta	l->2	
älte	 ->2	,->2	n->2	t->9	
ältn	i->1	
älts	i->1	
älut	b->1	v->2	
älv 	a->5	b->2	f->5	g->1	h->3	i->3	k->1	m->1	o->3	s->7	t->1	u->2	v->2	ä->3	
älv,	 ->5	
älv.	D->1	J->1	K->1	V->1	
älva	 ->61	,->3	.->5	n->1	
älvb	e->3	i->1	ä->1	
älvf	a->2	ö->1	
älvh	j->1	
älvk	l->20	o->1	
älvn	i->3	
älvp	l->1	
älvs	t->15	ä->1	
älvt	 ->5	
älvä	n->1	
ämbe	t->8	
ämd 	a->1	h->1	i->1	o->1	t->1	v->1	
ämda	 ->8	,->1	
ämde	 ->5	
ämdh	e->1	
ämel	s->1	
ämfö	r->18	
ämja	 ->36	.->1	n->17	r->6	s->1	t->1	
ämka	 ->1	r->1	
ämli	g->62	k->13	n->34	
ämma	 ->18	,->1	d->3	n->10	r->1	s->3	
ämme	l->122	r->39	
ämmi	g->4	
ämn 	s->1	
ämn,	 ->1	
ämn.	D->1	
ämna	 ->54	,->1	d->9	n->3	r->23	s->13	t->18	
ämnd	a->8	e->18	
ämne	 ->3	.->2	:->1	n->19	r->5	t->4	
ämni	n->17	
ämns	 ->8	.->1	
ämnt	 ->9	,->2	.->2	s->6	
ämnv	i->1	ä->1	
ämpa	 ->69	d->1	n->3	r->13	s->42	t->8	
ämpe	l->1	
ämpl	i->61	
ämpn	i->80	
ämra	 ->2	d->4	n->1	r->1	s->2	
ämre	 ->5	
äms 	u->1	
ämsi	d->1	
ämst	 ->39	.->1	a->13	ä->24	
ämt 	a->4	e->1	f->2	i->1	o->1	p->1	s->4	t->1	ö->2	
ämt,	 ->3	
ämt.	D->1	
ämta	 ->3	n->1	r->1	s->1	t->1	
ämtn	i->1	
ämts	a->1	
ämvi	k->2	
än 1	 ->2	0->3	6->1	
än 2	0->1	1->1	
än 3	0->2	
än E	u->1	
än F	o->1	
än W	a->1	
än a	c->1	l->2	t->13	v->1	
än b	a->2	
än d	e->20	i->2	
än e	j->1	l->1	n->30	t->4	
än f	a->2	e->3	r->1	ö->7	
än g	e->2	i->2	
än h	a->3	i->1	
än i	 ->14	n->3	
än j	a->1	
än k	a->2	o->4	
än l	i->1	o->1	ä->2	
än m	a->5	e->2	i->5	y->1	å->1	
än n	a->1	ä->2	å->6	
än o	c->13	m->3	
än p	.->1	e->1	o->1	å->4	
än r	a->2	e->4	
än s	a->1	k->2	o->10	t->3	ä->1	å->6	
än t	i->7	r->2	v->2	
än u	t->2	
än v	a->7	i->7	ä->3	å->1	
än ä	r->4	
än å	k->6	r->2	
än, 	e->1	m->1	
än.I	n->1	
än.J	a->2	
än.T	y->1	
än; 	d->1	
äna 	a->1	n->1	r->1	s->4	
änad	e->1	
änar	 ->14	.->2	
änd 	(->1	b->3	e->1	m->4	
änd,	 ->2	
änd.	K->1	
ända	 ->88	,->1	.->5	?->1	m->13	n->8	r->9	s->16	t->1	
ändb	a->9	
ände	 ->26	,->1	.->1	b->9	l->27	r->249	s->11	t->1	
ändi	g->232	
ändl	i->5	ö->1	
ändn	i->64	
ändp	u->6	
ändr	a->75	i->293	
änds	 ->20	k->26	
ändå	 ->51	,->1	.->1	
änfö	r->1	
äng 	g->1	k->2	o->1	å->1	
äng.	D->1	
änga	 ->13	,->1	n->3	r->6	s->4	
ängb	r->1	
ängd	 ->17	a->1	e->12	
änge	 ->35	l->1	r->18	s->1	t->1	
ängi	g->2	l->1	
ängl	i->23	
ängn	i->44	
ängr	e->62	
ängs	 ->2	l->1	y->2	
ängt	 ->6	a->1	e->8	
änhe	t->47	
änie	n->1	
änin	g->1	
änit	e->12	
änk 	b->1	p->1	t->1	
änka	 ->37	,->1	n->288	s->3	
änkb	a->4	
änke	n->1	r->41	
änkl	i->5	
änkn	i->15	
änks	 ->3	a->2	
änkt	 ->5	.->1	a->8	e->3	s->3	
änli	g->15	
änna	 ->69	,->1	.->2	g->9	n->26	s->8	
änne	 ->1	d->1	l->1	n->28	r->74	t->6	
änni	n->10	s->98	
änns	 ->3	.->1	
ännu	 ->72	.->4	;->1	
änny	t->2	
äns 	f->1	p->1	s->2	v->2	
änsa	 ->12	,->1	d->27	n->3	r->5	s->5	t->9	
änsc	h->2	
änse	e->8	n->4	r->30	
änsf	r->2	
änsk	a->1	l->42	o->7	
änsl	a->15	e->7	i->21	o->7	
änsn	i->12	
änso	m->1	
änsp	r->1	
änst	 ->6	,->1	.->2	e->124	f->1	g->3	r->1	
änsv	ä->1	
änsy	n->72	
änsö	v->12	
änt 	-->1	a->8	d->3	e->4	f->2	g->1	h->1	i->3	k->1	l->1	m->5	o->1	p->2	s->9	t->3	u->5	
änt,	 ->3	
änt.	J->1	V->1	
änt:	 ->1	
änta	 ->43	.->2	d->1	n->5	r->39	s->2	t->5	
äntl	i->20	
äntn	i->7	
änts	 ->13	
änvi	s->35	
äpad	e->1	
äpna	d->2	
äpni	n->1	
äpp 	a->1	k->1	
äpp,	 ->1	
äpp.	D->1	
äppa	 ->7	n->2	
äppe	n->3	r->2	t->1	
äpph	ä->1	
äpps	r->1	
äppt	e->3	
äpro	d->1	
är "	k->1	
är -	 ->13	
är 1	,->1	/->1	0->2	6->1	
är 2	5->1	9->1	
är 3	0->1	
är 5	0->1	
är 7	 ->1	
är 8	0->1	
är A	n->1	
är B	a->8	o->1	
är C	E->1	
är D	o->1	
är E	U->5	g->1	u->11	
är F	N->1	P->1	
är K	i->5	
är L	u->1	
är M	a->1	o->13	
är N	i->1	
är P	a->17	o->2	r->1	
är R	e->2	
är S	c->1	o->1	
är V	i->4	
är W	a->2	
är a	b->10	c->2	k->5	l->45	m->1	n->40	r->4	t->167	v->40	
är b	a->14	e->81	l->3	o->3	r->22	u->1	y->1	ä->7	å->5	ö->3	
är c	e->2	i->1	o->1	
är d	a->7	e->579	i->6	j->4	o->18	r->2	ä->29	å->5	ö->1	
är e	f->4	g->6	k->1	l->1	m->12	n->243	r->1	t->123	u->1	v->1	x->6	
är f	a->30	e->7	i->10	l->4	o->16	r->46	u->11	y->1	ä->1	å->1	ö->100	
är g	a->7	e->11	i->2	j->2	l->13	o->8	r->7	å->5	
är h	a->35	e->32	i->2	j->1	o->5	u->6	ä->4	å->2	ö->1	
är i	 ->89	b->2	d->2	l->1	n->156	s->1	
är j	a->51	u->18	ä->1	
är k	a->13	l->14	n->5	o->58	r->3	u->1	v->2	ä->7	
är l	a->6	e->6	i->21	o->2	y->2	ä->16	å->6	ö->4	
är m	a->48	e->50	i->15	o->4	u->1	y->56	ä->2	å->10	ö->21	
är n	a->18	e->5	i->8	o->2	u->11	y->6	ä->13	å->29	ö->34	
är o	a->5	b->4	c->55	e->8	f->10	j->1	k->2	l->4	m->15	n->1	r->6	s->2	t->3	u->3	
är p	a->7	e->3	l->6	o->10	r->22	u->2	å->18	
är r	e->28	i->12	o->2	u->3	ä->13	å->2	ö->1	
är s	a->16	e->4	i->5	j->9	k->20	l->3	n->3	o->17	p->6	t->23	u->2	v->11	y->7	ä->46	å->27	
är t	a->2	e->5	i->40	j->2	o->2	r->6	v->10	y->21	ä->3	
är u	n->10	p->23	r->1	t->26	
är v	a->13	e->17	i->161	u->1	ä->32	å->10	
är y	p->1	r->1	t->10	
är Ö	s->1	
är ä	g->1	l->2	n->12	r->15	v->4	
är å	r->2	t->3	
är ö	d->1	k->1	n->2	p->3	v->30	
är! 	1->1	B->1	C->1	D->2	E->3	F->1	I->2	J->6	L->2	N->2	O->1	T->1	U->1	V->4	Ä->1	
är!.	H->1	
är!D	e->1	
är!E	r->1	
är!J	a->1	
är, 	a->13	b->3	d->3	f->9	h->6	i->4	j->3	k->14	l->1	m->15	n->4	o->9	p->1	r->1	s->5	t->3	u->2	v->9	ä->10	
är. 	D->1	N->1	i->1	
är..	 ->1	
är.D	e->9	ä->1	
är.E	f->1	n->1	
är.F	ö->4	
är.G	e->1	
är.H	e->1	
är.I	 ->1	
är.J	a->11	
är.K	o->1	
är.R	a->1	
är.S	o->2	å->1	
är.V	a->1	i->7	
är.k	o->1	
är: 	F->1	h->1	n->1	v->1	Ä->1	
är; 	v->1	
är?D	e->1	
är?H	a->1	
är?J	a->1	
ära 	5->1	a->14	b->2	d->3	e->5	f->11	h->5	i->1	k->59	l->2	m->4	o->7	p->3	r->1	s->13	u->5	ä->2	å->1	
ära,	 ->2	
ära.	N->1	
ärad	e->22	
äran	 ->18	,->3	.->3	?->1	d->3	
ärar	e->2	t->1	
äras	 ->6	
ärav	 ->4	
ärbe	s->1	
ärd 	2->1	a->4	b->1	d->2	e->3	f->2	k->1	m->3	o->4	s->3	u->1	v->2	
ärd,	 ->8	
ärd.	D->3	H->1	I->1	J->1	
ärd;	 ->2	
ärda	 ->23	,->2	.->1	n->5	r->2	s->2	t->2	
ärde	 ->18	,->1	-->1	.->4	d->2	f->7	g->3	l->1	n->20	r->268	s->2	t->4	
ärdi	g->41	
ärdl	i->3	
ärdo	m->7	
ärds	 ->1	b->1	l->1	m->1	o->1	p->7	s->3	v->1	
äre 	k->1	
äref	t->12	
ärem	o->19	
ären	 ->41	,->6	.->2	?->1	d->21	s->3	
ärer	 ->14	!->1	,->5	.->1	n->14	
äret	 ->1	
ärfr	å->1	
ärfö	r->280	
ärg,	 ->2	
ärga	d->1	
ärhe	t->5	
ärhä	n->1	
äri 	s->1	v->1	
ärib	l->6	
ärif	r->2	
ärig	e->19	
ärin	g->12	
ärja	d->2	
ärka	 ->26	,->1	n->2	s->3	
ärkb	a->3	
ärke	 ->7	l->5	n->2	r->7	t->1	
ärki	l->1	
ärkl	i->5	
ärkn	i->19	
ärks	 ->3	.->3	a->53	
ärkt	 ->21	.->1	a->18	s->1	
ärl 	o->1	
ärld	 ->1	,->2	.->1	e->37	s->17	
ärle	d->1	k->2	
ärli	g->20	n->1	
ärma	 ->2	n->1	r->20	s->13	
ärme	d->49	l->1	
ärmi	n->10	
ärmn	i->5	
ärn-	 ->2	
ärna	 ->34	.->1	n->6	r->1	
ärne	n->8	
ärnf	r->2	
ärni	n->4	
ärnk	a->1	r->22	
ärnp	r->2	u->2	
ärns	t->1	ä->3	
ärnt	e->3	
ärnv	a->8	ä->15	
äro 	t->1	
äroa	n->1	
ärom	 ->1	
äros	a->1	
ärpa	 ->6	s->2	
ärpe	r->1	
ärpl	a->1	
ärpn	i->1	
ärpo	l->2	
ärpt	a->2	
ärpå	 ->2	
ärr 	a->1	b->3	d->3	f->3	g->1	h->6	i->4	k->3	n->1	o->2	s->4	ä->5	å->1	
ärr,	 ->2	
ärr.	V->1	
ärra	 ->1	r->2	s->2	t->1	
ärre	 ->8	,->1	
ärrä	t->1	
ärrö	r->4	
ärs 	f->2	h->1	m->1	n->1	s->1	
ärsk	i->158	t->1	
ärsm	ä->1	
ärst	 ->1	a->7	
ärsy	n->1	
ärt 	F->1	a->12	b->1	e->5	f->1	g->1	i->1	k->1	m->2	o->3	p->1	s->2	
ärt,	 ->5	
ärt.	J->1	O->1	S->1	V->1	
ärta	 ->3	d->1	n->2	r->1	t->14	
ärti	l->2	
ärtl	i->7	
ärto	m->17	
ärts	a->1	
ärut	ö->1	
ärv 	o->1	
ärva	 ->6	d->1	r->47	t->1	
ärvb	r->1	
ärvh	e->1	
ärvi	d->6	
ärvl	i->1	
ärvs	a->3	
ärvt	 ->2	
äs t	e->1	
äs u	n->1	
äs y	t->1	
äsa 	k->1	o->1	v->1	
äsba	r->2	
äsch	 ->1	e->1	
äsdu	k->1	
äsen	 ->2	,->2	d->6	t->26	
äser	 ->6	
äsfr	ä->1	
äsk.	H->1	
äsku	n->1	
äsni	n->2	
äson	g->1	
ässi	g->31	
äst 	D->1	a->1	d->2	e->2	f->1	g->1	k->1	r->1	s->1	t->1	
ästa	 ->97	.->4	n->19	r->2	
ästb	a->4	
äste	 ->3	l->1	n->1	r->8	s->1	
ästk	u->1	
ästm	a->1	
ästn	i->2	
ästr	a->3	
ästs	 ->1	
ästv	ä->1	
ät d	ä->1	
ät k	a->1	
ät m	i->1	
ät o	c->1	s->1	
ät s	i->1	k->2	o->2	
ät. 	D->1	
äta 	d->1	s->1	
äta,	 ->1	
ätar	e->2	
ätas	 ->2	
äte.	O->1	
äten	 ->4	
äter	 ->2	
ätet	 ->2	
äthe	t->1	
ätig	t->1	
ätor	 ->1	
ätsk	a->1	
ätst	r->1	
ätt 	(->2	-->2	H->1	a->55	b->9	e->7	f->18	g->7	h->8	i->18	k->23	l->3	m->5	n->4	o->24	p->9	r->6	s->47	t->22	u->8	v->11	ä->10	å->2	ö->2	
ätt,	 ->37	
ätt.	 ->2	A->2	B->1	D->13	E->3	F->2	H->6	I->1	J->7	K->2	L->1	M->5	N->2	S->4	V->5	Ä->1	
ätt:	 ->2	
ätt?	A->1	D->1	O->1	S->1	
ätta	 ->167	!->1	,->4	.->3	d->9	n->24	r->24	s->24	t->10	
ätte	 ->20	,->1	d->1	g->1	l->4	n->85	r->66	s->1	t->23	
ättf	r->1	ä->7	ö->1	
ätth	å->9	
ätti	g->122	l->2	
ättl	i->1	
ättm	ä->1	
ättn	a->1	i->213	
ättr	a->60	e->75	i->18	
ätts	 ->11	,->2	.->1	a->4	f->1	h->2	i->2	k->9	l->118	o->6	p->2	r->1	s->53	t->4	v->4	
ättv	i->74	
ättä	n->1	
ätve	r->11	
äv m	e->1	
äva 	4->1	a->8	d->4	e->9	f->3	i->2	j->1	k->1	m->2	s->1	t->3	å->2	ö->1	
ävad	e->4	
ävan	 ->8	.->1	d->7	s->1	
ävar	 ->4	e->1	
ävas	 ->11	,->1	.->1	
ävat	 ->1	
ävda	 ->7	d->3	r->12	t->5	
ävde	 ->1	,->1	s->2	
ävdv	u->1	
även	 ->266	t->9	
äver	 ->44	.->2	
äves	 ->1	
ävig	t->1	
ävja	s->1	
ävla	d->1	r->1	
ävli	n->1	
ävna	d->4	
ävni	n->10	
ävs 	a->2	b->1	d->11	e->12	f->8	h->1	i->2	k->1	m->2	o->1	p->1	r->1	s->4	u->1	v->3	ä->1	
ävs,	 ->3	
ävs.	E->2	
ävt 	e->1	s->1	
ävts	 ->1	.->1	
ävul	e->1	s->1	
äxa 	u->1	
äxa.	H->1	M->1	
äxan	?->1	d->6	
äxat	 ->1	
äxel	k->1	v->2	
äxer	 ->6	,->1	
äxla	n->1	r->1	
äxli	n->2	
äxor	.->1	
äxt 	a->1	o->4	s->1	ä->1	
äxt,	 ->2	
äxt.	K->1	O->1	
äxtb	r->1	
äxte	n->8	r->2	
äxth	u->7	
äxts	k->3	
å "m	e->1	
å - 	a->1	d->1	i->1	m->1	o->3	s->1	
å 10	 ->1	0->1	
å 13	 ->2	
å 14	0->1	
å 19	9->1	
å 20	 ->1	0->2	
å 22	,->1	
å 24	 ->1	
å 33	 ->1	
å 34	 ->1	
å 37	 ->1	
å 40	 ->1	
å 5 	m->1	
å 50	 ->1	-->1	
å 7,	2->1	
å 75	 ->1	
å 80	 ->2	
å 86	 ->1	
å 90	 ->1	
å 95	 ->1	
å Al	l->2	
å As	s->1	
å At	l->1	
å BS	E->1	
å Ba	l->5	
å Be	l->1	
å CE	N->1	
å CS	U->1	
å Da	 ->1	
å EG	-->4	
å EU	-->2	:->2	
å Er	i->2	
å Eu	r->18	
å Fl	a->1	
å Fö	r->1	
å Ge	n->1	
å Go	l->2	
å Ho	l->1	
å IS	P->1	
å In	t->6	
å Ir	l->1	
å Is	r->1	
å Ki	n->1	
å Ma	l->1	
å Mo	r->1	
å Ol	i->1	
å PP	E->1	
å Pa	p->1	
å Ri	c->2	
å Ro	i->1	
å Ty	s->1	
å Vä	s->2	
å ab	s->1	
å ac	c->1	
å ak	t->4	
å al	b->1	l->40	t->1	
å am	b->1	
å an	 ->1	d->22	g->1	l->1	m->1	n->1	s->10	t->3	v->1	
å ar	b->9	g->1	t->5	
å as	p->2	y->1	
å at	t->353	
å av	 ->18	f->1	g->4	s->2	t->1	
å ba	l->2	r->6	s->3	
å be	 ->1	f->4	g->1	h->10	k->4	r->4	s->5	t->9	
å bi	d->1	l->6	
å bl	e->1	i->8	o->1	y->1	
å bo	l->1	r->8	s->1	
å br	a->3	e->5	i->1	o->3	
å by	g->2	
å bä	r->3	s->8	t->2	
å bå	d->3	
å bö	r->10	
å ce	n->1	
å ci	v->1	
å cr	i->1	
å da	g->9	n->1	
å de	 ->69	b->2	f->2	l->6	m->9	n->124	r->4	s->16	t->166	
å di	r->2	s->2	
å dj	u->7	
å do	m->2	
å dr	a->1	u->1	
å du	b->3	m->1	
å dy	l->1	
å dä	r->3	
å då	l->1	
å ef	f->5	t->2	
å eg	e->3	
å ek	o->6	
å el	e->1	l->3	
å em	b->1	
å en	 ->130	a->12	d->1	g->1	h->3	i->1	k->1	l->2	o->1	s->1	
å er	 ->3	,->1	a->1	k->1	s->1	t->1	
å et	a->1	t->172	
å eu	r->14	
å ex	a->1	e->2	
å fa	k->2	l->4	m->2	r->4	s->9	
å fe	l->1	m->2	n->1	
å fi	n->12	s->2	
å fl	e->3	y->2	
å fo	k->1	l->2	r->5	
å fr	a->22	e->2	i->2	å->30	
å fu	l->2	n->1	
å fy	r->2	
å fä	l->5	r->1	
å få	 ->3	r->7	t->2	
å fö	l->5	r->129	t->2	
å ga	r->2	t->1	
å ge	 ->2	m->16	n->8	o->1	r->1	
å gi	v->1	
å gl	a->1	o->1	
å go	d->3	t->1	
å gr	a->3	u->83	ä->1	
å gä	l->2	r->2	
å gå	 ->1	n->5	r->3	
å gö	r->7	
å ha	 ->5	d->2	n->5	r->11	t->1	v->5	
å he	l->9	m->3	t->2	
å hi	n->1	
å hj	ä->6	
å ho	m->1	p->1	s->1	t->1	
å hu	r->19	v->1	
å hä	n->2	r->5	v->1	
å hå	l->1	
å hö	g->3	
å i 	A->1	S->1	T->1	b->1	c->1	d->11	e->9	f->5	g->1	k->4	l->2	n->1	p->1	r->1	s->7	v->3	
å ia	k->1	
å ic	k->1	
å id	é->1	
å ig	e->4	å->1	
å ih	o->1	
å il	l->2	
å im	p->1	
å in	 ->15	f->5	g->4	i->1	l->2	n->6	o->1	r->5	s->9	t->29	v->3	
å ir	l->1	
å it	a->1	
å ja	g->7	k->1	
å jo	r->2	
å ju	 ->1	s->2	
å jä	r->3	
å ka	d->1	l->11	m->2	n->26	t->2	
å kl	a->7	i->1	
å kn	u->1	
å ko	l->5	m->43	n->24	r->10	
å kr	a->2	i->4	ä->1	
å ku	n->3	
å kv	a->3	i->2	
å kä	n->1	r->2	
å kö	r->2	
å la	g->4	n->13	
å li	g->1	k->3	s->3	t->3	
å lo	b->1	k->2	s->1	v->1	
å ly	c->1	
å lä	g->2	m->4	n->25	s->1	t->2	
å lå	g->5	n->18	t->1	
å lö	r->1	
å ma	j->1	n->3	r->13	s->1	
å me	d->41	l->3	n->3	r->6	
å mi	g->2	l->13	n->21	s->1	t->1	
å mo	d->2	n->1	t->4	
å my	c->43	
å mä	n->2	
å må	l->3	n->24	s->17	t->2	
å mö	j->10	
å na	t->4	
å ne	d->2	
å no	g->1	r->3	t->3	
å ny	 ->2	a->4	c->1	s->1	t->21	
å nä	m->2	r->8	s->4	t->1	
å nå	g->31	t->1	
å nö	d->4	
å oa	c->2	
å ob	e->2	l->1	
å oc	h->48	k->7	
å oe	n->1	
å of	f->1	t->5	
å og	y->1	
å ol	i->3	j->3	
å om	 ->15	f->1	k->1	r->16	t->1	
å on	s->2	
å or	d->4	g->1	s->1	
å os	s->7	
å pa	p->1	r->4	s->2	
å pe	n->2	r->5	s->1	
å pl	a->11	
å po	l->2	s->2	ä->1	
å pr	e->1	i->8	o->7	
å pu	n->9	
å på	 ->16	m->3	p->2	t->1	v->1	
å ra	n->1	s->1	t->1	
å re	a->1	d->4	f->2	g->16	k->1	s->12	
å ri	k->4	s->2	
å ry	g->2	
å rä	c->2	d->1	k->2	t->12	
å rå	d->10	
å rö	d->1	s->2	
å sa	d->1	k->5	m->31	n->2	t->1	
å se	 ->13	d->1	k->3	m->1	n->8	r->2	s->1	
å si	f->1	g->8	k->7	n->17	s->1	t->5	
å sj	ä->3	
å sk	a->17	e->3	i->1	o->2	u->11	y->1	ä->2	
å sl	u->2	å->1	
å sm	i->1	å->7	
å sn	a->31	
å so	c->2	m->38	
å sp	e->10	r->1	å->1	
å st	a->13	e->2	o->13	r->8	u->2	ä->2	ö->9	
å su	b->2	
å sv	a->1	å->4	
å sy	d->1	f->1	s->3	
å sä	g->15	k->7	r->2	t->17	
å så	 ->26	d->3	v->2	
å ta	 ->12	c->7	l->13	n->1	r->1	s->2	
å te	k->1	m->1	r->1	x->1	
å ti	d->7	l->57	m->3	
å tj	ä->1	
å to	g->1	p->1	r->9	
å tr	a->4	e->6	o->4	ö->3	
å tv	i->1	ä->1	å->6	
å ty	c->1	d->1	s->1	
å tä	n->3	
å un	d->10	g->1	i->6	
å up	p->21	
å ut	 ->6	,->1	a->3	f->2	g->2	o->2	r->1	s->2	t->1	v->3	ö->1	
å va	d->12	k->1	l->2	n->1	r->27	t->1	
å ve	c->1	d->4	m->2	r->5	t->11	
å vi	 ->11	a->1	c->1	d->15	k->18	l->31	s->11	t->1	
å vr	e->1	
å vä	g->29	l->4	r->3	s->2	
å vå	r->26	
å yt	t->3	
å zi	g->2	
å Ös	t->2	
å äg	n->1	
å än	 ->2	d->7	n->2	t->1	
å är	 ->44	
å äv	e->3	
å åh	ö->1	
å år	 ->6	,->1	s->1	
å ås	i->1	
å åt	 ->1	a->1	e->4	g->4	m->2	
å ök	a->2	
å ön	 ->1	s->1	
å öp	p->6	
å öv	e->6	
å, a	l->1	t->3	
å, b	ö->2	
å, d	ä->1	
å, e	l->1	n->1	t->1	
å, f	r->3	ö->4	
å, g	e->1	
å, h	e->2	u->1	
å, i	 ->2	
å, l	ö->1	
å, m	e->7	
å, n	u->1	ä->3	
å, o	b->1	c->8	f->1	m->3	
å, r	i->1	ä->1	ö->1	
å, s	o->1	t->1	å->2	
å, t	i->1	
å, v	i->1	å->1	
å, ä	r->1	
å. D	e->2	
å...	.->1	
å.At	t->2	
å.Be	t->1	
å.Bi	s->1	
å.Br	i->1	
å.De	 ->1	n->2	t->10	
å.Do	c->1	
å.Dä	r->2	
å.En	 ->1	
å.Eu	r->2	
å.FP	Ö->1	
å.Fr	u->1	
å.Fö	r->2	
å.Ge	n->1	
å.Gr	a->1	
å.He	r->2	
å.I 	s->1	
å.In	t->1	
å.Ja	g->8	
å.Ju	s->1	
å.Jä	m->1	
å.Me	n->1	
å.Ni	 ->1	
å.No	r->1	
å.Nä	r->2	
å.Oc	h->1	
å.Om	 ->1	
å.Or	d->1	
å.På	 ->2	
å.Sl	u->1	
å.So	c->1	
å.Un	i->1	
å.Vi	 ->4	
å.Är	 ->2	
å: a	t->1	
å: d	e->2	
å: f	ö->2	
å: Ö	p->1	
å: å	 ->1	
å; d	e->1	
å?. 	(->1	
å?In	t->1	
å?Ja	g->1	
å?Se	r->1	
åbar	 ->2	
åber	o->1	
åbju	d->1	
åbör	j->11	
åd (	a->1	
åd -	 ->1	
åd a	n->1	t->1	
åd b	e->1	
åd f	r->2	ö->1	
åd i	 ->1	
åd n	ä->1	
åd o	c->2	m->3	
åd s	o->3	
åd, 	b->1	m->1	o->2	
åd.D	e->1	
åd.J	a->1	
åd.K	a->1	
åd.L	å->1	
åd.M	e->1	
åd?Ä	r->1	
åda 	a->1	b->3	d->6	e->5	f->7	g->1	h->1	i->1	l->2	m->3	n->1	o->3	p->2	s->3	
åda,	 ->1	
ådad	 ->1	e->2	
ådan	 ->57	,->2	.->2	?->1	a->49	d->5	t->54	
ådar	 ->1	.->1	e->1	n->1	
ådd 	m->1	
ådda	 ->4	
ådde	 ->3	s->1	
åde 	-->1	D->1	S->2	a->5	b->2	d->10	e->4	f->9	g->1	h->4	i->9	k->4	m->14	n->2	o->7	p->4	r->2	s->10	t->1	v->4	ä->5	å->1	ö->1	
åde,	 ->14	
åde.	 ->1	D->4	F->4	I->2	J->3	M->4	O->2	P->1	T->1	V->1	
åde:	 ->1	
åde;	 ->1	
åde?	D->1	
ådef	ö->1	
åden	 ->61	)->1	,->10	.->20	:->2	;->1	?->2	a->36	s->1	
åder	 ->26	)->7	a->3	
ådet	 ->212	)->1	,->47	.->52	:->1	?->4	s->99	
ådfr	å->6	
ådgi	v->26	
ådgö	r->1	
ådli	g->7	
ådni	n->1	
ådra	g->1	
ådsb	e->1	
ådsk	a->20	
ådsl	a->3	
ådsm	e->1	i->1	ö->1	
ådso	r->20	
ådsr	ä->1	
ådst	o->1	
åeli	g->6	
åels	e->8	
åend	e->136	
åer 	g->1	i->3	o->1	s->1	
åer,	 ->3	
åer.	D->2	K->1	M->1	
åer:	 ->1	
åern	a->1	
ået.	D->1	
åfre	s->1	
åföl	j->4	
åför	e->6	
åg I	r->1	
åg a	r->1	t->15	v->2	
åg d	e->5	ä->1	
åg e	l->1	t->1	
åg h	ö->1	
åg i	n->2	
åg n	i->2	å->1	
åg o	m->1	
åg r	e->1	
åg s	i->2	o->1	
åg t	i->1	
åg u	t->2	
åg Ö	s->1	
åg ä	r->1	
åg, 	v->1	
åg.E	u->1	
åga 	-->1	a->18	b->3	e->2	f->7	g->6	h->9	i->9	j->1	k->8	m->7	n->27	o->83	p->3	r->4	s->47	t->5	v->6	ä->9	ö->1	
åga!	F->1	
åga,	 ->26	
åga.	 ->1	-->1	A->1	D->8	E->2	F->2	H->3	I->2	J->8	M->2	N->1	O->2	S->1	T->1	U->1	V->5	Ä->1	
åga:	 ->7	
åga?	.->1	
ågad	e->8	
ågan	 ->173	,->14	.->16	:->5	;->1	?->1	d->1	
ågar	 ->24	.->1	
ågas	a->1	ä->19	
ågat	 ->3	,->1	a->1	s->2	
ågav	a->1	
ågek	o->1	
ågel	l->1	s->1	v->1	
ågen	 ->1	
åger	i->1	p->1	
åges	t->10	
åget	 ->1	e->2	
ågic	k->3	
ågkr	a->2	
ågla	r->6	
åglä	n->1	
ågni	n->8	
ågol	y->1	
ågon	 ->110	,->2	.->1	s->15	t->39	
ågor	 ->177	)->1	,->37	.->28	:->4	;->1	?->1	l->1	n->28	
ågot	 ->184	,->2	.->6	?->1	
ågra	 ->149	
ågru	p->3	
ågrä	l->1	
ågs 	i->1	m->1	
ågs.	J->1	L->1	
ågt 	s->1	v->1	
ågve	r->1	
ågå 	i->1	
ågåe	n->6	
ågår	 ->7	.->3	
ågåt	t->1	
åhun	d->1	
åhän	d->6	
åhär	.->1	
åhör	a->1	
åja,	 ->1	
åk f	ö->1	
åk p	å->3	
åk t	i->1	
åk. 	D->1	
åka 	e->1	
åkar	 ->5	e->3	n->1	
åket	 ->2	.->2	
åkig	t->3	
åkla	g->37	
åkli	g->3	
åkom	r->2	
åkra	t->30	
åkta	g->1	
åkte	 ->1	
ål (	B->1	
ål 1	 ->2	,->2	-->11	.->1	
ål 2	 ->5	,->1	-->3	.->1	
ål 5	b->2	
ål a	t->3	v->1	
ål b	e->2	
ål e	n->1	
ål f	i->1	ö->19	
ål g	å->1	
ål h	e->1	i->1	
ål i	 ->7	
ål j	a->1	
ål l	i->1	
ål n	å->1	
ål o	c->5	m->3	
ål p	å->2	
ål r	ö->1	
ål s	k->1	o->13	ä->1	
ål t	i->1	
ål u	p->2	
ål ä	r->4	
ål, 	R->1	f->2	g->1	h->1	m->2	n->1	o->1	p->1	s->6	u->1	
ål-2	-->1	
ål.B	ä->1	
ål.D	e->2	ä->1	
ål.E	t->1	
ål.F	r->1	
ål.H	e->2	
ål.I	 ->2	
ål.J	a->1	
ål.K	u->1	
ål.M	a->1	e->1	
ål.N	ä->2	
ål.Ä	v->1	
ål: 	V->1	a->1	
åla 	b->1	f->1	
åla,	 ->1	
ålag	d->1	o->1	t->2	
ålam	o->2	
ålar	e->2	f->1	
åld 	i->1	o->1	
ålde	r->12	t->2	
åldr	a->3	
ålds	a->3	h->2	u->1	
åldt	a->2	
åled	e->44	
ålen	 ->15	.->2	s->1	
ålet	 ->23	,->2	.->5	
ålfö	r->5	
ålge	m->1	
ålig	 ->5	a->8	g->5	h->1	t->8	
ålin	d->25	r->4	
ålit	l->1	
ålka	s->1	
åll 	a->1	f->2	h->1	i->3	k->2	o->3	r->1	s->4	t->1	v->1	
åll,	 ->5	
åll.	D->2	F->1	I->1	J->2	V->1	
åll:	 ->1	
åll?	.->1	
ålla	 ->85	,->1	n->84	r->1	s->11	
ållb	a->25	
ålle	n->1	r->94	t->27	
ålli	t->23	
ålln	a->1	i->66	
ålls	 ->4	,->1	.->1	a->2	l->2	m->2	r->2	t->7	v->1	
ålme	d->1	
ålni	n->3	
ålsd	o->1	
ålse	k->5	n->2	
ålsk	y->1	
ålss	i->1	
ålst	i->1	
ålsä	t->17	
ålun	d->4	
ålve	r->5	
åläg	g->6	
åmin	d->1	n->29	
ån (	H->21	
ån -	 ->2	
ån 1	0->1	5->1	9->5	
ån 2	8->1	
ån 3	,->1	
ån 5	 ->2	0->1	
ån 8	9->1	
ån 9	5->1	
ån A	f->1	l->2	m->4	t->2	u->1	
ån B	S->1	a->1	o->1	r->2	
ån C	E->2	a->1	
ån D	a->1	e->1	
ån E	G->2	U->1	r->2	u->24	
ån F	M->1	l->3	r->1	ö->1	
ån G	U->1	a->1	o->1	ö->1	
ån H	e->2	
ån I	R->1	n->3	s->1	
ån J	a->1	
ån K	o->1	y->2	ö->2	
ån L	a->1	i->1	o->1	
ån M	a->1	
ån N	a->3	
ån O	S->1	
ån P	P->2	S->1	a->1	o->3	
ån R	o->1	
ån S	a->3	h->1	y->2	
ån T	a->4	e->1	y->1	
ån U	N->1	S->1	
ån V	e->1	
ån W	i->1	u->1	
ån a	l->4	n->3	t->26	v->3	
ån b	e->1	i->4	o->2	u->2	ö->5	
ån d	a->3	e->89	i->4	o->1	r->1	ä->1	
ån e	n->19	r->3	t->17	u->1	x->3	
ån f	a->2	l->2	r->2	ö->39	
ån g	e->4	
ån h	a->4	e->1	ö->2	
ån i	 ->3	
ån j	u->4	
ån k	a->3	o->34	
ån l	a->1	e->3	i->1	ä->4	
ån m	a->4	e->7	i->8	o->2	å->2	
ån n	a->1	y->2	å->3	
ån o	b->1	c->11	f->1	l->4	m->1	p->1	r->2	s->2	
ån p	a->13	e->1	r->4	å->3	
ån r	a->1	e->3	å->13	
ån s	a->3	e->1	i->8	k->3	o->2	t->4	y->1	ä->3	å->1	ö->1	
ån t	.->1	i->5	o->2	r->16	u->1	
ån u	n->2	t->20	
ån v	a->2	e->1	i->5	ä->1	å->10	
ån Ö	s->1	
ån ä	r->1	
ån å	r->1	
ån ö	v->4	
ån, 	d->1	f->1	n->1	o->1	
ån.D	e->3	ä->1	
ån.H	ä->1	
ån.Ä	n->1	
åna 	m->1	o->3	
ånad	 ->9	,->2	.->3	e->59	s->1	
ånan	d->2	
ånar	 ->1	e->6	n->5	
ånas	 ->1	
ånbo	k->1	
ånd 	a->5	d->2	e->7	f->7	h->2	i->5	k->2	m->3	n->1	o->7	p->1	s->5	t->4	v->1	ä->1	å->1	
ånd,	 ->8	
ånd.	 ->1	A->1	D->3	F->1	H->1	J->1	V->2	
ånd?	.->1	J->1	
ånda	g->3	r->5	
ånde	.->1	l->1	n->10	t->19	
åndi	g->1	
åndp	u->97	
ånds	 ->1	d->12	p->2	r->1	s->1	t->2	
åner	 ->1	.->1	
ång 	-->1	a->9	b->5	d->6	e->6	f->12	h->6	i->7	k->4	l->1	m->2	n->1	o->6	p->6	r->4	s->20	t->34	u->6	v->6	ä->4	ö->1	
ång"	.->1	
ång,	 ->11	
ång.	D->5	F->1	H->1	J->1	N->2	O->1	T->1	V->2	
ånga	 ->157	,->2	.->2	r->16	s->1	
ångd	r->1	
ånge	l->1	n->45	r->26	t->1	
ångf	a->15	r->1	u->1	ä->2	
ångk	ö->1	
ångl	i->1	
ångm	å->1	
ångn	a->2	
ångr	a->2	e->1	
ångs	 ->3	a->8	b->3	f->1	i->10	p->15	r->15	s->9	t->8	ä->1	
ångt	 ->34	.->3	g->11	i->4	
ångv	a->6	
ångå	r->1	
ånin	g->7	
ånko	m->3	
ånsp	a->1	
ånta	r->1	s->1	
ånto	g->1	
ånva	r->8	
ånvä	n->1	
ånyo	 ->1	
åolj	a->1	
åpek	a->50	
åpsl	a->1	
år -	 ->1	
år 1	9->19	
år 2	0->33	
år B	a->1	
år M	a->1	
år O	L->1	
år a	d->1	k->1	l->5	n->3	r->1	t->32	v->15	
år b	a->1	e->11	i->1	o->2	r->2	u->1	
år d	e->49	i->5	j->1	o->1	r->1	u->1	ä->5	å->2	
år e	f->4	g->2	l->3	m->1	n->25	r->5	t->9	
år f	a->4	e->1	i->2	o->3	r->22	å->1	ö->26	
år g	e->8	i->1	l->1	r->16	ö->2	
år h	a->5	e->8	ä->3	å->1	ö->1	
år i	 ->42	b->1	d->1	f->2	g->3	n->72	
år j	a->13	u->1	
år k	a->3	l->9	o->14	r->1	u->1	v->1	
år l	a->2	e->2	i->4	o->2	y->1	ä->1	å->2	
år m	a->2	e->11	i->10	o->8	y->4	å->2	ö->2	
år n	a->1	i->1	o->1	u->2	y->1	ä->1	å->2	ö->2	
år o	c->17	f->2	m->3	r->4	s->1	
år p	a->1	e->1	l->3	o->4	r->3	å->19	
år r	e->8	o->3	ä->2	ö->2	
år s	a->3	e->18	i->5	j->2	k->6	l->1	n->3	o->13	p->1	t->14	v->1	ä->1	å->2	
år t	a->6	i->32	r->2	v->1	
år u	n->7	p->7	t->15	
år v	a->5	e->2	i->34	ä->4	
år y	t->1	
år ä	g->1	n->2	r->3	v->2	
år å	 ->1	s->3	t->5	
år ö	n->2	p->1	v->2	
år".	J->1	
år)?	 ->1	
år, 	E->1	a->1	d->2	e->2	f->1	i->1	k->3	m->4	n->2	o->6	p->1	s->2	t->1	u->3	v->1	ä->1	
år. 	E->1	J->1	
år.D	e->12	
år.E	n->1	
år.F	ö->2	
år.H	e->2	u->1	ä->1	
år.I	 ->2	
år.J	a->4	
år.K	ä->1	
år.L	a->1	y->1	
år.M	a->1	
år.O	m->1	
år.R	e->1	
år.S	a->1	
år.T	y->1	
år.V	e->1	i->4	å->1	
år.Ä	n->1	
år?N	ä->1	
år?S	o->1	
åra 	a->12	b->4	d->5	e->10	f->19	g->7	h->3	i->5	k->13	l->13	m->19	n->2	o->2	p->9	r->16	s->14	t->6	u->1	v->4	ä->5	å->6	ö->4	
åra,	 ->1	
åran	d->1	
årar	 ->1	e->4	
åras	,->1	
årat	a->1	
årba	r->3	
årbe	d->1	g->1	
ård 	g->1	k->1	o->2	p->1	t->1	
ård)	,->1	
ård,	 ->2	
årda	 ->7	g->2	r->5	s->2	
årde	n->1	
årdn	a->2	
årds	-->1	l->2	m->1	
åren	 ->27	,->5	.->6	s->2	
året	 ->30	,->8	.->3	s->4	
århu	n->7	
årig	a->7	h->31	t->7	
årin	g->1	
årkl	y->1	
årkö	t->1	
årli	g->8	
årlö	s->2	
årni	n->2	
års 	E->1	b->3	e->1	p->1	s->1	t->3	ö->1	
årsa	f->1	
årsb	e->2	
årsp	e->1	r->1	
årsr	a->2	
årss	k->2	
årst	i->1	
årt 	E->2	a->36	b->3	d->6	e->10	f->14	g->3	h->1	i->2	k->4	l->5	m->6	n->2	o->3	p->13	r->3	s->15	t->2	u->12	v->3	y->1	
årt,	 ->3	
årt.	M->1	
årta	l->1	
årti	o->1	
årtu	s->3	
åröv	e->1	
ås a	l->1	t->2	v->1	
ås b	l->2	ä->1	
ås d	e->2	ä->1	
ås e	n->2	
ås f	a->1	ö->3	
ås g	e->2	ö->1	
ås i	 ->13	g->1	n->1	
ås k	o->1	
ås m	o->1	
ås o	c->1	
ås p	å->1	
ås s	k->1	
ås t	i->2	
ås u	p->1	
ås v	a->1	
ås, 	i->1	
ås.D	e->1	
ås.F	ö->1	
ås.L	a->1	
ås: 	a->1	
åsam	k->3	
åsat	t->1	
åser	 ->3	
åsik	t->50	
åska	l->1	
åsky	n->7	
åskå	d->2	
åsom	 ->34	
åss 	m->1	
åst 	s->1	
åsta	 ->2	d->25	
åste	 ->693	,->3	
åstr	i->1	
åstå	 ->4	,->2	e->8	r->4	s->2	t->1	
åsyf	t->5	
åt E	u->1	
åt F	ö->1	
åt a	n->1	t->7	
åt b	e->1	
åt d	e->27	
åt e	g->1	n->3	r->2	t->2	
åt f	o->1	r->1	
åt g	e->1	
åt h	u->1	
åt i	 ->8	m->1	n->2	
åt j	ä->1	
åt k	o->4	v->1	
åt l	i->1	
åt m	a->1	e->2	i->55	o->1	
åt n	u->1	y->1	
åt o	c->2	s->26	
åt p	a->1	å->1	
åt r	e->1	ä->3	
åt s	a->1	i->4	y->1	
åt t	i->1	v->1	ä->1	
åt u	n->1	
åt v	e->1	å->1	
åt Ö	s->1	
åt ä	m->1	r->2	
åt å	t->1	
åt",	 ->1	
åt, 	i->1	k->1	m->2	u->1	
åt.D	a->1	e->1	ä->1	
åt.F	r->1	
åt.H	e->1	
åt.J	a->1	
åt.K	o->1	
åt.N	ä->1	
åt.V	a->1	
åta 	E->1	J->1	a->2	b->3	d->10	e->2	f->2	h->1	j->1	k->1	l->1	m->4	n->1	o->2	p->2	r->2	s->7	t->1	
åtag	a->28	i->2	l->4	
åtal	 ->6	.->1	a->10	s->7	
åtan	d->3	k->1	
åtar	 ->7	,->2	n->1	
åtas	 ->6	
åte 	s->1	
åten	 ->4	h->2	s->1	
åter	 ->41	,->1	.->1	a->18	b->1	e->1	f->13	g->7	h->4	i->25	k->8	l->2	n->11	s->33	t->9	u->32	v->71	
åtet	 ->1	
åtfö	l->12	
åtgä	r->240	
åtgå	n->1	
åtil	l->1	
åtit	 ->2	s->1	
åtli	g->5	
åtmi	n->27	
åtna	 ->5	.->1	
åtnj	u->1	
åtry	c->3	
åts 	e->1	f->1	m->1	å->1	
åtsa	s->2	
åtsk	i->3	
åtst	r->3	
ått 	-->1	8->1	9->1	E->1	K->1	a->7	b->3	d->5	e->22	f->6	g->1	h->5	i->12	j->1	k->3	l->1	m->10	n->7	o->4	p->2	s->5	t->11	u->4	v->8	y->3	ä->1	å->1	
ått,	 ->2	
ått.	D->2	F->1	I->2	P->2	
åtta	 ->4	,->1	
åttf	u->1	
åtto	 ->2	n->1	r->1	
åtts	 ->7	.->2	
åtvi	n->4	
åvar	 ->1	a->1	
åver	k->37	
åvid	a->3	
åvil	a->1	
åvis	a->2	b->1	
åvor	 ->1	.->1	
åväl	 ->41	
åzon	 ->1	
ça M	o->5	
çois	 ->1	
ère 	k->1	
ète 	s->1	
ève 	1->1	
ève,	 ->1	
èvek	o->1	
é - 	f->1	o->2	
é at	t->2	
é av	e->1	
é el	l->1	
é fö	r->3	
é ha	r->1	
é ja	g->1	
é ko	m->1	
é me	d->1	
é oc	h->3	
é om	 ->1	
é pe	r->1	
é so	m->5	
é ut	a->1	
é är	 ->1	
é, m	e->1	
éavt	a->1	
ébet	o->1	
ébé 	a->1	
écha	r->1	
ée, 	v->1	
éer 	a->1	i->2	m->1	o->2	s->3	t->1	
éer,	 ->3	
éer.	D->1	
éern	a->7	
éfér	e->1	
éför	f->2	
ékon	v->1	
én (	C->2	
én a	t->6	
én b	a->1	e->1	ö->1	
én f	ö->3	
én i	 ->1	
én k	o->1	
én l	a->1	
én m	e->1	
én o	c->4	m->11	
én s	a->1	i->1	
én v	a->1	i->1	
én ä	r->1	
én, 	k->1	o->1	s->1	u->1	v->1	
én.H	u->1	
én.M	e->1	
én.W	o->1	
én?V	i->1	
éns 	a->2	g->6	r->2	s->1	
éren	d->1	
érys	 ->1	
és R	u->1	
ésys	t->2	
étai	n->1	
éuni	o->2	
ête 	o->3	
êts 	(->1	
í är	 ->1	
íez 	G->1	
ínci	p->1	
ón C	r->2	
ón i	 ->1	
ón t	i->1	
ón v	i->1	
ónio	 ->1	
ône-	A->1	
ö fö	r->2	
ö i 	d->1	e->1	
ö ka	n->1	
ö mo	t->1	
ö sa	k->1	
ö so	m->1	
ö vi	n->1	
ö!De	t->1	
ö, f	o->7	ö->1	
ö, h	ä->1	
ö, l	i->1	
ö, s	m->1	
ö, u	p->1	
ö- o	c->2	
ö.De	t->3	
ö.Då	 ->1	
ö.Me	n->1	
ö.Un	d->1	
ö.Vi	l->1	
öanp	a->1	
öans	v->2	
öar 	s->1	
öarn	a->5	
öavt	a->1	
öbel	a->1	
öbes	k->1	t->1	
öble	r->2	
öbo 	v->1	
öbro	t->1	
öcke	r->3	
öd -	 ->2	
öd a	n->1	v->4	
öd b	i->1	
öd d	e->2	ä->1	
öd e	f->1	n->2	
öd f	r->7	ö->20	
öd g	e->1	
öd h	a->1	o->1	
öd i	 ->6	b->1	n->5	
öd k	a->4	o->1	
öd l	ö->1	
öd m	e->2	å->3	
öd o	c->14	m->4	
öd p	e->1	r->1	å->5	
öd s	k->1	o->18	å->1	
öd t	i->43	
öd v	a->2	i->4	
öd ä	n->2	
öd å	t->2	
öd ö	k->1	
öd, 	d->1	e->1	m->1	o->3	s->7	u->1	
öd."	J->1	
öd.-	 ->1	
öd..	(->1	
öd.A	l->1	t->1	
öd.D	e->10	ä->1	å->1	
öd.E	u->1	
öd.F	ö->2	
öd.H	a->1	e->4	
öd.I	 ->2	
öd.J	a->3	
öd.M	e->1	o->1	
öd.N	i->1	
öd.O	r->1	
öd.R	e->1	
öd.S	å->1	
öd.T	r->1	
öd.U	t->1	
öd.V	i->2	
öd.Ä	n->1	v->1	
öd.Å	 ->1	r->1	
öd; 	d->1	
öd?-	 ->1	
öda 	o->3	s->1	t->2	
öda"	 ->1	
öda,	 ->1	
ödad	e->3	
ödan	d->5	
ödas	 ->1	,->1	
ödat	s->1	
ödbe	d->1	
ödd.	M->1	
ödde	 ->1	s->2	
öde 	i->1	u->1	
öde,	 ->4	
öde.	D->1	
öde?	H->1	
ödel	a->1	s->5	
ödem	a->1	
öden	 ->23	,->2	.->4	a->1	s->4	
ödep	a->1	
öder	 ->59	,->1	.->1	m->2	
ödes	b->1	d->2	g->1	
ödet	 ->29	,->1	.->2	s->2	
ödfö	d->1	
ödgr	ö->1	
ödig	 ->2	.->1	a->3	t->7	
ödin	s->1	
ödir	e->1	
ödja	 ->62	.->2	s->7	
ödje	r->1	
ödme	d->1	
ödmo	t->1	
ödni	n->1	v->1	
ödor	.->1	
ödos	a->1	
ödoä	m->1	
ödpo	l->1	
ödra	 ->6	m->2	r->1	
öds 	a->5	b->1	e->1	g->1	j->1	t->1	
ödsd	ö->1	
ödsf	a->1	
ödsi	t->1	
ödsp	o->1	
ödsy	s->4	
ödvä	n->125	
ödåt	g->5	
öend	e->1	
öer 	f->1	i->1	s->1	
öern	a->1	
öfak	t->1	
öfar	l->1	t->8	
öfrå	g->4	
öfte	 ->3	n->8	
öför	b->1	h->1	s->2	
ög a	r->1	
ög b	e->1	
ög f	e->1	
ög g	r->6	
ög i	n->1	
ög k	v->1	
ög n	i->2	
ög p	r->2	
ög s	e->1	k->1	o->1	t->2	y->1	
ög, 	d->1	
öga 	f->1	g->1	k->3	m->1	n->1	p->1	r->3	s->1	t->2	å->2	
öga,	 ->1	
öga.	M->1	
ögak	t->1	
ögat	.->1	
öge 	k->1	r->1	
ögel	m->1	
öger	 ->2	,->1	e->6	m->1	n->19	p->1	v->1	
öghe	t->3	
öglj	u->1	
ögna	 ->1	
ögni	v->3	
ögon	 ->5	,->1	b->13	
ögra	 ->1	
ögre	 ->18	.->1	
ögsk	o->1	
ögst	 ->11	,->1	a->16	
ögt 	f->1	i->2	p->3	s->1	u->1	v->1	
ögt,	 ->1	
ögt.	S->1	
ögte	k->2	
ögti	d->4	
öinf	o->1	
öja 	J->1	d->4	f->1	k->1	l->1	m->1	o->5	s->2	t->1	
öja.	V->1	
öjad	e->1	
öjak	t->2	
öjan	d->2	
öjar	 ->3	e->1	
öjas	.->3	
öjd 	-->1	a->1	g->1	m->1	p->1	s->1	u->1	
öjda	 ->6	,->3	
öjde	 ->2	n->1	r->3	
öjdp	u->2	
öje 	B->1	E->1	f->1	o->1	
öjel	s->1	
öjer	 ->5	
öjet	 ->2	
öjev	ä->3	
öjli	g->309	
öjni	n->2	
öjor	.->1	
öjs 	t->1	
öjsm	å->2	
öjt 	o->1	s->1	
öjts	 ->1	,->1	
ök a	t->4	
ök b	e->1	
ök i	 ->5	
ök o	m->1	
ök s	o->1	
ök, 	d->1	o->1	s->1	
öka 	F->1	a->11	b->3	d->4	e->3	f->12	g->2	h->3	i->2	j->1	k->8	m->4	o->3	s->8	t->1	u->5	v->4	å->1	
öka,	 ->1	
öka.	O->1	R->1	T->1	
ökad	 ->28	e->9	
ökan	d->11	
ökar	 ->12	,->3	.->1	l->6	
ökas	 ->5	,->2	.->3	t->1	
ökat	 ->16	.->1	a->10	
öke 	d->1	
öke.	M->1	
öken	 ->2	
öker	 ->21	
öket	 ->4	
ökmo	d->1	
ökni	n->43	
ökon	f->1	s->5	
ökra	v->8	
öks,	 ->1	
öksb	o->1	
ökst	ä->1	
ökt 	F->1	a->5	b->1	d->1	e->1	f->1	h->1	o->1	u->1	v->1	
ökte	 ->6	
ökva	l->1	
öl n	ä->1	
öl o	c->1	
öl, 	s->1	
ölag	s->1	
ölar	.->1	
öld 	m->1	
öld,	 ->1	
öldb	e->1	
öldg	r->1	
ölja	 ->31	,->1	.->1	k->14	n->37	r->1	s->6	
öljd	 ->18	.->1	e->21	r->1	s->2	å->1	
ölje	l->3	r->17	
öljn	i->10	
öljs	 ->4	,->1	
öljt	 ->2	s->2	
öll 	K->1	a->3	d->3	e->4	i->2	m->1	n->1	o->2	s->1	t->1	ö->1	
öll.	H->1	
ölls	 ->4	
öln 	a->1	i->1	
öm a	v->2	
öm b	e->1	
öm i	n->1	
öm t	a->1	
öm, 	s->1	
öm: 	N->1	
öma 	H->2	a->3	d->4	e->2	f->2	h->2	i->1	o->3	p->1	r->1	s->2	t->1	v->2	
öma,	 ->1	
öma.	D->1	
öman	d->7	
ömas	 ->2	
ömba	r->1	
ömd,	 ->2	
ömde	.->1	s->1	
öme.	K->1	
ömer	 ->9	
ömes	g->1	
ömin	i->1	
ömli	g->2	
ömma	 ->15	:->1	n->3	r->3	s->1	
ömme	n->4	r->5	
ömni	n->34	
öms 	e->2	v->1	
ömse	s->5	
ömsk	a->1	
ömt 	A->1	W->1	a->1	b->3	e->1	p->1	s->1	v->1	
ömts	 ->2	
ömtå	l->1	
ömvä	r->1	
ömän	 ->2	
ömäs	s->11	
ömål	 ->2	s->1	
ön N	o->1	
ön e	l->1	n->1	
ön f	ö->2	
ön h	å->1	
ön i	 ->1	
ön o	c->6	
ön p	å->1	
ön s	o->2	
ön t	i->1	
ön v	ä->2	
ön ä	r->1	
ön!D	e->1	
ön, 	a->1	d->1	h->1	m->1	o->3	s->1	u->1	
ön.D	e->2	ä->1	
ön.E	n->1	
ön.F	r->1	
ön.J	a->1	
ön.L	å->1	
ön.M	a->1	
ön.U	n->1	
ön.V	i->1	å->1	
öna 	e->1	f->1	g->2	h->2	i->1	m->1	n->1	o->1	p->1	s->2	
öna/	E->1	
önar	 ->1	e->1	
önas	 ->2	,->1	
önbo	k->1	
önde	r->7	
öne-	 ->1	
önea	r->1	
önen	 ->3	
öner	 ->2	
önhe	t->1	
önit	z->1	
önk 	h->1	r->1	u->1	
önk.	D->1	
önor	m->2	
öns 	f->1	s->1	
önsa	m->5	
önsg	r->1	
önsk	a->54	e->3	n->2	v->10	
önst	e->2	r->1	
önt 	a->1	l->1	
önta	g->3	
öomr	å->4	
öovä	n->1	
öp a	v->2	
öpa 	d->1	e->1	u->1	
öpan	d->6	
öpar	e->3	n->1	
öpen	h->1	
öper	 ->12	.->1	s->1	
öpkr	a->1	
öpol	i->8	
öppe	n->65	t->14	
öppn	a->16	i->4	
öpro	b->3	g->1	
öpsb	e->1	
öpsl	a->1	
öpt 	i->1	u->5	
öpte	 ->3	
öpåv	e->1	
ör "	K->1	a->2	f->1	i->1	n->1	
ör -	 ->6	,->1	
ör 1	9->17	
ör 2	0->5	7->1	9->1	
ör 3	 ->1	3->1	
ör 5	 ->1	,->1	
ör 7	5->1	6->1	
ör 8	1->1	
ör A	g->1	l->3	
ör B	e->1	i->1	o->1	r->3	
ör C	S->1	e->1	
ör D	a->2	e->1	
ör E	C->1	G->4	U->9	r->1	u->60	
ör F	P->1	o->2	ö->2	
ör G	e->1	o->1	
ör H	a->1	
ör I	M->1	N->1	n->1	s->1	
ör K	a->3	o->1	u->2	y->1	
ör L	a->1	e->1	
ör M	o->1	
ör O	L->1	
ör P	P->1	a->1	o->2	
ör S	a->2	ã->1	
ör T	a->1	i->6	u->1	
ör V	o->1	
ör W	T->1	a->1	
ör a	b->2	c->1	i->1	l->141	m->2	n->46	r->15	s->3	t->778	v->26	
ör b	a->3	e->44	i->11	j->1	l->6	o->3	r->4	u->14	ä->1	å->3	ö->6	
ör c	e->2	h->1	i->4	
ör d	a->4	e->684	i->11	j->1	o->4	u->2	ä->7	å->4	ö->1	
ör e	f->1	g->4	k->16	l->5	m->1	n->149	r->34	t->57	u->1	v->2	x->3	
ör f	a->11	e->3	i->12	j->1	l->5	o->10	r->33	u->3	y->1	å->8	ö->68	
ör g	a->1	e->23	i->3	l->1	o->4	r->16	u->2	ä->1	ö->8	
ör h	a->39	e->23	i->1	j->3	o->6	u->12	ä->10	å->3	ö->5	
ör i	 ->19	c->1	h->2	k->1	l->1	n->62	
ör j	a->14	o->11	u->4	ä->3	
ör k	a->19	l->1	n->1	o->104	r->10	u->23	v->9	ä->6	
ör l	a->9	e->3	i->28	o->3	ä->15	å->7	ö->1	
ör m	a->34	e->52	i->60	o->6	y->15	ä->14	å->29	ö->3	
ör n	a->11	e->2	i->2	o->9	u->3	y->7	ä->42	å->19	ö->3	
ör o	c->19	f->13	l->5	m->14	p->1	r->7	s->56	t->1	v->2	
ör p	a->23	e->26	l->1	o->6	r->19	u->1	å->5	
ör r	a->2	e->60	i->4	o->1	ä->28	å->9	ö->6	
ör s	a->16	e->10	i->54	j->5	k->31	l->2	m->5	n->4	o->5	p->4	t->59	v->3	y->20	ä->17	å->13	
ör t	.->2	a->7	e->2	i->53	j->7	o->1	r->26	u->3	v->8	y->4	å->1	
ör u	n->40	p->12	r->2	t->67	
ör v	a->39	e->12	i->76	o->1	u->1	ä->5	å->43	
ör y	n->1	r->1	t->2	
ör Ö	s->2	
ör ä	g->1	n->8	r->26	v->4	
ör å	k->1	r->12	t->26	
ör ö	a->1	g->7	k->3	p->5	r->1	s->1	v->34	
ör".	O->1	
ör, 	1->1	B->1	a->6	e->2	f->3	h->1	i->2	k->3	m->1	o->4	s->3	t->1	u->1	v->1	ä->2	
ör. 	D->1	E->1	
ör.(	L->1	
ör..	.->1	
ör.D	e->6	i->1	
ör.E	t->1	
ör.F	ö->1	
ör.H	e->1	
ör.J	a->1	
ör.K	o->1	
ör.M	a->1	e->2	
ör.V	i->4	å->1	
ör: 	D->1	F->1	a->1	
ör; 	d->1	
ör?D	ä->1	
ör?F	r->2	
ör?I	 ->1	
ör?Ä	r->1	
öra 	-->1	E->3	a->27	b->7	d->101	e->72	f->24	g->8	h->6	i->12	k->14	l->5	m->41	n->25	o->7	p->10	r->6	s->38	t->10	u->16	v->15	y->2	ä->5	å->2	ö->2	
öra,	 ->9	
öra.	D->5	E->2	H->1	I->1	J->4	L->1	N->1	O->1	P->1	S->1	
öra?	J->1	
örak	t->1	
öral	l->1	
öran	d->389	k->4	l->2	s->1	
örar	b->1	l->1	n->1	
öras	 ->60	!->2	,->5	.->16	;->1	
örba	n->2	r->12	
örbe	h->6	r->27	
örbi	 ->1	f->2	g->6	n->22	s->1	
örbj	u->14	
örbl	e->1	i->14	
örbr	u->1	y->2	ä->2	
örbu	d->26	n->12	
örbä	t->78	
örd 	a->2	f->1	k->1	m->1	o->1	
örd,	 ->1	
örd.	D->2	
örda	 ->29	,->2	.->3	?->1	d->2	g->1	n->9	r->1	t->2	
örde	 ->19	,->1	.->2	l->42	n->7	s->11	
ördh	e->1	
ördj	u->11	
ördn	a->1	
ördo	m->2	r->2	
ördr	a->164	ö->1	
ördu	b->2	n->1	
ördä	r->4	
ördö	m->20	
öre 	2->1	A->1	K->1	d->5	e->1	m->3	n->2	o->3	s->2	u->4	v->2	å->1	ö->1	
öreb	i->1	r->2	y->23	
öred	r->166	ö->2	
öref	a->20	ö->1	
öreg	i->8	r->1	å->17	
öreh	a->1	
örek	o->22	
örel	e->1	i->26	s->21	
örem	å->13	
ören	 ->1	,->1	a->25	i->12	k->8	l->9	s->1	t->28	
örer	 ->6	,->3	.->4	n->10	
öres	a->6	k->28	l->104	p->10	t->15	ä->1	
öret	a->200	r->73	
örfa	l->1	r->76	t->7	
örfi	n->1	
örfj	o->1	
örfl	u->14	y->4	
örfo	g->18	
örfr	y->1	å->4	
örfä	k->1	r->2	
örfå	n->1	
örfö	l->5	
örg 	H->14	
örgl	ö->2	
örgr	u->3	
örgä	v->1	
örha	n->92	s->3	
örhi	n->31	
örho	p->12	
örhå	l->56	
örhö	l->1	
örig	 ->2	a->2	h->15	t->2	
örin	g->16	t->5	
örir	r->1	
örja	 ->68	d->8	n->19	r->17	t->12	
örjd	e->1	
örje	r->2	
örjn	i->4	
örk 	d->1	
örka	s->9	
örkl	a->76	ä->1	
örkn	i->3	
örko	r->2	
örkr	o->1	
örku	n->2	
örla	g->3	
örle	g->2	
örli	g->39	k->45	n->1	s->2	t->10	v->19	
örlo	r->20	
örlu	s->10	
örlä	g->2	n->4	
örlå	t->4	
örme	d->3	n->2	
örmi	d->3	
örmo	d->12	
örmy	n->1	
örmå	 ->2	g->31	n->14	r->1	
örmö	g->1	
örn 	d->1	f->1	
örna	m->1	
örne	d->2	k->8	
örni	n->7	
örns	t->1	
örnu	f->14	
örny	a->4	b->39	e->6	
örol	ä->2	
öron	,->1	m->2	
öror	d->44	e->28	s->6	
örpa	c->5	s->1	
örpl	i->21	
örr 	d->1	e->2	ö->1	
örr,	 ->2	
örra	 ->42	r->3	
örre	 ->77	n->4	s->2	
örrg	å->3	
örri	n->1	
örrä	d->1	n->4	
örrå	d->1	
örs 	a->17	b->1	d->1	e->6	f->7	i->8	k->1	m->2	o->1	p->5	t->1	u->1	ä->1	ö->2	
örs,	 ->7	
örs.	 ->1	.->1	D->2	H->1	J->2	O->1	V->1	
örsa	m->12	
örse	 ->2	n->28	r->2	s->1	
örsi	k->67	
örsk	a->2	i->2	j->1	o->2	r->4	ä->1	å->1	
örsl	a->492	
örso	m->1	n->5	
örsp	o->1	
örst	 ->75	.->2	a->246	e->1	k->1	o->3	ä->30	å->83	ö->21	
örsu	m->9	
örsv	a->62	i->15	u->4	å->2	
örsä	k->44	l->5	m->10	n->1	
örså	g->1	
örsö	k->61	r->4	
ört 	-->2	D->1	a->1	d->5	e->7	f->6	i->3	k->1	l->1	m->12	n->2	o->2	p->3	s->6	t->2	u->2	v->2	
ört,	 ->3	
ört.	J->1	K->1	
örte	c->3	
örti	d->6	
örtj	u->1	ä->20	
örtn	i->1	
örtr	o->60	y->2	ä->3	ö->1	
örts	 ->27	,->3	.->4	
örtv	i->1	
örty	d->3	
örtä	c->1	
örun	d->1	
örut	 ->2	.->1	b->1	o->15	s->63	v->2	
örva	l->49	n->6	r->1	
örve	r->22	
örvi	r->12	s->9	
örvr	ä->1	
örvä	g->14	n->29	r->11	
örvå	n->6	
örän	d->74	
öråd	e->1	
örål	d->3	
öröd	a->3	e->2	
örör	e->2	
öröv	a->3	
ös -	 ->1	
ös d	a->1	e->1	
ös e	n->1	
ös k	ä->1	
ös o	c->2	
ös p	o->1	
ös r	a->1	
ös s	k->1	u->1	
ös u	t->1	
ös, 	k->1	
ös.D	e->1	
ösa 	a->1	d->9	e->2	f->1	g->2	h->1	i->1	k->2	m->8	n->1	o->3	p->8	r->1	s->4	u->2	v->4	
ösa,	 ->4	
ösa.	A->1	F->1	I->1	M->1	
ösar	 ->1	e->2	
ösas	 ->5	.->1	
ösek	t->1	
öser	 ->1	i->3	
öses	 ->1	
ösgö	r->1	
öshe	t->44	
ösid	a->1	
öska	d->2	
öske	l->3	
ösky	d->11	
öskä	l->2	
ösni	n->52	
ösry	c->1	
öss 	o->1	p->1	ä->1	
öss)	 ->1	
össo	r->1	
öst 	-->2	a->2	d->2	f->2	h->3	i->4	l->1	m->1	o->5	p->2	r->1	s->3	t->2	v->1	
öst,	 ->3	
öst.	J->1	Ä->1	
östa	 ->47	,->1	.->4	d->15	r->15	t->15	
östb	l->1	
öste	d->4	n->1	r->72	s->1	u->3	
östf	ö->7	
östl	ä->1	
östn	i->57	
östr	a->3	ä->3	
östs	.->1	
östt	o->1	
östu	t->2	
östv	i->3	
östö	d->1	
ösyn	p->6	
öt 9	3->1	
öt a	t->1	
öt d	e->1	
öt h	a->1	
öt l	o->1	
öt t	a->4	
öt v	i->1	
öt.D	e->1	
öta 	E->1	d->8	e->1	m->2	p->1	s->3	v->1	
ötan	d->1	
ötar	 ->1	
ötas	 ->1	
öte 	d->1	i->4	k->1	m->4	o->1	p->1	s->1	
öteb	o->1	
öten	 ->2	a->2	
öter	 ->43	!->14	,->7	.->1	n->24	s->1	
ötes	 ->1	.->1	g->3	t->1	
ötet	 ->19	.->2	
ötfå	n->1	
ötkö	t->3	
ötra	n->1	
öts 	a->1	b->1	i->1	k->2	m->1	
öts.	V->1	
ötse	l->5	
ötsk	a->1	
ötsl	i->4	
ött 	B->1	F->1	d->2	k->1	o->1	p->2	s->3	t->1	u->1	v->2	ä->1	
ött.	D->2	J->1	
ötta	 ->1	,->1	t->2	
ötte	 ->2	r->8	s->1	
öttk	r->1	
öttr	a->1	
ötts	 ->2	-->1	p->1	
öuts	k->1	
öva 	E->1	a->1	d->1	e->3	f->1	g->3	h->1	k->2	l->1	n->1	p->3	r->1	s->2	t->1	u->2	v->1	ö->1	
övad	e->2	
övan	d->1	
övar	 ->5	e->2	
övas	 ->6	.->3	
övat	 ->1	s->1	
övde	 ->2	
över	 ->311	,->5	.->10	a->9	b->9	c->1	d->14	e->71	f->23	g->41	h->4	i->1	k->6	l->35	m->2	n->4	o->1	p->1	r->4	s->70	t->54	v->71	
övit	t->1	
övla	d->1	
övli	g->1	
övni	n->12	
övoå	r->1	
övra	d->1	n->1	r->1	
övri	g->65	
övs 	d->3	e->6	f->2	i->3	m->1	n->1	o->1	p->1	s->2	
övs,	 ->2	
övs.	D->1	F->1	I->1	S->2	
övsk	o->1	
övst	a->1	
övt 	f->1	s->1	t->1	
övts	 ->1	
övän	l->7	
övär	d->3	
öw f	ö->1	
öy -	 ->1	
ööw 	f->1	
øn, 	i->1	m->1	
ørge	n->2	
ührk	o->1	
ünch	e->1	
ürkd	a->1	
üsse	l->4	
