 "	A->2	B->1	D->4	E->4	J->1	K->7	L->1	M->2	O->2	P->1	T->3	U->1	a->8	b->1	c->1	d->5	e->9	f->2	g->2	h->2	i->3	j->1	k->4	l->3	m->1	n->4	o->3	p->2	r->6	s->5	t->1	u->2	v->2	å->1	ö->2	
 '	V->1	
 (	"->1	1->4	5->1	8->2	9->1	A->35	B->7	C->11	D->1	E->29	F->16	H->22	I->4	K->10	P->16	S->2	U->2	a->9	d->2	e->4	f->8	h->1	i->4	k->6	m->3	o->1	r->2	s->2	t->2	u->1	Ö->5	å->1	
 ,	 ->5	
 -	 ->551	(->1	,->9	e->1	o->3	
 0	 ->1	0->27	1->1	5->1	6->1	
 1	 ->28	,->8	-->12	.->1	/->1	0->29	1->18	2->28	3->20	4->16	5->22	6->14	7->13	8->10	9->223	
 2	 ->19	,->8	-->3	.->4	0->117	1->10	2->8	3->3	4->7	5->18	6->7	7->7	8->12	9->7	
 3	 ->9	,->3	-->3	.->3	0->12	1->7	2->4	3->8	4->7	5->8	6->3	7->8	8->6	9->4	:->1	
 4	 ->13	,->4	.->4	0->18	1->5	2->4	3->2	4->3	5->9	6->3	7->1	8->5	
 5	 ->13	,->5	.->2	0->12	1->1	2->4	3->1	4->1	5->2	6->2	7->1	b->3	
 6	 ->16	,->3	.->1	0->4	2->1	7->1	8->2	
 7	 ->18	)->1	,->7	.->1	0->6	3->1	5->3	6->1	7->1	9->1	
 8	 ->9	,->2	0->14	1->16	2->8	3->1	5->4	6->3	7->3	8->5	9->2	
 9	 ->8	,->2	.->1	0->6	1->1	2->1	3->2	4->7	5->5	6->5	7->2	8->1	
 :	 ->1	
 A	.->1	B->4	D->1	K->1	c->1	d->5	f->4	g->2	h->7	i->1	k->3	l->36	m->44	n->7	p->1	r->8	s->5	t->8	u->3	v->5	z->2	
 B	 ->2	N->16	P->1	R->1	S->6	a->41	e->51	i->6	l->3	o->15	r->39	u->4	y->3	
 C	.->2	4->6	5->15	E->11	S->2	a->17	e->13	h->2	l->1	o->20	r->2	u->3	y->1	
 D	 ->1	D->1	a->43	e->146	i->7	o->2	u->12	ä->7	å->2	í->1	ü->1	
 E	-->1	C->3	D->3	E->3	G->53	I->1	K->5	L->3	M->6	U->138	c->1	d->1	f->11	g->2	h->2	i->1	k->3	l->7	m->1	n->12	q->9	r->29	t->5	u->794	v->7	x->3	
 F	B->1	E->2	M->1	N->11	P->14	R->1	a->2	e->2	i->12	l->19	o->9	r->65	u->1	ä->1	å->2	ö->71	
 G	A->2	U->3	a->17	e->15	i->3	o->18	r->34	u->6	ö->1	
 H	a->50	e->56	i->10	o->4	u->26	ä->5	å->1	
 I	 ->33	-->1	C->3	I->8	M->2	N->4	R->1	S->1	V->3	X->2	l->1	m->3	n->34	r->21	s->40	t->17	z->1	
 J	a->152	e->3	o->19	u->2	ä->1	ö->14	
 K	a->25	f->1	i->36	o->102	u->13	v->2	y->7	ä->4	ö->3	
 L	T->1	a->50	e->15	i->23	l->1	o->17	u->7	y->3	å->12	ö->1	
 M	A->1	a->35	c->6	e->38	i->15	o->38	u->1	ü->1	
 N	a->12	e->11	i->13	o->5	u->1	y->3	ä->14	å->1	
 O	C->1	F->1	L->16	M->1	S->1	b->1	c->5	f->2	i->1	l->3	m->6	n->1	r->1	s->4	u->1	z->2	
 P	P->12	R->1	S->4	V->3	a->70	e->6	l->3	o->38	r->32	u->1	å->5	é->1	
 Q	u->1	
 R	E->2	I->2	a->21	e->13	h->1	i->7	o->18	u->2	y->4	å->6	é->2	
 S	E->4	O->1	P->1	S->1	a->29	c->35	e->16	h->10	i->1	j->6	k->7	l->1	o->19	p->9	r->3	t->27	u->3	v->7	w->3	y->27	á->1	ã->2	å->2	ö->2	
 T	V->4	a->40	e->6	h->23	i->28	o->13	r->4	s->3	u->37	y->20	å->1	
 U	C->2	E->1	N->4	S->11	l->1	n->9	p->1	r->3	t->4	z->2	
 V	 ->1	D->1	I->3	a->27	e->11	i->53	l->1	o->2	ä->7	å->5	
 W	T->1	a->20	e->2	i->11	o->18	u->5	y->4	
 X	 ->1	X->2	
 Y	a->1	o->1	
 Z	e->2	i->1	
 [	K->2	S->1	
 a	 ->3	)->2	b->45	c->58	d->40	f->4	g->47	i->5	j->1	k->81	l->1083	m->39	n->1759	p->12	r->558	s->56	t->6147	u->16	v->3225	x->2	
 b	)->2	a->384	e->2334	i->391	j->2	l->389	o->183	r->317	u->116	y->88	ä->147	å->78	é->1	ö->329	
 c	 ->1	)->1	a->17	e->62	h->26	i->36	o->17	r->1	
 d	)->1	a->422	e->9379	i->476	j->53	o->203	r->153	u->33	v->45	y->23	ä->521	å->172	ö->61	
 e	)->1	-->1	.->1	c->2	d->2	f->487	g->170	j->14	k->261	l->357	m->124	n->3131	p->4	r->381	t->1404	u->391	v->24	x->278	
 f	.->2	a->693	e->117	i->546	j->23	l->217	o->494	r->2386	u->209	y->44	ä->33	å->471	ö->6507	
 g	a->173	e->1084	i->80	j->112	l->99	n->3	o->256	r->627	u->6	y->11	ä->438	å->317	ö->438	
 h	a->2624	e->683	i->146	j->117	o->260	u->289	y->21	ä->571	å->180	ö->230	
 i	 ->3677	,->2	.->6	a->9	b->20	c->34	d->68	f->37	g->57	h->28	k->5	l->19	m->26	n->4011	r->18	s->32	t->37	v->5	
 j	a->1120	e->1	o->76	u->252	ä->73	
 k	a->1129	e->11	i->15	l->223	m->4	n->36	o->3361	r->437	u->464	v->171	y->3	ä->232	ö->26	
 l	'->1	a->427	e->317	i->506	j->13	o->93	u->21	y->108	ä->573	å->183	ö->142	
 m	.->1	a->1029	e->3252	i->1172	j->1	o->498	u->25	y->565	ä->196	å->1110	ö->322	
 n	a->339	e->103	i->316	j->1	o->142	r->29	u->273	y->367	ä->661	å->534	ö->159	
 o	a->50	b->87	c->5149	d->6	e->29	f->195	g->5	h->3	i->7	j->7	k->31	l->216	m->2354	n->25	p->36	r->532	s->344	t->31	u->13	v->16	ä->4	ö->7	
 p	.->1	a->575	e->327	h->2	i->5	l->157	o->522	r->1009	s->1	u->181	y->1	å->2004	
 q	u->4	
 r	a->302	e->1607	i->296	o->83	u->67	y->17	ä->609	å->384	é->1	ö->225	
 s	.->4	a->1008	c->9	e->667	i->1117	j->244	k->1981	l->263	m->82	n->153	o->3645	p->233	r->1	t->2200	u->79	v->197	y->440	ä->1002	å->784	ö->33	
 t	.->26	a->1249	e->152	h->3	i->2856	j->126	o->163	r->618	u->77	v->264	y->306	ä->103	å->8	ö->1	
 u	-->1	l->3	m->1	n->1041	p->1011	r->110	t->1857	
 v	a->1345	e->645	i->3872	o->58	r->7	u->6	ä->619	å->422	ö->1	
 w	a->1	e->1	o->1	
 y	n->2	p->2	r->20	t->134	
 z	i->4	o->4	
 º	 ->1	
 Ä	m->1	n->3	r->3	v->11	
 Å	 ->3	r->1	t->3	
 Î	l->1	
 Ö	V->4	p->1	s->82	
 ä	c->1	g->80	k->1	l->9	m->36	n->649	r->2647	t->1	v->275	
 å	 ->26	b->1	h->1	k->38	l->22	n->1	r->284	s->86	t->657	v->1	
 ö	a->6	b->1	d->13	g->20	k->124	l->1	m->8	n->64	p->98	r->11	s->59	v->673	
! 	1->1	A->6	B->4	C->1	D->56	E->16	F->20	G->5	H->2	I->20	J->112	K->6	L->11	M->7	N->14	O->3	P->6	R->4	S->13	T->13	U->8	V->31	Ä->10	Å->4	Ö->1	
!"	.->1	D->1	J->1	O->1	
!(	P->1	
!.	 ->1	(->1	H->1	
!A	l->2	m->1	n->1	v->1	
!D	e->20	ä->1	
!E	f->2	n->1	r->1	u->1	
!F	r->3	ö->2	
!G	e->1	
!H	a->1	e->9	ä->1	
!I	 ->1	
!J	a->18	
!K	u->1	
!L	e->1	å->1	
!M	e->5	i->2	y->1	ä->1	
!N	i->1	ä->3	
!O	m->2	
!P	r->1	
!R	ö->1	
!S	a->1	k->1	
!T	a->1	i->3	r->1	v->1	
!U	n->1	
!V	i->5	
!Ä	v->2	
" 	(->1	-->1	a->3	b->1	e->1	f->2	g->2	h->1	i->1	m->4	o->6	p->1	s->9	t->2	v->1	Ä->1	ä->1	
"!	I->1	
")	,->1	
",	 ->23	
".	.->1	B->2	D->10	E->2	H->1	I->1	J->5	K->2	N->1	O->2	R->1	V->1	
";	 ->1	
"A	m->1	t->1	
"B	i->1	
"D	e->6	
"E	U->1	q->1	u->2	
"I	 ->1	
"J	a->4	
"K	u->4	v->3	
"L	o->1	
"M	e->1	i->2	
"O	l->1	m->2	
"P	o->1	
"T	i->2	y->1	
"U	r->1	
"a	f->1	l->3	n->3	v->1	
"b	a->1	
"c	o->1	
"d	e->4	i->1	ö->1	
"e	g->1	k->1	n->4	u->3	
"f	o->1	ö->1	
"g	e->2	
"h	e->2	
"i	n->3	r->1	
"j	a->1	
"k	o->2	r->1	u->1	
"l	ä->3	
"m	e->1	
"n	a->1	e->1	o->1	å->1	
"o	b->1	r->1	v->1	
"p	a->1	å->1	
"r	e->5	i->1	
"s	e->1	h->1	k->1	p->1	v->1	
"t	i->1	
"u	t->2	
"v	a->2	
"å	t->1	
"ö	p->1	v->1	
'V	a->1	
'e	a->1	
("	d->1	
(1	4->2	9->13	
(5	7->1	
(8	0->2	
(9	6->1	8->1	9->2	
(A	5->36	p->5	r->1	
(B	5->4	e->1	r->2	
(C	5->7	E->3	N->9	O->15	
(D	A->2	E->3	
(E	G->1	I->1	L->3	N->34	S->1	U->3	
(F	I->2	P->1	R->18	U->1	
(G	e->1	
(H	-->21	o->1	
(I	C->1	F->1	M->1	T->3	h->1	n->1	
(K	O->8	u->2	
(L	i->2	
(N	L->4	
(P	P->1	T->16	a->16	r->1	
(S	E->1	P->1	Y->1	a->4	
(T	a->8	
(U	t->2	
(a	r->7	t->1	v->1	
(d	e->2	
(e	f->1	l->1	n->2	
(f	i->4	o->1	ö->3	
(h	ä->1	
(i	 ->2	n->2	
(k	o->4	r->2	
(m	a->2	e->1	
(o	c->1	
(r	e->1	å->1	
(s	e->1	å->1	
(t	.->1	y->1	
(u	n->1	
(Ö	V->1	s->4	
(å	t->1	
) 	"->1	(->7	-->3	0->3	1->1	3->1	5->3	A->1	B->1	C->1	D->8	E->2	F->9	H->23	I->5	J->16	K->1	L->3	M->1	N->4	O->1	S->1	T->6	U->1	V->5	a->33	b->1	e->1	f->9	h->3	i->9	l->1	m->1	o->13	p->1	s->4	t->1	z->1	Ä->1	ä->2	
)(	G->1	P->9	T->1	
))	 ->5	(->8	.->6	F->1	H->1	o->1	
),	 ->12	
).	 ->1	(->1	)->1	.->4	D->5	F->3	H->5	J->3	K->2	L->1	V->2	
)0	0->3	5->2	6->1	
):	A->19	
);	 ->2	
)?	 ->1	
)A	n->5	
)B	e->8	
)D	e->1	
)F	r->8	ö->2	
)G	e->1	
)H	e->3	
)J	a->3	u->1	
)K	o->1	
)N	ä->3	
)O	l->1	
)R	e->1	
)S	ä->1	
)T	a->1	
)U	t->1	
)]	.->3	
)o	c->1	
)Å	t->1	
, 	"->5	(->1	,->1	1->21	2->9	3->9	4->6	5->3	6->1	7->2	8->2	9->3	A->8	B->9	C->2	D->6	E->18	F->3	G->4	H->4	I->8	J->4	K->7	L->10	M->3	N->2	O->3	P->6	R->5	S->14	T->7	U->1	V->2	W->5	Z->1	a->273	b->123	c->2	d->388	e->319	f->429	g->65	h->291	i->294	j->67	k->212	l->74	m->538	n->172	o->808	p->101	r->57	s->769	t->178	u->209	v->350	y->1	Î->1	ä->185	å->32	ö->11	
,0	7->1	
,2	 ->3	
,3	 ->1	
,4	 ->1	2->1	8->1	
,5	 ->3	
,6	 ->1	
,7	 ->1	
,8	 ->4	
,9	 ->1	
- 	"->1	'->1	(->15	,->1	1->26	2->1	3->1	6->1	8->1	A->2	C->21	D->2	E->1	F->1	H->3	K->2	P->1	R->3	S->2	a->44	b->4	c->1	d->58	e->27	f->24	g->5	h->15	i->28	j->16	k->12	l->5	m->23	n->14	o->171	p->9	r->6	s->54	t->10	u->11	v->23	Ö->2	ä->17	å->2	ö->5	
-(	E->1	
-,	 ->12	
-0	0->39	1->14	2->3	3->12	7->13	8->8	
-1	9->4	
-2	 ->1	-->1	0->22	
-4	 ->1	
-9	8->1	
-A	l->3	r->1	t->1	
-B	e->7	
-C	a->1	l->1	
-D	E->8	e->1	
-E	x->1	
-F	i->3	r->2	
-H	a->1	e->1	
-I	)->1	I->1	s->1	
-J	ø->2	
-K	e->1	
-L	e->1	o->1	
-M	a->3	
-N	o->1	
-P	M->1	l->4	
-R	o->2	
-S	S->1	h->6	y->1	
-a	f->3	l->1	n->7	v->4	
-b	e->7	i->4	r->1	u->2	
-d	a->2	e->3	i->5	o->22	
-e	f->1	l->1	n->1	r->1	
-f	a->1	o->2	r->5	ö->23	
-g	e->2	r->20	
-h	o->1	
-i	n->9	r->1	s->1	
-k	a->4	o->25	r->4	
-l	a->2	e->3	i->2	o->1	ä->5	
-m	a->2	e->7	
-n	a->1	i->1	o->1	y->1	
-o	l->1	m->8	r->4	
-p	o->1	r->27	
-r	a->2	e->7	ä->4	å->4	
-s	h->1	i->1	k->1	o->2	p->3	t->18	y->1	ä->3	
-t	a->9	e->2	r->1	
-u	p->1	t->1	
-v	a->1	ä->1	
-z	o->3	
. 	(->38	-->1	1->20	2->3	7->2	A->2	D->62	E->14	F->8	G->1	H->10	I->5	J->10	K->3	L->1	M->17	N->3	O->6	P->3	R->1	S->7	T->2	U->1	V->17	W->1	a->19	b->1	d->8	e->6	f->10	g->3	h->2	i->11	j->1	k->3	m->8	n->6	o->7	p->3	s->7	t->1	u->2	v->4	Ä->4	Å->1	Ö->1	ä->2	ö->1	
."	 ->1	D->1	I->1	J->1	M->1	
.(	A->6	D->4	E->13	F->6	I->4	L->2	N->4	P->7	S->4	T->7	
.)	 ->4	.->2	A->3	B->8	F->7	G->1	H->2	J->1	O->1	R->1	S->1	Å->1	
.,	 ->3	
.-	 ->15	
..	 ->34	(->25	)->1	.->10	F->1	H->5	L->1	T->1	V->1	
.0	0->13	5->1	
.1	 ->8	)->1	.->3	2->1	4->1	5->1	8->1	9->1	
.2	 ->6	)->1	5->1	
.3	 ->3	,->1	0->1	;->1	
.4	 ->1	.->2	
.5	0->1	5->1	
.8	 ->1	
.9	0->1	
.?	A->1	
.A	c->1	h->1	k->1	l->47	m->2	n->18	r->5	t->23	v->43	
.B	a->6	e->35	i->6	l->7	o->3	r->6	u->1	y->1	ä->1	å->5	
.C	S->1	e->2	o->1	u->1	
.D	E->1	a->7	e->1402	i->8	o->5	ä->121	å->23	
.E	G->3	K->1	U->5	f->41	k->2	m->8	n->101	r->8	t->43	u->51	v->1	x->4	
.F	E->1	P->4	a->9	e->2	i->4	l->7	o->4	r->103	y->1	å->1	ö->234	
.G	e->30	i->2	o->1	r->6	ä->1	å->1	ö->2	
.H	a->27	e->273	i->7	o->4	u->33	y->1	ä->32	ö->1	
.I	 ->221	b->3	d->1	l->1	m->1	n->47	r->1	s->1	t->1	
.J	a->772	o->2	u->10	ä->2	
.K	a->19	i->3	n->1	o->131	r->3	u->7	v->2	ä->6	
.L	a->3	e->3	i->15	y->3	ä->3	å->50	
.M	a->63	e->244	i->48	o->9	y->4	ä->5	å->13	ö->2	
.N	a->17	e->1	i->37	o->1	u->28	y->2	ä->65	å->5	ö->1	
.O	K->1	L->2	M->2	a->2	b->2	c->62	f->3	m->108	n->1	r->17	z->1	
.P	P->2	a->22	e->4	l->4	o->2	r->24	u->2	å->42	
.R	a->4	e->27	i->5	o->3	u->1	ä->3	å->16	
.S	a->31	c->3	e->16	i->5	j->3	k->10	l->38	m->2	n->2	o->48	t->28	u->2	v->1	y->7	ä->4	å->42	
.T	V->1	a->34	e->1	h->3	i->39	o->5	r->22	u->1	v->5	y->17	ä->1	
.U	n->38	p->6	r->4	t->19	
.V	a->89	e->7	i->557	o->1	ä->3	å->26	
.W	o->1	
.Y	t->3	
.a	.->28	
.d	.->3	
.e	x->20	
.g	.->1	
.k	.->4	o->1	
.m	.->8	
.o	.->7	
.Ä	n->24	r->18	v->31	
.Å	 ->13	r->6	t->5	
.Ö	V->1	g->2	k->1	s->2	v->3	
/0	0->7	1->6	2->3	3->6	8->4	
/1	/->2	9->41	
/2	0->26	1->2	
/3	 ->1	5->4	
/4	0->1	3->1	
/5	5->2	9->2	
/6	0->1	
/7	1->2	2->1	5->1	
/9	2->1	5->1	8->2	9->28	
/E	G->8	K->2	u->1	
/N	G->2	o->2	
/O	i->1	
/d	e->1	
/e	l->1	
/h	a->1	
/i	n->1	
/r	i->1	
/s	a->1	
/å	r->2	
0 	-->6	0->11	E->1	a->5	b->2	d->4	e->4	f->8	g->2	h->4	i->10	j->3	k->9	l->1	m->22	n->2	o->8	p->38	r->1	s->5	t->11	u->2	v->1	º->1	ä->12	å->11	
0"	 ->3	.->2	
0(	C->5	
0)	 ->23	.->2	:->1	
0,	 ->13	
0-	 ->1	2->17	b->1	p->4	t->9	
0.	(->2	)->2	2->1	4->1	D->6	F->4	J->2	K->1	M->2	O->1	S->3	T->2	V->1	
0/	1->4	2->3	9->5	
00	 ->76	"->5	)->26	,->7	-->26	.->24	0->141	1->14	2->15	3->7	4->9	5->1	6->31	7->6	8->4	9->4	N->1	
01	 ->1	,->1	/->2	0->14	1->3	2->6	3->1	6->3	8->5	9->2	
02	 ->2	)->2	,->2	.->5	/->1	0->3	1->1	2->3	4->2	
03	 ->2	(->1	/->4	0->1	1->1	2->2	3->4	4->2	5->4	7->4	?->1	
04	 ->1	.->2	/->4	0->1	1->1	5->2	
05	 ->3	(->1	/->4	0->1	5->1	9->2	
06	 ->11	(->2	,->5	.->9	/->5	5->1	6->2	9->1	
07	 ->1	,->1	/->6	1->1	3->1	7->1	8->7	9->5	
08	 ->2	/->5	0->6	1->3	2->3	3->1	7->1	
09	 ->1	/->2	0->1	4->2	5->3	
0N	ä->1	
1 	0->2	4->1	a->1	d->1	e->1	f->3	g->1	i->5	j->11	m->6	o->20	p->7	r->1	s->3	u->3	v->1	ä->2	å->1	ö->1	
1(	C->2	
1)	 ->1	
1,	 ->9	2->2	3->1	4->1	
1-	2->1	o->4	r->5	s->2	
1.	0->4	1->6	3->5	5->1	A->1	E->1	F->1	J->1	K->1	V->1	
1/	1->5	2->3	3->1	9->4	E->3	
10	 ->19	,->1	.->1	/->2	0->9	4->2	5->4	6->3	7->2	8->2	
11	 ->6	,->4	.->6	/->2	0->1	3->1	5->1	
12	 ->9	(->1	,->4	.->7	/->6	0->2	2->1	3->2	4->3	5->1	6->1	7->1	
13	 ->14	(->1	,->2	.->2	/->2	0->1	3->1	8->1	
14	 ->15	,->1	/->1	0->3	3->1	
15	 ->14	,->2	.->2	/->1	0->2	8->4	
16	 ->7	)->1	,->1	4->1	6->1	7->4	9->2	
17	 ->6	,->2	.->2	/->1	0->1	4->1	6->2	
18	 ->9	(->1	,->1	/->3	0->3	
19	 ->6	.->1	/->1	1->1	2->1	3->2	4->5	5->3	6->7	7->2	8->6	9->251	
1:	a->1	
2 	(->1	-->4	0->1	4->1	a->1	b->2	d->2	e->3	f->3	h->1	i->14	j->1	m->6	o->9	p->5	r->1	s->4	u->2	å->1	
2(	C->2	
2)	 ->3	.->1	
2,	 ->23	4->1	5->1	6->1	8->1	
2-	o->3	s->1	
2.	 ->1	0->7	1->1	2->1	D->1	H->1	I->2	J->1	M->3	P->1	V->1	Ä->1	
2/	1->3	2->5	4->1	9->4	
20	 ->19	,->1	.->1	/->2	0->145	1->2	8->2	
21	 ->7	.->2	2->3	:->1	
22	 ->3	,->4	.->1	/->3	6->1	8->1	
23	 ->3	(->1	,->2	
24	 ->5	0->2	4->3	5->1	8->1	
25	 ->13	(->2	.->2	0->1	5->4	
26	 ->7	0->1	2->1	
27	 ->6	(->1	,->1	/->2	
28	 ->4	(->1	,->2	/->1	0->5	:->1	
29	 ->4	,->1	/->1	9->2	
3 	(->2	-->3	0->5	A->1	E->1	a->2	b->1	d->1	f->4	h->2	i->5	j->2	m->1	n->1	o->7	p->9	s->1	u->1	ä->1	
3(	C->3	
3,	 ->6	7->1	8->2	9->1	
3-	1->2	4->1	l->2	
3.	0->1	1->1	2->1	8->1	F->2	I->1	O->1	T->1	
3/	1->4	2->4	7->1	9->2	
30	 ->11	,->2	-->1	0->1	5->1	
31	 ->6	4->1	8->1	
32	 ->1	,->3	.->1	7->2	
33	 ->7	.->1	/->2	2->1	3->2	4->2	
34	 ->4	,->1	.->1	/->2	1->2	4->1	
35	 ->6	.->1	/->4	0->2	1->1	2->2	
36	 ->1	,->1	7->1	
37	 ->3	,->2	.->1	/->1	0->3	1->2	
38	 ->4	,->1	.->1	:->1	
39	 ->3	,->1	
3:	 ->1	
3;	 ->1	
3?	F->1	H->1	
4 	-->1	0->1	c->1	e->3	f->6	h->1	i->8	j->2	l->2	m->5	n->3	o->9	p->5	r->1	s->2	t->4	å->1	
4(	C->2	
4,	 ->8	
4-	0->6	1->1	
4.	1->1	2->1	D->3	F->1	I->3	J->2	K->1	
4/	1->8	2->1	5->2	7->1	
40	 ->13	(->2	,->1	/->1	0->6	9->3	
41	 ->4	/->3	0->1	
42	 ->5	
43	 ->2	.->2	
44	 ->5	.->2	
45	 ->5	,->1	.->5	/->2	
46	 ->2	2->1	
47	 ->1	
48	 ->5	,->1	.->1	7->1	
5 	(->1	-->1	0->5	a->2	c->1	f->3	g->3	h->1	i->6	k->1	m->21	o->10	p->14	r->2	s->3	t->4	v->1	å->3	
5(	C->3	
5)	U->1	
5,	 ->8	5->1	8->1	
5-	0->62	1->1	
5.	 ->1	"->1	)->1	0->2	4->1	D->1	E->1	F->2	H->1	S->1	V->1	
5/	0->1	1->6	2->1	3->1	9->5	E->6	
50	 ->13	,->1	-->3	/->2	0->1	
51	/->1	9->1	
52	 ->2	(->1	/->1	0->2	2->1	
53	 ->1	
54	0->1	
55	 ->6	)->1	/->2	0->1	
56	 ->1	,->1	
57	 ->1	,->1	.->1	1->1	
58	 ->2	)->1	.->1	
59	1->2	8->2	
5b	 ->1	-->1	.->1	
6 	"->1	-->2	0->1	[->1	d->1	e->3	f->4	g->1	h->2	i->11	k->1	l->2	m->2	n->1	o->16	p->7	r->1	s->1	t->2	v->2	ä->1	å->3	
6(	C->2	
6)	 ->1	
6,	 ->12	0->1	
6.	D->3	E->2	F->1	H->1	J->3	M->2	O->1	S->1	T->1	Å->1	
6/	0->2	1->1	2->2	3->3	7->2	9->2	
60	 ->2	-->1	/->2	0->1	
61	4->1	
62	 ->5	.->1	
64	 ->1	
65	2->1	
66	 ->2	2->1	
67	 ->10	,->1	/->1	
68	 ->1	5->1	
69	 ->1	(->2	/->1	
7 	(->2	-->3	0->1	d->5	f->4	g->2	h->3	i->12	l->3	m->8	n->1	o->13	p->7	s->1	t->2	u->1	ä->1	å->1	
7(	C->1	
7)	 ->1	.->1	
7,	 ->15	2->1	4->1	5->1	
7.	-->1	.->1	1->1	2->2	3->1	B->1	D->2	E->1	F->1	I->1	M->1	N->1	S->2	V->2	
7/	0->7	1->6	2->3	6->1	9->3	
70	 ->4	(->2	0->4	
71	 ->1	(->2	/->1	3->1	5->1	
72	8->1	
73	,->1	/->1	
74	 ->1	
75	 ->4	
76	 ->2	2->2	
77	 ->2	8->1	
78	/->2	0->1	1->1	2->1	5->1	6->1	8->1	
79	/->1	1->1	3->1	5->1	6->1	8->1	
7?	D->1	
7N	ä->1	
8 	-->4	4->1	a->1	b->1	d->1	f->4	g->2	h->2	i->7	j->1	k->1	m->7	n->4	o->12	p->1	r->2	s->1	t->4	u->3	v->2	ä->5	
8(	C->1	S->1	
8)	 ->3	.->1	0->1	
8,	 ->10	
8-	2->2	9->1	
8.	 ->1	1->1	4->1	D->1	P->1	S->1	
8/	0->5	1->5	2->2	5->2	9->5	E->1	
80	 ->19	.->1	/->3	1->1	3->1	5->2	7->1	8->1	9->2	
81	 ->6	.->10	/->1	3->1	7->1	9->1	
82	 ->2	)->1	,->5	.->2	/->1	5->2	9->1	
83	 ->2	
85	 ->4	/->2	
86	 ->5	.->1	/->1	
87	 ->1	,->1	.->2	/->1	
88	 ->3	/->3	
89	 ->2	,->1	
8:	 ->1	e->1	
9 	(->1	-->28	a->4	b->1	d->4	e->1	f->7	g->1	h->5	i->7	j->1	k->4	l->1	m->5	n->1	o->8	p->4	r->1	s->2	t->2	u->3	v->3	ä->2	å->1	ö->1	
9"	.->1	
9(	C->2	
9)	 ->19	.->1	0->5	:->18	A->2	
9,	 ->12	
9-	2->2	
9.	 ->1	.->1	1->1	2->2	5->1	D->3	E->2	F->3	J->2	K->1	U->1	V->1	
9/	0->11	1->1	2->4	4->1	9->2	
90	 ->7	(->1	-->1	.->1	
91	 ->4	/->3	7->1	
92	 ->4	,->1	/->1	3->1	
93	 ->5	,->1	-->2	.->1	/->2	0->1	?->1	
94	 ->7	(->2	,->2	-->1	.->1	/->5	5->1	8->1	
95	 ->11	,->2	-->1	.->1	/->5	7->2	
96	 ->11	,->2	.->5	/->6	1->1	7->6	9->1	
97	 ->20	)->1	,->2	.->11	/->8	6->1	7->1	?->1	N->1	
98	 ->22	)->4	,->3	-->3	.->3	/->6	2->2	6->3	9->1	
99	 ->72	"->1	)->45	,->7	-->2	.->17	/->13	0->2	1->3	2->4	3->8	4->6	5->9	6->18	7->42	8->33	9->126	:->1	
9:	 ->1	
: 	"->14	A->6	D->9	E->3	F->11	G->3	H->3	I->4	J->8	K->8	M->1	N->5	O->2	P->3	R->1	S->2	T->2	U->4	V->14	a->12	b->2	d->28	e->10	f->16	g->3	h->7	i->6	j->5	k->4	m->4	n->3	o->5	p->2	r->1	s->2	t->3	u->6	v->22	Ä->2	Å->2	Ö->1	å->1	ö->1	
:A	n->19	
:D	e->2	
:F	ö->2	
:a	 ->1	
:e	 ->3	
:s	 ->74	.->1	
; 	D->1	J->1	a->8	b->1	d->33	e->7	f->10	h->1	i->7	j->4	k->1	l->1	m->5	o->5	p->3	s->3	u->1	v->6	ä->1	å->1	ö->1	
? 	2->1	D->2	H->2	I->1	M->1	O->1	R->1	
?"	J->1	
?,	 ->2	
?-	 ->3	
?.	 ->9	(->2	H->2	
?A	n->4	t->2	v->2	
?B	o->1	
?D	a->1	e->31	ä->3	
?E	f->1	l->1	n->2	t->3	u->2	
?F	i->1	o->1	r->9	ö->8	
?H	a->4	e->16	u->10	ä->2	
?I	 ->8	n->2	
?J	a->23	o->4	
?K	a->5	o->7	ä->1	
?M	a->1	e->3	
?N	a->1	e->6	i->3	ä->4	
?O	c->3	l->1	m->2	
?P	a->1	r->1	å->2	
?R	I->1	e->1	
?S	e->2	k->3	o->2	v->1	
?T	a->1	i->1	y->1	ä->1	
?U	t->1	
?V	a->7	e->3	i->26	
?Ä	r->11	v->2	
A 	-->1	O->1	a->1	e->1	h->3	p->1	v->1	
A)	 ->2	
A,	 ->3	
A-	i->1	s->1	
A.	 ->1	J->1	V->1	
A5	-->36	
A:	s->1	
AB	B->3	C->1	
AD	R->1	
AF	 ->6	,->8	.->4	:->2	
AK	T->1	
AN	D->1	
AR	P->1	
AS	 ->1	P->1	
AT	T->1	
Ac	c->1	t->1	
Ad	a->1	e->1	o->2	r->1	
Af	r->4	
Ag	r->1	u->1	
Ah	e->8	
Ai	d->1	
Ak	k->3	t->1	
Al	a->2	b->4	d->1	e->2	g->1	i->1	l->51	p->2	s->6	t->18	
Am	e->2	o->7	s->39	
An	d->7	g->23	h->1	k->1	l->2	m->1	n->5	s->9	t->3	v->2	
Ap	a->1	p->5	
Ar	a->3	b->4	d->1	i->4	t->3	
As	i->2	s->2	t->1	
At	a->2	l->4	t->29	
Au	s->1	t->1	v->1	
Av	 ->30	b->1	f->1	g->1	i->1	s->17	
Az	o->2	
B 	A->1	o->1	t->1	
B-	A->2	
B5	-->4	
BA	T->1	
BB	 ->1	-->2	
BC	 ->1	
BI	 ->1	
BN	I->7	P->9	
BP	,->1	
BR	Å->1	
BS	E->6	
Ba	k->2	l->8	n->1	r->33	s->3	
Be	d->4	f->1	h->7	k->1	l->9	n->1	r->42	s->5	t->32	v->1	
Bi	g->1	l->5	s->7	
Bl	a->9	o->1	
Bo	e->1	l->1	n->1	r->5	s->1	u->6	w->4	
Br	a->4	e->9	i->5	o->9	u->1	y->19	
Bu	d->2	l->1	s->2	
By	g->1	r->3	
Bä	s->1	
Bå	d->5	
C 	d->1	
C,	 ->1	
C-	l->1	
C.	 ->2	V->1	
C4	-->6	
C5	-->22	
CA	F->1	
CE	C->1	N->12	R->1	S->4	
CH	 ->1	O->3	
CK	 ->1	
CL	A->1	
CM	.->1	
CN	S->9	
CO	D->13	S->2	
CS	U->3	
Ca	d->6	m->2	n->5	r->2	s->2	u->1	v->1	
Ce	n->13	r->1	y->1	
Ch	a->1	i->1	
Cl	a->1	i->1	
Co	c->2	l->1	n->2	r->2	s->9	u->1	x->4	
Cr	e->2	
Cu	n->1	r->1	s->1	x->1	
Cy	p->1	
D 	b->1	f->1	k->1	
D)	)->12	]->1	
D,	 ->1	
D-	g->2	
DA	)->2	
DD	,->1	-->2	R->1	
DE	 ->1	)->4	-->7	B->1	
DR	 ->1	)->1	-->1	.->1	:->1	
DS	K->1	
Da	 ->3	g->8	l->7	m->3	n->26	r->1	v->3	
De	 ->153	l->6	m->2	n->268	r->2	s->61	t->1117	u->1	
Di	m->5	r->9	s->1	
Do	c->2	k->1	m->3	r->1	
Du	b->7	h->1	i->3	t->1	
Dä	r->132	
Då	 ->25	
Dí	e->1	
Dü	h->1	
E 	F->1	h->2	o->2	t->1	ä->1	
E)	 ->3	.->1	J->1	
E-	 ->2	D->8	g->12	k->4	l->1	t->1	
E/	N->2	
EB	A->1	
EC	A->1	H->3	
ED	D->3	
EE	G->3	
EG	 ->7	,->7	-->52	.->1	:->3	?->1	
EI	F->2	
EK	 ->1	(->4	S->8	
EL	)->3	D->3	L->1	
EM	-->1	U->6	
EN	 ->4	)->36	,->2	-->1	:->4	
EO	 ->3	
EP	 ->2	
ER	N->1	R->3	
ES	)->2	-->3	
EU	 ->39	,->5	-->44	.->11	:->44	?->1	G->3	
Ec	e->1	
Ed	i->1	
Ef	f->5	t->50	
Eg	y->2	
Eh	u->2	
Ei	e->1	
Ek	o->5	
El	i->1	l->4	m->2	s->1	
Em	e->8	i->1	
En	 ->67	b->1	d->11	k->1	l->37	
Eq	u->10	
Er	 ->1	a->1	f->2	i->30	k->2	t->2	
Et	i->3	t->48	
Eu	r->851	
Ev	a->7	e->1	
Ex	c->1	e->1	p->2	u->1	x->3	
F 	g->1	h->1	i->2	k->2	s->1	
F)	 ->1	,->1	
F,	 ->8	
F.	A->1	F->1	H->1	M->1	
F:	s->2	
FA	F->1	
FB	I->1	
FE	O->3	
FI	)->1	L->1	P->1	
FJ	)->2	:->1	
FM	I->1	
FN	,->1	-->1	.->1	:->8	
FO	P->1	
FP	Ö->19	
FR	)->18	Å->1	
FS	R->1	
FU	F->1	
Fa	c->4	k->4	r->2	s->1	
Fe	i->2	l->1	m->1	
Fi	n->16	r->1	s->4	
Fl	a->2	e->4	o->19	é->1	
Fo	U->2	g->1	l->6	n->1	r->4	
Fr	a->60	e->1	i->3	u->85	ä->2	å->44	
Fu	n->1	
Fy	r->1	
Fä	s->1	
Få	r->3	
Fö	l->6	r->313	
G 	a->1	o->2	s->1	t->2	u->1	
G(	P->1	
G,	 ->9	
G-	d->24	f->14	i->1	k->16	r->3	
G.	(->1	V->1	
G:	s->3	
G?	,->1	
GA	-->1	S->1	
GF	J->3	
GL	-->2	
GO	R->1	
GU	E->2	S->1	
Ga	l->3	m->3	r->5	z->6	
Ge	m->6	n->41	r->1	
Gi	l->2	n->1	v->2	
Go	e->1	l->13	m->1	n->1	o->1	r->1	t->1	
Gr	a->10	e->14	o->3	u->11	ö->2	
Gu	a->1	i->1	l->1	s->1	t->2	
Gä	l->1	
Gå	 ->1	
Gö	r->2	t->1	
H 	B->1	
H-	0->21	
HO	 ->1	,->1	.->1	
Ha	a->1	d->3	g->1	i->37	m->1	n->25	r->12	t->2	v->1	
He	a->1	b->1	d->2	i->2	l->26	m->1	n->1	r->329	
Hi	c->1	l->1	m->1	s->2	t->12	
Ho	l->3	n->4	p->1	w->1	
Hu	h->1	l->25	r->36	v->7	
Hy	c->1	
Hä	n->4	r->36	
Hå	l->1	
Hö	g->1	
I 	-->4	A->1	E->4	F->2	H->1	I->3	N->1	R->1	S->1	T->3	a->11	b->9	d->86	e->21	f->15	g->3	h->2	i->3	j->1	k->5	l->7	m->10	n->4	o->9	p->5	r->12	s->31	t->1	u->3	v->19	ä->1	ö->3	
I)	 ->2	;->1	
I,	 ->2	
I-	p->3	
I.	 ->2	
I:	e->2	
IC	E->4	
IF	 ->1	)->1	I->1	O->1	
II	 ->7	)->1	,->1	-->2	.->1	:->2	I->5	
IK	,->1	.->2	
IL	,->1	
IM	O->3	
IN	A->3	G->2	T->4	
IP	O->1	
IR	A->1	
IS	P->1	
IT	)->3	
IV	 ->3	
IX	 ->1	,->1	
Ib	l->3	
Id	é->1	
Ih	å->1	
Il	e->1	l->1	
Im	b->3	m->1	
In	d->6	f->4	g->18	i->3	n->2	o->10	r->3	s->2	t->36	
Ir	l->22	
Is	a->2	l->1	r->38	t->1	
It	a->18	
Iz	q->1	
J)	 ->1	,->1	
J:	s->1	
Ja	 ->3	,->8	c->7	g->953	n->1	p->3	v->1	
Je	a->1	r->2	
Jo	 ->1	,->3	n->16	r->4	s->1	
Ju	 ->1	g->1	n->1	s->10	
Jä	m->3	
Jö	r->14	
Jø	r->2	
K 	(->1	n->1	
K(	1->3	9->1	
K,	 ->2	
K.	D->2	
KA	N->1	
KO	M->10	
KS	G->8	
KT	U->1	
Ka	f->1	l->3	n->26	r->12	s->1	t->1	u->4	z->1	
Ke	e->1	
Kf	o->1	
Ki	n->34	r->5	
Kn	a->1	
Ko	c->15	d->1	l->1	m->122	n->22	r->4	s->64	u->12	
Kr	a->3	
Ku	l->25	m->1	n->1	
Kv	a->1	i->5	ä->1	
Ky	o->7	
Kä	n->1	r->10	
Kö	l->2	p->1	
L 	(->1	
L)	 ->7	,->1	
L,	 ->1	
L-	g->2	
LA	 ->1	F->18	S->1	
LD	R->3	
LF	A->1	
LL	A->1	
LT	C->1	
La	 ->2	a->7	m->7	n->35	p->2	
Le	 ->1	a->5	d->5	i->8	o->1	
Li	b->8	i->3	k->13	l->1	s->8	t->2	v->5	
Ll	o->1	
Lo	i->3	m->2	n->4	r->4	t->3	u->1	y->2	
Lu	t->1	x->6	
Ly	c->2	n->4	
Lä	g->2	n->1	
Lå	n->2	t->61	
Lö	ö->1	
M 	A->1	s->1	
M(	1->8	9->2	
M-	2->1	
M.	A->1	
MA	R->1	
MI	 ->1	K->3	
MO	)->1	.->1	:->1	
MR	Ö->2	
MU	,->1	-->2	:->3	
Ma	a->6	c->1	d->6	i->1	j->1	l->7	n->58	r->18	t->2	x->2	
Mc	C->1	N->5	
Me	d->55	l->20	n->214	r->3	x->1	
Mi	c->1	d->2	l->1	n->55	s->2	t->6	
Mo	n->19	r->10	s->1	t->8	u->9	
Mu	l->1	
My	c->1	l->1	n->3	
Mä	n->5	r->1	
Må	h->1	l->2	n->10	
Mö	j->2	
Mü	n->1	
N 	e->1	h->1	k->1	o->1	
N)	 ->37	)->1	
N,	 ->3	
N-	g->1	u->1	
N.	H->1	
N:	s->12	
NA	 ->2	,->1	
ND	E->1	
NG	(->1	.->1	L->2	
NI	 ->6	,->1	F->1	N->2	
NL	)->4	
NM	I->3	
NP	 ->7	,->2	
NS	)->9	
NT	E->4	
Na	l->5	n->1	p->1	r->1	t->27	
Ne	d->9	j->8	w->1	
Ni	 ->45	e->6	k->2	v->1	
No	g->1	i->1	r->7	
Nu	 ->27	m->1	v->1	
Ny	a->3	l->1	t->1	
Nä	r->83	s->26	
Nå	g->5	j->1	
Nö	d->1	
O 	b->2	i->1	ä->1	
O)	.->1	
O,	 ->1	
O.	D->2	
O:	s->1	
O?	E->1	
OC	H->1	
OD	)->13	
OF	S->1	
OK	,->1	
OL	 ->1	)->1	A->18	F->1	
OM	 ->1	(->10	R->2	
OP	)->1	
OR	N->1	
OS	)->2	S->1	
Oa	v->2	
Ob	e->3	
Oc	h->68	k->2	
Of	f->4	t->1	
Oi	l->2	
Ol	i->2	j->3	y->1	
Om	 ->104	a->1	r->15	
On	e->1	ö->1	
Or	a->1	d->11	k->2	o->2	s->2	
Os	l->3	m->1	
Ou	v->1	
Oz	 ->2	,->1	
P 	(->3	a->2	j->1	m->3	o->1	p->4	r->1	å->1	
P)	 ->1	.->1	
P,	 ->3	
PA	-->1	
PE	 ->2	-->13	
PM	 ->1	
PO	L->2	
PP	E->15	
PR	-->1	
PS	E->4	
PT	)->16	
PV	C->3	
Pa	c->3	d->2	k->5	l->26	p->2	r->46	t->23	y->2	
Pe	a->1	i->2	k->1	r->4	t->2	
Pl	a->9	o->1	ä->1	
Po	e->5	h->1	l->2	m->1	n->1	o->1	r->27	w->3	
Pr	e->8	i->1	o->50	í->1	
Pu	n->2	r->1	
PÖ	 ->13	)->2	-->2	:->4	
På	 ->48	s->1	
Pé	t->1	
Qu	e->1	
R 	-->1	a->1	
R)	 ->19	
R-	e->1	g->1	
R.	S->1	
R:	s->1	
RA	 ->1	
RE	G->3	P->2	
RI	N->3	
RN	)->1	ä->1	
RP	O->1	
RR	E->3	
Ra	c->2	f->3	n->4	p->14	s->2	
Re	a->2	d->11	f->7	g->7	n->2	p->1	s->7	t->1	v->4	
Rh	ô->1	
Ri	c->3	i->2	k->5	o->1	s->1	
Ro	b->2	i->1	j->1	m->5	o->1	p->1	t->9	v->2	y->1	
Ru	i->1	m->1	s->1	
Ry	s->4	
RÅ	D->1	G->1	
RÖ	S->2	
Rä	k->1	t->2	
Rå	d->22	
Ré	u->2	
Rö	s->1	
S 	(->1	o->1	
S)	 ->2	)->9	]->2	
S-	z->3	
S:	s->1	
SA	 ->5	,->2	.->2	:->1	
SD	 ->1	
SE	 ->3	)->1	-->7	K->5	M->1	
SG	,->2	-->6	
SK	A->1	
SO	L->1	
SP	 ->2	A->1	Ö->2	
SR	 ->1	
SS	 ->1	:->1	E->1	
ST	N->2	
SU	-->1	:->2	
SY	N->1	
Sa	g->1	i->1	l->1	m->43	n->10	v->9	
Sc	h->38	
Se	a->4	b->1	d->20	g->2	i->5	r->1	t->1	
Sh	a->6	e->10	
Si	m->1	s->2	t->3	
Sj	u->2	ä->3	ö->4	
Sk	a->5	o->6	u->8	y->1	ä->1	
Sl	o->1	u->38	
Sm	å->2	
Sn	a->2	
So	a->1	c->4	k->1	l->6	m->56	u->1	
Sp	a->7	e->2	
Sr	i->3	
St	.->1	a->11	o->21	r->9	ä->1	å->1	ö->11	
Su	a->1	b->2	d->2	
Sv	a->1	e->8	
Sw	o->3	
Sy	d->5	f->6	r->24	
Sá	n->1	
Sã	o->2	
Sä	g->1	k->2	r->2	
Så	 ->34	d->2	l->4	n->1	s->2	v->1	
Sö	d->2	
T 	O->1	
T)	 ->19	
TC	M->1	
TE	 ->1	R->3	
TN	I->2	
TO	?->1	
TT	 ->1	
TU	E->1	
TV	 ->1	-->4	
Ta	 ->1	c->40	d->5	i->1	l->10	m->22	n->5	u->1	
Te	r->4	s->1	x->2	
Th	e->21	y->5	
Ti	b->21	d->2	l->49	t->1	
To	d->1	m->3	n->1	p->2	r->5	t->6	
Tr	a->3	e->2	i->1	o->20	ä->1	
Ts	a->3	
Tu	r->37	s->1	
Tv	ä->4	å->2	
Ty	 ->8	c->1	d->1	s->20	v->9	
Tä	n->2	
Tå	g->1	
U 	"->1	I->1	a->3	b->2	d->1	f->1	g->2	h->2	i->4	k->3	m->3	o->4	p->1	r->1	s->6	u->2	ä->2	
U,	 ->7	
U-	a->1	b->2	e->1	f->6	g->2	i->5	k->7	l->5	m->6	n->1	o->1	p->2	r->3	s->3	t->1	u->1	v->1	
U.	.->1	A->1	D->3	F->1	N->1	R->1	V->3	
U:	s->49	
U?	H->1	
UC	K->1	L->1	
UE	/->2	L->1	N->1	
UF	)->1	
UG	F->3	
UN	I->1	M->3	
US	A->10	D->1	P->1	
Ul	s->1	
Un	d->37	g->3	i->8	
Up	p->7	
Ur	 ->4	b->2	q->1	s->1	
Ut	a->3	b->2	d->1	e->1	f->3	g->2	i->1	m->2	n->2	s->6	t->1	v->3	
Uz	b->2	
V 	-->2	a->1	i->2	
V-	b->1	k->1	p->1	s->1	
VC	,->1	-->1	.->1	
VD	 ->1	
VI	 ->1	I->4	
VP	 ->5	)->1	
Va	d->76	l->9	n->5	p->1	r->30	t->3	
Ve	l->1	m->9	n->4	r->4	t->3	
Vi	 ->558	,->1	a->1	c->1	d->21	k->1	l->30	n->1	s->16	t->10	v->1	
Vl	a->1	
Vo	d->1	l->1	n->1	
Vä	r->4	s->6	
Vå	r->31	
WT	O->1	
Wa	f->2	l->15	s->3	
We	b->1	s->1	
Wi	d->1	e->9	l->1	
Wo	g->18	r->1	
Wu	l->2	r->3	
Wy	e->3	n->1	
X 	o->2	
X,	 ->1	
XV	I->2	
XX	V->2	
YN	)->1	
Ya	s->1	
Yo	r->1	
Yt	t->3	
Ze	e->2	
Zi	m->1	
[K	O->2	
[S	E->1	
].	)->1	H->2	
a 	"->6	(->2	-->63	1->14	2->8	3->4	4->1	5->2	6->2	7->1	8->9	9->1	A->7	B->9	C->9	D->2	E->82	F->15	G->3	H->8	I->5	J->6	K->6	L->7	M->14	N->3	O->1	P->9	R->8	S->7	T->7	U->1	W->1	Z->2	a->1135	b->659	c->22	d->1171	e->937	f->1704	g->443	h->492	i->934	j->41	k->918	l->324	m->1114	n->329	o->1324	p->866	r->718	s->1860	t->705	u->782	v->603	y->19	Ö->6	ä->456	å->226	ö->124	
a!	 ->2	A->1	D->4	F->4	H->2	J->1	L->1	M->1	O->1	Ä->1	
a"	 ->3	,->1	.->7	;->1	i->1	
a)	 ->2	
a,	 ->721	
a-	,->1	I->1	R->1	o->1	
a.	 ->46	(->4	)->2	-->4	.->7	1->1	A->19	B->10	C->1	D->172	E->37	F->36	G->3	H->44	I->42	J->100	K->16	L->9	M->54	N->21	O->22	P->17	R->5	S->26	T->12	U->12	V->101	Ä->11	Å->3	Ö->1	
a/	E->1	h->1	s->1	
a:	 ->31	F->1	
a;	 ->12	
a?	"->1	.->1	A->2	D->8	E->1	F->2	H->3	I->3	J->4	M->1	N->2	P->2	S->1	V->7	Ä->1	
aH	e->1	
aN	ä->2	
aa	f->1	m->1	n->7	r->1	s->6	
ab	 ->1	a->2	b->122	e->51	i->35	l->29	o->13	r->5	s->47	u->4	v->1	
ac	 ->3	"->1	-->1	a->5	c->88	e->21	i->23	k->228	o->3	q->4	t->1	è->1	
ad	 ->641	,->20	-->1	.->50	:->1	;->1	?->3	a->36	d->7	e->1297	g->29	i->52	j->2	k->24	l->11	m->28	o->34	r->7	s->66	t->1	v->8	z->5	ö->1	
ae	l->61	
af	 ->1	a->4	e->1	f->81	i->23	l->1	o->2	r->17	t->187	
ag	 ->2672	,->109	.->106	:->3	;->1	?->4	a->442	b->15	d->12	e->534	f->5	g->29	h->13	i->139	l->35	m->2	n->122	o->71	r->9	s->227	t->125	u->1	å->10	
ah	a->1	u->1	å->43	
ai	 ->7	d->42	l->3	n->38	r->1	v->2	w->1	
aj	 ->5	,->1	.->2	o->43	
ak	 ->52	,->6	.->8	:->1	?->1	a->102	d->1	e->74	f->1	g->31	i->12	k->2	l->13	n->54	o->32	p->1	r->9	s->15	t->555	u->4	ä->1	å->3	
al	 ->290	!->1	"->2	,->24	-->13	.->30	:->2	;->1	F->1	a->679	b->23	d->119	e->173	f->44	i->287	j->35	k->14	l->2023	m->428	n->16	o->33	p->48	r->9	s->58	t->152	u->29	v->29	y->63	ö->1	
am	 ->381	!->1	,->36	.->31	?->2	a->113	b->78	e->739	f->186	g->53	h->170	i->42	k->14	l->97	m->724	n->58	o->115	p->59	r->14	s->62	t->336	u->2	v->9	å->35	ö->86	
an	 ->3158	!->242	"->4	,->247	-->3	.->88	:->7	;->3	?->9	N->1	a->200	b->23	c->9	d->3886	e->155	f->65	g->192	h->112	i->132	j->8	k->201	l->86	m->56	n->245	o->30	p->15	r->6	s->1466	t->598	u->17	v->189	y->3	z->4	ç->1	ö->20	
ao	 ->1	r->1	s->2	
ap	 ->76	"->3	,->16	.->17	:->1	a->358	e->274	i->35	k->11	l->38	n->2	o->2	p->168	r->9	s->92	t->2	
ar	 ->4406	!->24	"->2	)->1	,->215	-->1	.->242	:->13	;->4	?->6	a->1337	b->567	c->3	d->52	e->1039	f->54	g->50	h->27	i->331	j->91	k->346	l->761	m->74	n->574	o->15	p->5	r->16	s->177	t->622	v->30	y->1	z->1	ä->1	å->2	é->1	ó->2	
as	 ->1420	!->4	"->1	,->90	.->140	:->2	;->1	?->2	a->9	b->5	c->16	e->25	h->5	i->41	k->21	m->5	n->3	o->2	p->37	s->78	t->590	u->4	y->21	ä->20	å->4	
at	 ->728	,->55	.->80	:->3	;->1	?->2	a->130	c->2	e->598	f->4	h->6	i->1145	j->1	l->115	n->1	o->77	p->11	r->1	s->424	t->6798	u->216	z->2	ä->1	ö->10	ü->1	
au	 ->9	"->1	,->7	.->1	M->1	b->1	c->1	d->2	e->3	f->1	k->9	m->1	n->4	r->2	s->10	t->11	x->1	
av	 ->2738	,->11	.->13	?->1	a->18	b->14	d->8	e->89	f->26	g->96	h->5	i->14	k->3	l->24	m->1	o->1	p->1	r->5	s->313	t->92	u->1	v->42	
aw	,->1	.->1	
ax	 ->3	-->3	a->2	b->1	e->2	i->17	l->1	
ay	 ->3	,->4	.->1	D->1	a->9	b->1	e->3	s->4	
az	a->7	i->16	
aç	a->5	
b 	S->2	e->1	h->2	k->1	o->3	s->1	v->1	
b)	 ->2	
b,	 ->4	
b-	o->1	
b.	A->1	D->1	
ba	 ->12	-->1	c->4	d->33	g->2	i->1	k->112	l->48	n->105	r->488	s->45	t->184	x->1	y->1	
bb	 ->6	,->2	a->77	e->7	i->1	l->11	p->1	t->43	v->1	y->12	
be	 ->19	a->32	b->3	d->104	f->167	g->180	h->350	i->1	k->152	l->109	m->18	n->15	o->1	r->391	s->543	t->1249	u->3	v->121	x->1	
bi	 ->2	b->13	d->111	e->2	f->5	g->8	h->1	k->2	l->348	n->42	o->10	s->37	t->31	
bj	e->2	u->42	ö->2	
bl	.->27	a->135	e->216	i->349	o->16	u->4	y->8	å->3	
bn	i->1	
bo	 ->3	a->1	c->2	d->3	e->4	g->1	j->1	k->60	l->22	m->10	n->10	r->310	s->14	t->13	u->5	v->2	x->1	
bp	l->1	
br	a->89	e->32	i->114	o->74	u->103	y->24	ä->17	å->23	ö->11	
bs	e->2	i->23	o->41	t->7	u->3	
bt	 ->34	,->3	.->6	
bu	 ->1	d->173	g->1	k->2	l->4	n->28	r->14	s->3	t->2	
bv	a->1	e->12	ä->1	
by	,->1	a->1	b->1	e->1	g->147	i->2	m->1	n->3	r->35	t->20	v->1	x->1	
bä	l->10	n->1	r->145	s->42	t->153	v->10	
bå	d->72	t->9	
bé	 ->1	b->1	
bö	c->3	d->1	j->2	l->1	r->364	t->1	
c 	-->1	B->1	b->2	d->1	i->2	l->1	o->1	s->1	
c"	,->1	
c)	 ->1	
c,	 ->1	
c-	d->1	s->1	t->1	
c.	 ->3	D->1	E->1	
c?	A->1	
cC	a->1	
cN	a->5	
ca	 ->6	,->1	.->1	l->2	n->4	o->1	p->11	s->2	y->6	
cc	e->94	
ce	 ->21	,->1	.->7	d->2	k->2	l->2	m->22	n->243	p->102	r->99	s->114	u->1	
ch	 ->4627	!->1	)->1	,->14	.->2	/->1	:->1	?->1	I->2	a->19	e->43	h->1	i->2	l->4	n->12	o->5	r->18	s->1	t->9	u->3	w->3	y->1	ö->1	ü->4	
ci	a->220	d->1	e->55	f->29	l->3	n->1	o->19	p->209	r->10	s->66	t->24	v->19	
ck	 ->213	"->1	,->28	-->1	.->12	a->308	b->7	d->8	e->664	f->8	h->18	i->1	l->363	n->77	o->40	p->3	r->6	s->637	t->39	u->5	v->3	ö->5	
cl	i->1	
co	,->1	-->1	b->2	m->3	n->3	p->1	r->6	s->5	u->2	v->1	
cq	u->4	
cr	i->1	
ct	.->1	n->1	o->2	
cu	 ->1	,->1	
cy	,->1	a->1	c->1	d->1	f->1	k->7	
cè	t->1	
d 	"->3	(->5	-->11	1->7	2->9	3->2	5->1	7->2	8->2	A->4	B->8	C->1	D->2	E->29	F->5	G->3	H->5	I->5	J->1	K->6	L->8	M->5	O->2	P->2	R->1	S->7	T->4	U->4	V->2	W->1	a->482	b->105	c->2	d->383	e->213	f->292	g->102	h->110	i->166	j->24	k->135	l->28	m->222	n->67	o->221	p->111	r->64	s->367	t->211	u->69	v->136	y->8	Ö->2	ä->63	å->17	ö->39	
d!	 ->2	
d)	 ->1	,->3	
d,	 ->166	
d-	 ->1	a->1	f->1	k->1	
d.	 ->3	"->2	(->1	,->1	-->1	.->2	A->4	B->1	D->55	E->6	F->8	G->1	H->16	I->10	J->23	K->7	L->2	M->13	N->7	O->18	P->2	R->3	S->5	T->3	U->4	V->16	Ä->2	Å->3	
d:	 ->4	
d;	 ->5	
d?	 ->1	-->2	.->1	D->1	F->1	H->1	J->1	V->1	Ä->1	
da	 ->683	!->1	"->1	,->39	.->38	?->4	b->2	c->5	d->40	f->3	g->372	h->43	i->1	k->6	l->15	m->264	n->741	p->1	r->247	s->144	t->123	
db	a->9	e->20	o->170	r->58	u->1	ä->10	
dd	 ->69	)->1	,->4	.->8	a->86	e->134	h->1	i->5	n->4	s->17	
de	 ->4583	!->9	"->1	(->1	,->172	-->5	.->211	:->39	;->5	?->7	H->1	P->1	a->7	b->181	c->41	d->2	e->4	f->58	g->5	h->1	i->2	k->15	l->959	m->356	n->3369	o->5	p->9	r->2020	s->847	t->4843	u->3	v->8	z->3	
df	i->3	r->10	u->1	ä->4	ö->249	
dg	a->67	e->127	i->28	n->71	o->1	r->2	ä->2	å->5	ö->3	
dh	e->25	i->1	j->1	å->4	ö->1	
di	 ->20	,->1	.->3	:->1	;->1	a->60	c->3	d->14	e->32	f->10	g->701	k->40	l->3	m->13	n->18	o->9	p->11	r->251	s->252	t->40	u->4	v->18	z->5	ä->1	
dj	a->91	e->83	o->1	u->58	ä->9	
dk	a->1	o->25	u->3	v->1	ä->94	
dl	a->182	e->356	i->395	ä->79	ö->1	
dm	a->1	e->4	i->28	o->4	ä->1	å->3	
dn	a->38	i->408	
do	 ->5	,->1	.->4	c->61	e->1	f->1	g->15	k->45	l->11	m->186	n->70	r->39	s->7	u->1	v->4	x->6	ä->1	
dp	e->1	o->1	r->1	u->119	
dr	a->1121	e->72	i->420	o->19	u->6	y->4	ä->40	å->1	ö->9	
ds	 ->102	,->4	-->6	.->5	/->1	;->1	N->1	a->41	b->56	c->1	d->19	e->23	f->24	g->1	h->6	i->9	j->1	k->89	l->20	m->33	n->8	o->31	p->64	r->16	s->39	t->20	u->5	v->5	y->5	ä->1	å->3	ö->1	
dt	 ->8	,->4	a->108	e->15	i->1	o->4	y->7	
du	 ->6	a->1	b->17	c->35	e->8	g->7	k->55	m->8	n->2	p->4	r->1	s->115	t->2	
dv	a->26	e->61	i->44	o->5	r->13	s->45	u->1	ä->129	
dw	i->1	
dy	k->7	l->3	n->5	r->8	s->1	
dz	i->4	j->5	
dä	c->1	m->2	r->523	
då	 ->204	,->3	.->2	?->1	l->19	t->6	v->1	
dé	 ->10	,->1	e->9	n->15	
dö	 ->1	d->21	e->1	l->10	m->90	p->4	r->14	s->1	t->3	v->1	
e 	"->9	(->37	-->43	1->17	2->8	3->1	4->3	8->1	9->1	A->6	B->7	C->3	D->4	E->29	F->6	G->7	H->4	I->4	J->2	K->8	L->2	M->5	N->2	O->3	P->23	Q->1	R->6	S->6	T->2	V->2	W->1	a->759	b->457	c->11	d->436	e->392	f->878	g->278	h->420	i->511	j->94	k->557	l->212	m->607	n->254	o->605	p->447	q->2	r->321	s->943	t->478	u->273	v->538	y->14	Ö->1	ä->264	å->136	ö->99	
e!	 ->7	A->1	D->1	J->1	M->1	N->1	S->1	Ä->1	
e"	 ->2	,->3	
e(	A->1	
e)	 ->3	
e,	 ->370	
e-	 ->7	A->3	F->2	L->2	M->1	N->1	a->4	d->5	f->3	l->2	m->2	p->2	s->14	
e.	 ->12	-->2	.->5	A->9	B->3	D->93	E->19	F->21	G->3	H->21	I->13	J->60	K->9	L->8	M->35	N->9	O->11	P->7	R->5	S->20	T->13	U->4	V->36	d->1	Ä->5	Å->4	Ö->1	
e:	 ->46	
e;	 ->6	
e?	D->2	E->1	F->2	H->6	I->1	J->1	K->1	O->1	S->1	V->2	
eE	n->1	
eF	r->1	
eH	e->1	
eN	ä->2	
eP	r->1	
ea	 ->4	d->8	g->16	k->54	l->23	m->8	n->2	r->4	t->30	u->6	
eb	,->1	a->175	b->2	e->21	i->1	o->8	r->21	u->9	y->25	ä->119	å->1	ö->8	
ec	 ->1	e->42	i->135	k->339	o->1	t->1	u->2	y->1	
ed	 ->1610	,->15	.->14	a->598	b->187	d->126	e->389	f->22	g->27	h->1	i->35	j->77	k->6	l->378	m->3	n->83	o->31	r->227	s->84	t->18	u->5	v->74	ö->55	
ee	-->2	.->1	l->8	n->68	r->17	s->1	x->1	
ef	 ->1	a->39	e->24	f->149	i->83	l->8	o->226	r->25	t->373	u->20	ä->22	ö->23	
eg	 ->56	,->3	.->2	a->136	d->1	e->616	i->366	l->151	n->46	o->14	r->152	u->1	ä->60	å->30	
eh	a->95	i->1	o->67	r->7	ä->1	å->120	ö->171	
ei	d->2	j->2	k->5	l->1	n->16	r->5	s->715	v->1	x->5	z->1	
ej	 ->13	,->10	.->4	d->4	o->3	u->4	ä->3	
ek	 ->3	a->122	e->10	h->4	i->9	l->62	n->52	o->395	r->48	s->6	t->793	u->7	v->86	y->16	ä->42	
el	 ->494	!->4	,->54	-->11	.->45	:->5	;->1	?->2	a->422	b->38	e->133	f->6	g->20	h->33	i->66	k->3	l->1282	m->6	n->63	o->24	p->4	r->12	s->764	t->265	u->3	v->68	y->4	z->1	ä->36	ö->6	
em	 ->355	,->35	.->68	:->5	;->2	?->2	a->52	b->55	e->647	f->1	h->14	i->43	l->17	m->27	o->258	p->125	s->334	t->28	v->1	y->1	ä->43	å->20	ö->15	
en	 ->10552	!->7	"->12	)->11	,->715	-->1	.->907	:->25	;->17	?->32	F->3	H->2	I->1	J->2	N->5	a->377	b->76	c->1	d->588	e->191	f->9	g->100	h->228	i->110	j->2	k->58	l->135	n->637	o->485	p->1	r->5	s->2065	t->1674	u->7	v->14	z->19	Ä->1	ä->3	å->1	è->3	ö->3	
eo	g->8	l->5	m->3	n->3	r->3	s->2	t->1	
ep	 ->2	a->67	e->1	h->3	n->1	o->12	p->33	r->28	s->2	t->126	u->19	
er	 ->6908	!->85	"->7	)->9	,->476	-->15	.->508	:->19	;->7	?->16	H->1	J->1	M->1	N->2	a->1780	b->70	c->1	d->66	e->381	f->110	g->197	h->324	i->1028	k->645	l->213	m->33	n->1708	o->104	p->8	r->729	s->743	t->292	u->39	v->187	y->2	ä->57	å->13	ö->52	
es	 ->403	"->1	,->17	-->7	.->17	;->1	a->35	b->2	d->2	e->67	f->6	g->5	h->4	i->31	k->185	l->353	m->15	n->4	o->105	p->111	q->1	r->3	s->835	t->428	u->173	v->35	y->2	ä->6	ö->11	
et	 ->7761	!->6	"->9	)->14	,->512	-->2	.->565	:->13	;->6	?->25	J->1	a->594	b->1	c->6	d->1	e->1198	f->11	h->1	i->14	j->1	k->17	l->36	m->2	n->31	o->78	p->14	r->196	s->812	t->2596	u->11	v->30	y->131	ä->299	å->10	ê->2	ö->1	
eu	g->2	m->1	n->3	r->416	s->1	t->12	
ev	 ->25	.->1	a->67	d->2	e->45	i->140	l->4	n->12	o->1	s->6	t->4	ä->17	å->2	
ew	 ->1	i->1	o->2	
ex	 ->24	,->1	.->21	a->39	c->5	e->117	i->50	k->3	m->1	p->60	t->90	u->3	v->1	
ey	 ->3	e->3	h->1	
ez	 ->4	,->2	-->2	u->1	
eä	g->2	
eå	t->1	
f 	-->1	H->2	a->1	e->2	f->5	h->3	i->3	k->1	l->1	n->1	o->5	s->4	t->1	u->1	ä->1	
f,	 ->5	
f-	 ->2	M->2	
f.	D->2	E->1	J->1	d->2	
fa	 ->25	,->2	.->1	b->2	c->4	d->11	e->3	i->1	k->136	l->251	m->15	n->72	r->419	s->138	t->268	u->1	v->1	x->1	
fb	e->1	
fd	r->1	
fe	b->16	d->12	k->162	l->39	m->57	n->114	r->249	s->9	t->1	
ff	 ->3	,->1	-->2	a->145	b->1	e->257	i->7	l->3	p->2	r->66	ä->12	
fh	j->1	
fi	 ->3	,->1	.->2	c->74	d->2	e->61	k->41	l->12	n->566	q->1	r->3	s->61	t->5	
fj	o->13	ä->11	
fk	r->1	
fl	a->34	e->158	i->22	o->9	u->14	y->61	ä->2	ö->4	
fm	a->1	
fo	b->1	d->10	g->58	k->5	l->122	n->128	r->725	s->4	t->4	
fp	r->2	
fr	a->732	e->116	i->222	o->23	u->87	y->5	ä->173	å->1433	
fs	i->1	t->6	
ft	 ->102	!->1	,->13	.->14	:->1	?->2	a->146	b->1	e->588	f->12	i->49	l->8	n->113	o->5	s->21	t->5	v->8	
fu	l->150	n->116	s->10	t->1	
fy	l->62	r->28	s->9	
fä	d->1	k->1	l->121	n->2	r->67	s->25	
få	 ->206	,->3	.->3	g->9	n->14	r->186	s->1	t->58	
fé	r->1	
fö	d->9	g->2	l->165	n->1	r->8138	t->3	
g 	(->6	-->25	1->22	2->9	3->6	4->8	5->2	6->4	8->2	D->1	E->3	F->1	G->1	H->14	I->4	O->1	T->1	V->1	[->1	a->714	b->145	c->2	d->111	e->117	f->463	g->93	h->286	i->379	j->11	k->199	l->58	m->250	n->77	o->394	p->163	r->94	s->636	t->482	u->147	v->405	y->2	Ö->2	ä->187	å->39	ö->28	
g!	"->1	H->1	J->1	
g"	 ->3	,->2	.->3	
g)	 ->4	,->1	.->1	N->1	
g,	 ->416	
g-	P->1	
g.	 ->10	(->2	)->3	.->4	A->13	B->4	D->115	E->18	F->29	G->5	H->27	I->23	J->63	K->15	L->6	M->25	N->12	O->23	P->7	R->3	S->12	T->7	U->2	V->37	a->1	Ä->4	
g:	 ->9	D->2	
g;	 ->8	
g?	D->5	F->3	H->2	J->2	O->1	T->1	V->1	Ä->1	
gN	ä->1	
ga	 ->1833	!->6	,->91	.->86	/->1	:->11	;->1	?->3	d->67	g->35	k->1	l->54	m->34	n->762	p->1	r->1360	s->142	t->97	u->18	v->21	
gb	a->15	e->1	l->1	o->1	r->1	y->1	
gd	 ->29	,->1	.->2	a->9	e->46	o->27	p->4	r->2	s->10	y->1	
ge	 ->210	,->4	.->6	?->1	d->6	f->10	k->1	l->112	m->399	n->2476	o->10	r->1013	s->50	t->474	
gf	a->15	l->1	o->21	r->2	u->1	ä->2	ö->5	
gg	 ->31	"->1	,->8	.->6	;->1	a->273	b->1	d->4	e->149	h->6	i->3	j->13	l->1	n->47	o->2	r->14	s->24	t->5	å->2	ö->21	
gh	 ->2	.->1	e->851	t->3	å->2	
gi	 ->34	,->6	-->1	.->10	a->7	b->3	c->23	e->35	f->106	g->10	i->1	k->47	l->28	m->5	n->22	o->254	p->8	s->169	t->149	u->3	v->122	z->5	ä->1	å->1	ö->4	
gj	o->136	
gk	r->3	u->1	ö->1	
gl	a->62	e->134	i->89	j->1	o->12	u->1	ä->41	ö->21	
gm	 ->1	a->4	e->6	ä->3	å->1	
gn	 ->4	a->182	e->16	i->229	o->4	u->2	ä->1	
go	 ->3	d->238	f->1	g->5	i->2	l->6	m->8	n->226	r->355	s->2	t->214	u->1	
gp	l->4	o->2	
gr	a->617	e->160	i->72	o->5	u->482	y->1	ä->142	å->2	ö->21	
gs	 ->99	,->5	-->12	.->3	a->42	b->37	c->13	d->5	e->16	f->329	g->16	h->3	i->23	j->2	k->197	l->76	m->29	n->16	o->14	p->110	r->44	s->99	t->191	u->8	v->46	y->2	ä->8	å->6	ö->1	
gt	 ->1229	!->2	,->73	.->83	:->1	;->1	?->1	a->1	e->12	g->11	i->8	o->5	r->2	s->39	v->112	
gu	d->2	e->5	l->2	m->18	r->1	s->1	v->1	
gv	a->7	e->1	
gy	n->19	p->2	
gä	c->1	l->406	n->24	r->338	v->1	
gå	 ->94	.->7	e->101	n->259	r->160	s->6	t->36	v->2	
gö	m->4	r->622	
h 	"->3	(->1	-->6	0->1	1->21	2->13	3->7	4->10	5->3	6->2	7->6	8->11	9->4	A->4	B->6	C->4	D->4	E->36	F->15	G->7	H->3	I->14	J->2	K->9	L->8	M->5	N->2	O->2	P->17	R->3	S->27	T->8	U->1	V->2	W->1	X->1	a->292	b->119	c->10	d->609	e->212	f->321	g->92	h->164	i->234	j->162	k->198	l->94	m->280	n->85	o->99	p->115	r->188	s->448	t->153	u->106	v->237	y->7	Ö->7	ä->55	å->37	ö->43	
h!	 ->1	
h)	D->1	
h,	 ->16	
h-	B->7	a->1	
h.	D->1	E->1	F->1	J->1	V->1	
h/	e->1	
h:	 ->1	
h?	F->1	
hI	 ->1	I->1	
ha	 ->190	,->1	.->1	b->2	d->85	f->37	g->2	k->1	l->27	m->43	n->808	p->2	r->1722	s->5	t->5	u->1	v->54	
he	 ->5	,->1	a->22	b->1	c->1	d->8	e->14	f->17	i->5	j->2	k->2	l->393	m->42	n->49	p->3	r->231	s->1	t->1789	u->2	z->1	
hh	o->1	
hi	e->7	g->1	l->1	n->91	p->1	q->1	s->36	t->63	
hj	a->1	ä->135	
hl	e->4	
hn	e->13	
ho	 ->4	.->1	b->2	c->6	e->1	f->1	k->1	l->8	m->7	n->57	p->125	r->6	s->51	t->40	v->80	w->1	
hr	e->10	k->1	o->14	ö->1	
hs	 ->1	
ht	 ->4	.->1	a->1	e->2	f->3	i->1	s->1	
hu	 ->1	d->2	g->3	l->4	m->9	n->21	r->212	s->27	v->47	
hw	a->1	e->1	i->1	
hy	 ->1	c->5	g->2	l->2	p->2	r->2	s->14	
hä	f->2	l->119	m->14	n->226	r->308	s->1	v->39	
hå	g->18	l->477	n->2	r->29	v->1	
hô	n->1	
hö	g->143	j->23	l->18	n->1	r->129	s->1	v->148	
hü	s->4	
i 	"->1	-->11	1->16	2->13	5->1	8->2	A->29	B->30	C->9	D->14	E->203	F->30	G->13	H->15	I->22	J->1	K->45	L->34	M->26	N->6	O->2	P->13	R->4	S->40	T->41	U->5	V->4	W->5	Y->1	a->338	b->243	c->3	d->794	e->315	f->528	g->134	h->402	i->253	j->32	k->332	l->83	m->372	n->88	o->163	p->128	r->147	s->687	t->152	u->136	v->341	y->5	z->2	Ö->38	ä->107	å->25	ö->35	
i!	 ->3	H->1	J->1	
i"	 ->1	
i,	 ->84	
i-	 ->10	,->1	g->1	i->1	r->1	
i.	(->1	.->2	A->3	B->1	D->12	E->4	F->4	H->4	I->1	J->3	K->2	L->1	M->3	N->1	S->3	U->1	V->6	
i:	 ->1	
i;	 ->1	
i?	 ->1	.->1	
ia	 ->51	,->4	-->1	.->2	g->1	k->8	l->279	n->19	r->21	s->7	t->88	
ib	a->7	b->1	e->95	i->12	l->33	u->1	y->1	
ic	 ->3	a->3	e->85	h->12	i->15	k->141	y->4	
id	 ->441	,->19	.->18	:->1	a->236	d->21	e->264	g->109	h->5	i->227	k->1	l->7	m->1	n->23	o->11	p->10	r->115	s->66	t->70	u->10	é->33	
ie	 ->4	,->1	-->2	b->3	c->1	d->4	f->8	k->1	l->137	m->3	n->182	p->1	r->267	s->7	t->91	u->1	ä->2	
if	a->10	e->7	f->27	i->102	o->4	r->61	t->266	u->1	ö->4	
ig	 ->1066	!->2	"->1	,->50	.->55	:->3	;->1	?->4	a->1254	d->12	e->597	g->144	h->836	i->9	j->1	l->5	m->1	n->21	o->6	r->13	s->4	t->1337	v->1	å->13	ö->6	
ih	a->3	e->116	j->1	o->12	ä->1	å->16	
ii	k->3	m->1	n->2	s->2	
ij	-->1	s->2	
ik	 ->155	!->1	"->1	,->35	-->2	.->34	:->1	?->2	a->403	e->485	g->2	h->39	i->57	l->22	m->2	n->66	o->12	r->17	s->58	t->914	v->9	ä->37	
il	 ->28	,->2	-->5	.->6	a->108	b->4	d->175	e->18	f->2	h->1	i->84	j->536	k->345	l->3466	m->3	o->16	p->7	r->2	s->16	t->180	u->1	v->9	ä->2	å->1	ö->1	
im	a->38	b->1	e->27	i->72	l->23	m->21	o->1	p->18	s->9	t->4	u->18	y->1	å->1	ö->1	
in	 ->550	!->1	"->1	,->31	-->3	.->33	:->1	?->1	a->360	b->36	c->203	d->336	e->98	f->290	g->4451	h->14	i->255	j->93	k->57	l->111	m->1	n->929	o->322	p->1	r->213	s->600	t->1989	u->24	v->76	z->2	ä->12	ö->1	
io	 ->40	,->3	-->4	.->2	:->1	;->1	d->86	e->4	f->2	g->1	l->7	n->3256	p->4	r->42	s->6	t->12	x->7	
ip	 ->29	,->3	.->4	a->42	e->172	i->10	l->32	n->10	o->5	p->5	r->7	s->2	
iq	u->4	
ir	 ->112	,->2	:->1	a->12	e->272	g->5	i->1	k->13	l->11	m->2	o->2	r->22	t->1	
is	 ->330	!->1	)->1	,->22	-->5	.->16	:->1	;->1	?->1	a->283	b->18	c->26	d->8	e->254	f->4	h->4	i->99	k->2383	l->2	m->104	n->16	o->16	p->5	r->20	s->1482	t->639	u->4	v->1	y->1	ä->11	
it	 ->309	,->8	-->5	.->10	a->107	b->53	e->415	h->1	i->874	l->15	n->1	o->25	r->9	s->63	t->389	u->312	y->5	z->2	ä->7	
iu	m->27	t->1	
iv	 ->229	,->27	.->29	:->2	;->1	?->2	a->284	b->2	e->307	f->4	i->146	k->3	l->15	n->20	r->6	s->119	t->125	ä->3	å->111	
iw	a->1	
ix	.->1	a->5	e->1	t->1	
iz	 ->4	,->2	-->1	i->5	
iä	k->1	r->17	
iå	l->1	t->1	
iè	r->1	
ié	 ->1	
iö	s->24	
j 	1->3	2->1	L->1	a->3	b->3	f->3	i->1	k->1	l->2	m->1	n->1	o->1	t->1	ä->1	ö->1	
j,	 ->13	
j-	v->1	
j.	(->1	D->1	E->1	I->1	J->1	R->1	T->1	V->1	
ja	 ->444	,->11	.->8	d->18	g->1088	k->24	l->7	m->1	n->129	p->1	r->71	s->35	t->23	
jd	 ->25	.->1	a->12	e->28	o->1	p->2	r->1	s->2	å->1	
je	 ->169	,->4	-->1	.->2	:->1	b->15	d->7	f->3	i->3	j->3	k->70	l->11	m->1	n->4	r->149	s->2	t->15	u->2	v->3	å->1	
jf	l->1	
ji	k->5	
jk	a->1	o->3	
jl	i->309	
jn	i->19	
jo	b->4	c->2	l->4	n->66	r->262	s->1	u->3	v->17	
js	 ->6	,->1	.->1	m->2	
jt	 ->5	s->4	
ju	 ->78	,->3	a->1	b->1	d->52	g->5	k->17	l->13	n->29	p->39	r->64	s->121	t->35	v->2	
jä	l->286	m->71	n->173	r->66	t->21	v->2	
jö	 ->8	!->1	,->11	-->2	.->6	a->4	b->4	d->4	e->4	f->18	i->1	k->26	l->1	m->17	n->44	o->5	p->14	r->5	s->32	t->1	u->1	v->10	
k 	-->6	D->1	J->1	K->1	T->1	a->59	b->32	c->2	d->23	e->21	f->76	g->17	h->30	i->62	j->11	k->55	l->21	m->48	n->29	o->95	p->46	r->24	s->125	t->38	u->32	v->35	ä->14	å->16	ö->5	
k!	A->1	O->1	
k"	 ->3	
k,	 ->101	
k-	 ->3	b->1	d->1	f->1	i->1	p->1	s->1	
k.	 ->7	.->1	A->3	B->2	D->23	E->3	F->6	G->1	H->12	I->4	J->7	K->2	M->3	N->1	O->2	R->2	S->1	T->4	V->10	Ä->2	
k:	 ->2	
k?	H->1	N->1	R->1	V->1	
ka	 ->2418	"->1	,->44	-->1	.->35	:->2	?->2	b->7	d->169	f->27	g->4	k->2	l->794	m->99	n->1377	o->2	p->705	r->354	s->161	t->301	v->4	y->11	
kb	a->12	e->8	i->1	o->1	ä->1	
kd	a->1	e->8	o->1	ö->1	
ke	 ->231	!->1	)->2	,->24	-->19	.->27	:->1	E->1	F->1	N->1	b->1	d->29	f->2	g->1	k->1	l->176	m->15	n->393	o->2	p->19	r->706	s->71	t->790	v->2	
kf	a->8	o->1	r->3	y->1	ö->11	
kg	i->2	r->33	
kh	 ->1	-->1	.->2	a->6	e->55	o->3	u->7	ä->9	
ki	 ->2	.->1	c->17	d->1	e->38	f->6	g->5	l->265	n->22	p->12	r->1	s->88	t->7	v->2	
kj	u->31	
kk	a->1	i->2	o->2	u->4	ö->1	
kl	.->21	a->542	e->7	i->578	o->10	u->25	y->6	ä->1	ö->1	
km	 ->2	,->1	.->1	e->4	o->1	
kn	a->342	e->3	i->403	o->4	u->8	y->9	ä->2	
ko	 ->5	,->1	.->1	a->14	d->15	e->1	f->5	g->40	h->5	k->2	l->272	m->2390	n->1344	o->1	p->17	r->331	s->122	t->179	u->1	v->3	
kp	a->10	r->4	
kr	a->472	e->105	i->358	o->59	y->9	ä->216	å->2	ö->1	
ks	 ->39	,->1	.->5	;->1	a->131	b->2	c->2	d->3	e->2	f->4	i->3	k->1	l->2	o->60	p->9	r->4	s->6	t->25	v->1	w->1	ä->1	å->587	ö->1	
kt	 ->773	!->1	"->1	,->47	.->69	:->4	;->2	?->3	a->236	b->7	d->2	e->495	f->3	h->3	i->1135	k->1	l->95	m->3	n->55	o->145	p->2	r->13	s->23	t->8	u->257	y->9	ä->9	ö->23	
ku	b->2	g->3	l->641	m->48	n->326	p->6	r->304	s->98	t->85	u->2	y->2	
kv	a->102	e->65	i->66	o->16	ä->50	å->3	
ky	 ->1	d->109	f->1	h->1	l->37	m->17	n->15	r->1	v->1	
kä	l->100	m->51	n->265	r->127	
kå	d->10	l->1	r->1	t->3	
kö	k->1	l->5	n->10	p->11	r->17	t->29	v->1	y->1	
l 	"->1	(->3	-->14	1->38	2->28	3->10	4->10	5->9	6->13	7->12	8->18	9->7	A->1	B->6	C->3	D->2	E->35	F->7	G->2	H->2	I->3	K->17	L->2	M->4	N->3	O->1	P->7	R->2	S->8	T->5	U->1	V->1	W->4	a->545	b->187	c->5	d->360	e->235	f->350	g->132	h->144	i->191	j->118	k->186	l->53	m->152	n->81	o->232	p->108	r->103	s->436	t->136	u->107	v->184	y->5	Ö->1	ä->71	å->29	ö->31	
l!	 ->2	H->2	J->1	M->1	T->1	
l"	 ->2	,->2	.->1	
l'	e->1	
l,	 ->183	
l-	 ->18	2->1	D->1	F->3	H->1	I->2	R->1	S->7	f->1	p->1	s->2	
l.	 ->24	1->1	A->3	B->3	D->47	E->10	F->15	G->1	H->11	I->10	J->22	K->7	L->1	M->12	N->4	O->2	P->3	R->1	S->13	T->4	U->1	V->25	a->27	Ä->4	
l:	 ->12	
l;	 ->3	
l?	.->1	D->1	E->1	H->1	J->2	K->1	
lF	i->1	
la	 ->1598	!->1	"->5	,->24	.->29	:->1	?->4	a->1	b->3	c->32	d->138	f->1	g->1037	i->7	k->26	m->614	n->1096	p->8	r->817	s->172	t->188	u->9	v->7	w->2	y->3	
lb	a->119	e->13	i->1	l->1	o->3	r->7	u->15	y->1	
ld	 ->43	,->10	.->5	a->111	b->2	e->163	g->1	h->23	i->77	j->1	n->66	o->1	r->49	s->23	t->2	
le	 ->538	,->3	-->2	.->2	d->439	f->2	g->268	h->3	i->2	j->2	k->45	l->17	m->555	n->287	o->1	r->1455	s->105	t->342	u->4	v->91	w->2	x->33	z->1	
lf	 ->2	-->2	a->1	e->6	i->1	k->1	o->24	r->41	s->3	t->4	u->3	ä->106	å->4	ö->42	
lg	a->2	e->3	i->18	j->1	o->1	r->4	ä->21	å->26	ö->2	
lh	a->47	e->25	j->8	o->1	ö->8	
li	 ->138	!->1	,->3	.->1	a->8	b->33	c->52	d->46	e->45	f->15	g->2866	h->1	k->426	l->6	m->25	n->639	o->2	p->2	r->117	s->279	t->763	v->193	x->1	
lj	 ->3	,->2	.->1	a->377	d->44	e->112	f->1	k->2	n->13	o->65	s->5	t->5	u->14	ö->190	
lk	 ->14	,->1	.->8	a->132	e->257	f->1	g->2	h->9	l->5	n->57	o->135	p->10	r->10	s->6	u->1	v->3	y->1	ä->12	ö->2	
ll	 ->3368	!->2	"->3	,->71	-->4	.->86	:->3	?->5	a->1441	b->87	d->118	e->2158	f->153	g->52	h->54	i->137	k->87	m->138	n->192	o->53	p->1	r->99	s->275	t->597	u->15	v->195	y->6	ä->199	å->59	ö->2	
lm	 ->1	,->1	.->1	a->432	e->7	o->1	s->1	y->2	ä->131	å->2	ö->6	
ln	 ->19	,->2	.->1	a->46	i->213	s->2	ä->6	
lo	 ->9	,->3	a->1	b->22	c->10	d->5	g->99	j->7	k->53	l->2	m->20	n->4	o->1	p->21	r->93	s->15	t->16	v->24	y->1	
lp	 ->48	,->2	.->5	a->49	e->8	l->2	o->45	r->4	s->1	t->3	u->2	v->1	
lr	a->11	e->15	i->7	o->1	u->1	y->1	ä->88	
ls	 ->145	,->4	-->1	.->10	?->1	a->64	b->2	d->2	e->441	f->8	h->3	i->26	k->58	l->10	m->16	n->3	o->20	p->15	r->5	s->53	t->190	u->5	v->7	y->9	ä->124	ö->6	
lt	 ->745	,->24	.->28	:->1	;->2	?->1	a->186	b->1	e->78	f->40	h->8	i->141	j->3	m->1	n->48	o->3	r->12	s->83	u->146	ä->4	
lu	c->5	d->6	f->3	g->6	k->5	m->5	n->21	p->1	r->4	s->34	t->761	x->1	
lv	 ->44	,->5	.->4	a->152	b->5	e->127	f->3	h->2	i->43	k->21	m->1	n->3	o->2	p->1	r->6	s->16	t->10	v->2	ä->36	å->5	ö->3	
ly	 ->2	!->1	,->2	.->2	b->1	c->125	d->8	f->13	g->18	k->17	m->6	r->1	s->107	t->30	v->1	w->1	
lz	 ->3	e->1	m->2	
lä	c->8	d->43	g->376	k->11	m->314	n->327	p->21	r->24	s->24	t->61	x->3	
lå	 ->34	d->13	e->1	g->15	n->124	r->47	s->33	t->124	
lé	c->1	
lö	d->4	f->11	j->9	k->1	m->21	n->15	p->25	r->1	s->179	t->7	v->1	
lø	n->2	
m 	"->8	-->19	1->6	2->4	3->6	4->4	5->2	6->1	8->1	A->9	B->12	C->4	D->8	E->101	F->9	G->8	H->7	I->6	J->4	K->6	L->8	M->4	N->1	O->1	P->9	R->3	S->10	T->12	V->1	W->3	a->644	b->231	c->7	d->745	e->425	f->493	g->170	h->389	i->367	j->159	k->323	l->144	m->365	n->172	o->193	p->137	r->245	s->563	t->216	u->170	v->504	y->5	Ö->4	ä->242	å->54	ö->41	
m!	D->2	M->1	T->1	
m"	.->1	
m)	 ->1	;->1	
m,	 ->164	
m-	 ->1	e->1	
m.	 ->12	(->1	,->1	.->2	A->5	B->2	D->43	E->5	F->8	G->3	H->12	I->6	J->17	K->3	L->1	M->14	N->8	O->7	P->2	R->3	S->9	T->3	U->1	V->21	m->1	Ä->2	
m/	r->1	
m:	 ->7	
m;	 ->2	
m?	D->1	J->1	M->1	V->2	
mI	.->1	
ma	 ->476	,->10	.->10	:->2	c->1	d->11	f->1	g->10	i->8	j->49	k->54	l->30	n->1575	p->1	r->515	s->50	t->185	v->3	x->8	
mb	 ->1	.->1	a->56	e->65	i->27	l->6	n->1	o->10	r->3	u->22	y->1	ä->4	
md	 ->7	,->2	a->9	e->9	h->1	i->1	r->6	ö->2	
me	 ->17	,->1	-->1	.->1	d->2510	g->1	k->11	l->437	n->1992	r->1248	s->50	t->249	u->4	x->2	
mf	a->84	i->1	l->1	o->4	u->5	ä->1	å->2	ö->362	
mg	e->1	i->4	r->4	ä->1	å->66	
mh	e->100	u->1	ä->54	å->17	ö->16	
mi	 ->20	,->3	.->3	?->1	b->2	d->17	e->8	f->1	g->248	i->1	k->15	l->306	n->713	p->1	r->6	s->1503	t->192	u->3	x->2	ä->10	å->1	
mj	a->62	u->3	
mk	a->6	o->10	r->15	
ml	a->65	e->2	i->185	o->2	ä->13	ö->5	
mm	 ->1	a->859	e->1168	i->1265	o->11	u->34	ö->1	
mn	 ->12	,->3	.->4	a->195	b->1	d->26	e->38	i->85	k->2	s->9	t->19	u->4	v->2	
mo	,->2	b->7	c->1	d->84	f->1	g->7	k->142	l->1	m->9	n->68	r->116	s->3	t->515	u->1	
mp	 ->14	.->1	a->157	e->157	i->2	l->123	n->85	o->17	r->56	s->1	t->1	u->7	å->1	
mr	a->24	e->7	i->1	u->3	ä->1	å->325	ö->57	
ms	 ->11	-->4	a->8	b->3	e->5	f->4	g->1	h->2	i->3	k->15	l->42	n->11	o->10	p->3	r->4	s->284	t->326	v->2	y->6	ä->8	å->1	
mt	 ->156	,->6	.->4	a->30	e->16	i->179	l->25	n->1	o->5	r->2	s->4	v->2	y->6	ä->1	å->1	
mu	g->1	l->44	m->4	n->63	r->1	s->9	t->5	
mv	a->5	e->6	i->6	ä->13	
my	c->452	g->1	l->1	n->164	t->1	
má	n->1	
mä	d->1	k->3	l->21	n->367	r->132	s->33	t->9	
må	 ->59	,->2	.->1	e->2	f->6	g->32	h->5	l->205	n->269	r->5	s->697	t->28	
mé	 ->3	a->1	k->1	n->2	s->1	
mö	b->2	d->5	g->2	j->307	n->2	r->9	s->1	t->143	v->2	
n 	"->16	(->45	,->1	-->72	1->96	2->29	3->15	4->5	5->6	6->1	7->3	8->3	9->4	A->19	B->15	C->10	D->11	E->71	F->13	G->10	H->29	I->24	J->6	K->20	L->7	M->2	N->7	O->1	P->20	R->7	S->17	T->11	U->4	V->8	W->24	X->1	a->1400	b->530	c->26	d->756	e->680	f->1282	g->526	h->683	i->1141	j->171	k->727	l->221	m->839	n->328	o->1302	p->541	r->399	s->1549	t->685	u->374	v->648	w->2	y->8	z->2	Ö->3	ä->408	å->109	ö->150	
n!	 ->228	A->1	D->3	E->2	H->1	J->6	M->1	N->2	R->1	S->1	T->2	U->1	V->2	
n"	 ->8	,->5	.->5	
n)	 ->6	(->2	,->1	.->3	J->1	N->1	
n,	 ->1122	
n-	 ->4	C->1	H->1	K->1	S->1	g->1	r->3	
n.	 ->27	"->1	(->5	)->13	.->14	1->2	A->27	B->6	C->2	D->287	E->42	F->61	G->4	H->81	I->45	J->138	K->33	L->14	M->64	N->25	O->35	P->18	R->9	S->58	T->24	U->15	V->121	W->1	Ä->9	Å->3	Ö->3	
n/	N->2	å->2	
n:	 ->35	F->1	
n;	 ->23	
n?	 ->3	.->1	A->1	D->8	E->1	F->5	H->4	I->1	J->4	K->5	N->1	O->1	P->1	S->1	V->11	Ä->5	
nF	r->3	
nH	e->2	
nI	 ->1	
nJ	a->2	
nN	ä->7	
na	 ->3086	!->3	"->3	,->258	-->1	.->307	/->2	:->3	;->5	?->14	H->1	b->73	c->10	d->552	f->2	g->10	i->2	k->4	l->258	m->27	n->245	p->20	r->436	s->436	t->590	u->1	v->6	z->16	
nb	a->69	e->24	i->9	j->7	l->32	o->3	r->2	u->9	y->1	
nc	 ->1	,->1	a->2	e->46	h->3	i->208	k->14	
nd	 ->501	!->2	)->1	,->49	-->1	.->47	?->4	a->615	b->11	e->4107	f->9	g->5	i->462	k->1	l->456	m->4	n->78	o->25	p->105	r->883	s->174	t->8	u->118	v->67	z->4	ä->1	å->58	é->1	ö->1	
ne	 ->72	!->1	,->9	-->5	.->4	:->1	a->2	b->117	d->66	e->1	f->14	g->26	h->85	j->5	k->13	l->290	m->4	n->1671	o->2	p->5	r->1209	s->43	t->53	u->2	v->2	z->2	
nf	a->14	e->174	i->7	l->29	o->92	r->22	ä->1	ö->226	
ng	 ->1506	!->1	"->6	)->6	,->215	-->1	.->271	:->4	;->4	?->7	a->952	b->1	d->53	e->1269	f->42	g->2	i->16	k->1	l->39	m->7	n->52	o->4	p->2	r->102	s->1073	t->78	u->2	v->6	ä->1	å->85	ö->3	
nh	a->50	e->246	i->1	o->6	u->1	ä->43	å->56	ö->4	
ni	 ->240	,->16	.->3	a->1	c->2	e->70	f->3	g->21	k->33	l->2	m->28	n->2453	o->465	p->5	r->1	s->385	t->156	u->5	v->114	é->1	
nj	 ->3	.->1	e->95	o->1	u->4	ä->2	ö->2	
nk	 ->8	"->1	-->1	.->1	a->364	b->4	e->180	f->9	i->3	l->51	n->20	o->28	r->132	s->7	t->409	u->285	ä->1	ö->3	
nl	a->11	e->124	i->247	y->1	ä->45	å->2	ö->6	
nm	a->27	ä->34	ö->2	
nn	 ->5	,->2	-->1	a->1279	d->1	e->540	h->1	i->229	l->7	o->105	s->353	u->80	y->2	ä->3	
no	 ->8	,->2	.->2	c->24	d->3	g->43	i->1	k->3	l->15	m->1062	n->13	p->19	r->201	s->7	t->31	v->20	w->1	
np	a->14	o->2	r->4	u->31	å->1	
nr	 ->29	a->14	e->91	i->57	y->2	ä->56	å->1	ö->7	
ns	 ->1493	!->1	,->43	-->6	.->26	/->1	:->1	;->1	?->3	a->359	b->15	c->9	d->14	e->644	f->33	g->1	h->13	i->165	j->17	k->903	l->129	m->25	n->23	o->8	p->226	r->59	s->44	t->720	u->77	v->335	y->85	ä->16	å->14	ö->23	
nt	 ->460	!->1	,->41	-->1	.->47	:->2	a->499	e->2606	f->6	i->246	k->2	l->249	n->8	o->42	p->3	r->550	s->66	t->1	u->26	v->4	y->19	ä->7	ó->1	ö->3	
nu	 ->281	,->6	.->8	:->1	;->1	?->1	a->16	c->1	e->2	f->14	l->2	m->12	n->1	p->4	s->7	t->27	v->45	
nv	a->39	e->56	i->59	o->9	ä->223	å->9	
ny	 ->39	a->173	b->41	c->8	d->1	e->8	f->2	h->13	k->3	l->30	m->5	n->6	o->4	p->1	s->14	t->131	v->1	å->1	
nz	 ->17	)->2	,->3	F->1	b->1	e->1	á->1	
nÄ	r->1	
nä	c->2	e->1	g->1	l->2	m->137	r->736	s->48	t->23	v->1	
nå	 ->67	,->1	.->4	b->2	d->8	g->505	l->5	r->17	s->7	t->20	
nç	o->1	
nè	v->3	
nö	d->140	j->29	r->4	s->19	t->6	v->3	
o 	(->2	-->3	1->1	C->5	E->1	L->1	P->2	R->1	S->1	T->3	V->4	a->10	b->5	d->3	e->1	f->24	g->6	h->5	i->12	k->5	l->2	m->13	n->5	o->21	p->8	r->1	s->22	t->7	u->4	v->5	ä->10	å->9	ö->2	
o!	A->1	
o,	 ->45	
o-	 ->1	P->4	a->2	p->1	r->1	
o.	 ->1	-->1	A->2	B->1	D->6	E->1	F->4	H->3	J->5	K->2	L->1	M->1	N->2	O->4	S->1	T->2	V->5	m->7	
o/	O->1	
o:	 ->1	
o;	 ->1	
o?	 ->1	H->1	
oN	ä->1	
oU	,->1	-->1	
oa	 ->3	c->31	d->5	k->15	l->14	n->17	r->7	t->1	v->12	
ob	 ->2	a->21	b->16	e->75	i->8	j->1	l->198	o->3	s->2	
oc	-->2	a->1	e->204	h->4577	i->212	k->699	o->1	
od	 ->91	,->5	.->3	?->1	a->50	d->10	e->137	f->1	i->53	j->2	k->89	l->17	o->5	s->39	t->46	u->85	w->1	
oe	b->1	d->14	f->4	g->5	k->10	l->2	n->138	r->13	t->8	
of	 ->25	,->4	.->4	a->3	d->1	e->63	f->114	h->1	i->12	o->1	r->4	s->4	t->55	u->2	ö->25	
og	 ->98	,->3	.->11	a->75	b->1	e->54	g->12	i->49	j->1	k->1	m->2	r->257	s->49	u->1	y->1	å->1	ö->9	
oh	a->3	e->1	j->2	o->1	ä->1	ö->1	
oi	g->1	j->1	n->6	r->4	s->6	
oj	a->7	e->64	k->2	o->1	u->6	ä->7	
ok	 ->24	,->5	.->5	a->52	e->39	i->2	l->16	o->35	r->143	s->2	t->13	u->57	ä->2	
ol	 ->26	,->7	-->2	.->6	;->1	a->67	b->2	d->7	e->76	f->12	i->752	j->42	k->161	l->498	m->3	n->1	o->36	p->1	s->18	t->11	u->145	v->11	y->53	z->2	ä->5	ö->2	
om	 ->6192	!->1	"->1	)->2	,->58	-->1	.->36	/->1	I->1	a->54	b->37	d->10	e->62	f->252	g->22	h->1	i->317	k->15	l->23	m->2289	n->45	o->14	p->101	r->361	s->215	t->2	u->1	v->17	á->1	ä->1	å->3	é->5	ö->16	
on	 ->629	"->1	)->2	,->72	-->2	.->103	/->2	:->3	;->1	?->9	N->1	a->215	b->16	c->56	d->149	e->2424	f->193	g->5	h->1	i->46	j->3	k->343	l->35	m->5	n->2	o->338	r->1	s->436	t->312	v->33	y->5	z->1	ä->248	å->1	ö->11	
oo	 ->1	d->4	i->1	l->1	m->1	p->1	s->1	
op	 ->12	,->6	-->1	.->4	a->480	e->727	i->10	l->1	o->47	p->182	r->8	t->8	u->7	y->1	å->1	é->10	
or	 ->688	)->1	,->83	.->83	:->4	;->1	?->4	a->215	b->18	c->5	d->832	e->162	f->2	g->319	h->2	i->238	k->7	l->7	m->463	n->152	o->87	p->8	r->51	s->177	t->844	u->6	v->6	w->1	ä->13	ê->1	ö->4	
os	 ->94	!->1	,->3	a->7	e->3	f->1	i->89	j->1	k->9	l->2	m->4	n->2	o->66	p->2	s->334	t->167	v->6	y->5	ä->17	å->1	
ot	 ->539	!->8	,->20	.->11	?->1	a->83	b->2	e->100	f->3	g->1	h->11	i->53	j->1	n->17	o->42	p->6	r->3	s->140	t->296	u->4	v->9	y->4	ä->1	å->4	
ou	 ->2	c->12	k->1	l->6	m->4	n->7	p->2	r->24	s->2	t->4	x->1	
ov	 ->51	"->1	,->3	.->5	a->32	e->67	i->32	j->1	k->2	o->63	s->9	v->2	y->1	ä->23	å->3	
ow	 ->1	-->1	e->5	i->3	n->3	
ox	 ->2	!->1	,->2	a->5	i->8	n->1	
oy	a->1	d->1	o->2	
oä	m->1	n->16	
oå	r->1	
oö	n->1	v->6	
p 	(->2	,->1	-->3	C->1	E->1	J->1	T->1	a->100	b->7	d->48	e->25	f->39	g->4	h->13	i->47	k->8	l->5	m->18	n->7	o->34	p->18	r->7	s->39	t->23	u->12	v->10	ä->15	ö->2	
p"	 ->1	!->1	,->2	
p,	 ->53	
p-	s->1	
p.	 ->3	.->1	A->1	D->16	E->2	F->1	H->1	I->4	J->12	M->1	P->1	S->3	T->1	V->8	g->1	Ä->2	
p:	 ->1	
p?	H->1	
pa	 ->411	!->2	"->1	,->39	.->62	;->1	?->3	N->1	c->10	d->27	g->6	k->13	l->12	m->1	n->96	p->171	r->842	s->261	t->41	v->3	y->2	
pb	a->1	r->3	y->20	ä->1	å->1	
pd	a->3	e->3	r->22	
pe	 ->2	a->2	c->85	d->3	g->13	h->13	i->712	k->222	l->177	n->565	r->497	s->10	t->158	
pf	a->53	y->54	ö->24	
pg	i->80	o->1	r->1	å->15	ö->2	
ph	a->1	e->7	o->13	t->1	ä->6	å->3	ö->10	
pi	a->1	c->2	e->12	l->5	n->5	o->1	r->4	s->2	t->37	
pj	a->1	
pk	a->11	o->7	r->1	
pl	a->206	e->61	i->177	o->13	u->4	y->4	ä->2	å->15	ö->8	
pm	a->58	j->2	u->21	ä->55	ö->12	
pn	a->19	e->2	i->119	å->93	
po	,->1	e->1	k->4	l->590	n->19	o->1	p->7	r->324	s->103	t->14	u->5	ä->12	
pp	 ->285	,->24	.->22	?->1	a->140	b->26	d->28	e->298	f->130	g->91	h->33	j->1	k->7	l->45	m->148	n->126	o->120	r->111	s->94	t->42	u->1	v->10	y->1	
pr	a->49	e->202	i->322	o->860	u->20	y->1	ä->45	å->26	ö->20	
ps	 ->6	-->1	.->2	a->9	b->6	d->1	f->1	i->16	k->35	l->5	m->20	n->11	o->2	p->9	r->21	s->7	t->39	v->2	y->1	ä->3	å->2	
pt	 ->23	.->2	a->57	e->75	i->30	o->5	r->10	ä->11	
pu	b->26	l->13	m->2	n->346	r->1	s->5	
pv	e->2	i->7	ä->2	
py	 ->1	r->2	
pä	n->11	r->3	
på	 ->1768	,->16	.->16	:->3	?->2	b->12	d->1	f->5	g->21	l->4	m->30	p->50	r->13	s->28	t->16	v->40	
pé	 ->1	e->9	r->1	
pö	k->4	
qa	l->2	
qu	a->10	e->7	i->5	o->2	q->2	
r 	"->8	(->7	-->87	1->90	2->73	3->16	4->11	5->6	6->2	7->6	8->6	9->5	A->14	B->34	C->9	D->6	E->151	F->18	G->12	H->5	I->16	J->6	K->22	L->17	M->22	N->6	O->5	P->37	R->9	S->22	T->18	U->5	V->6	W->6	[->1	a->2806	b->563	c->26	d->2496	e->1327	f->1370	g->368	h->552	i->1322	j->369	k->735	l->355	m->1135	n->477	o->1328	p->591	r->394	s->1831	t->1029	u->510	v->1055	y->20	Ö->8	ä->315	å->105	ö->172	
r!	 ->119	"->2	.->1	D->7	E->2	J->5	M->3	T->1	V->2	
r"	 ->6	)->1	,->1	.->3	
r)	 ->5	.->1	?->1	F->2	J->1	K->1	T->1	
r,	 ->980	
r-	 ->5	b->1	k->1	n->1	p->11	r->1	
r.	 ->29	(->3	)->2	-->4	.->11	9->1	A->14	B->13	C->1	D->245	E->36	F->60	G->8	H->37	I->40	J->119	K->34	L->11	M->41	N->19	O->28	P->10	R->11	S->27	T->25	U->8	V->109	k->1	Ä->13	Å->2	Ö->1	
r:	 ->45	
r;	 ->14	
r?	,->1	-->1	.->1	B->1	D->3	E->1	F->2	H->6	I->2	J->3	K->3	M->2	N->3	P->1	S->1	T->1	V->3	Ä->3	
rH	e->1	
rJ	a->1	
rM	e->1	
rN	ä->2	
ra	 ->3175	!->2	"->2	,->73	.->74	:->7	;->2	?->3	b->66	c->5	d->441	e->58	f->217	g->432	h->2	i->2	k->126	l->172	m->1021	n->1312	o->1	p->111	r->581	s->487	t->635	u->1	v->111	x->11	y->1	ç->5	
rb	,->1	a->28	e->625	i->40	j->34	l->18	r->24	u->38	ä->78	ö->12	
rc	e->4	o->1	y->4	
rd	 ->102	)->1	,->18	-->2	.->14	:->2	;->3	a->170	b->67	e->615	f->223	h->1	i->58	j->11	k->1	l->9	m->1	n->186	o->79	r->203	s->25	t->2	u->3	v->3	ä->4	ö->21	
re	 ->1120	!->1	"->3	,->88	-->1	.->86	:->2	?->4	a->70	b->30	c->54	d->618	e->7	f->183	g->752	h->2	i->1	j->7	k->385	l->157	m->78	n->1105	p->128	r->262	s->795	t->532	u->6	v->54	x->6	y->6	z->1	
rf	a->116	e->7	i->7	j->1	l->21	o->109	r->14	u->2	ä->4	å->1	ö->368	
rg	 ->34	,->6	.->4	a->273	e->40	h->1	i->132	l->5	m->2	n->1	o->39	r->22	s->1	u->17	ä->2	å->20	ö->17	
rh	a->102	e->311	i->32	o->16	u->10	ä->5	å->72	ö->18	
ri	 ->75	!->1	,->21	-->10	.->6	a->72	b->11	c->15	d->114	e->139	f->44	g->310	h->118	k->587	l->9	m->61	n->1524	o->131	p->69	r->1	s->371	t->372	u->13	v->155	ä->4	è->1	ö->8	
rj	a->126	d->1	e->93	n->4	
rk	 ->67	,->7	-->1	.->8	?->1	a->321	b->4	d->1	e->124	i->48	k->2	l->297	m->2	n->229	o->26	r->3	s->132	t->72	u->6	ä->42	ö->1	
rl	 ->5	-->1	a->645	d->59	e->16	i->508	o->20	s->2	u->13	y->2	ä->89	å->15	ö->2	ø->2	
rm	 ->62	,->9	-->1	.->7	:->1	a->210	e->229	f->3	i->26	n->31	o->36	p->15	r->2	s->4	t->19	u->18	y->15	ä->1	å->50	é->3	ö->3	
rn	 ->82	)->1	,->24	-->2	.->22	/->2	?->1	a->2252	b->1	d->3	e->36	f->3	h->1	i->68	k->23	o->2	p->6	s->23	t->9	u->14	v->23	y->49	ä->1	ö->2	
ro	 ->72	!->1	,->15	-->1	.->18	a->36	b->183	c->205	d->132	e->146	f->103	g->255	i->1	j->71	k->14	l->269	m->45	n->45	o->1	p->1234	r->288	s->21	t->200	u->3	v->60	
rp	a->17	e->4	l->22	n->1	o->24	r->6	t->4	u->5	å->2	
rq	u->1	
rr	 ->536	,->4	.->1	?->1	a->118	e->424	g->4	i->167	o->14	u->9	v->1	ä->7	å->15	ó->3	ö->5	
rs	 ->258	,->20	-->1	.->24	a->69	b->7	c->1	d->8	e->110	f->56	h->1	i->110	k->284	l->497	m->5	o->312	p->50	r->2	s->3	t->636	u->12	v->90	y->3	ä->111	å->2	ö->114	
rt	 ->771	!->2	)->1	,->49	-->3	.->46	:->2	?->1	N->1	a->77	b->3	d->1	e->235	f->100	g->9	h->3	i->305	j->21	k->19	l->9	m->2	n->31	o->35	p->3	r->79	s->186	u->104	v->2	y->111	z->3	ä->3	
ru	 ->149	,->1	a->16	b->5	c->2	e->5	h->2	i->1	k->283	l->6	m->107	n->341	p->238	s->20	t->112	v->16	
rv	 ->3	,->3	.->3	a->170	b->1	e->47	h->1	i->113	j->3	l->2	r->2	s->6	t->3	u->3	ä->103	å->6	
rw	e->1	
ry	 ->2	,->1	.->1	c->105	f->1	g->19	k->43	m->16	o->1	p->6	r->2	s->27	t->21	
rz	w->1	
rä	 ->2	c->153	d->193	f->147	g->43	k->66	l->3	m->153	n->348	p->2	r->2	s->3	t->756	v->175	
rå	 ->3	d->776	e->2	g->859	k->59	l->8	n->628	o->1	p->1	r->12	s->2	t->3	z->1	
ré	b->1	f->1	
rê	t->1	
rí	n->1	
ró	n->5	
rö	d->13	g->1	j->16	k->3	m->22	n->21	r->151	s->192	t->15	v->24	
s 	"->2	(->3	-->21	1->5	2->5	3->1	4->1	8->1	A->2	B->7	C->1	D->4	E->17	F->1	G->3	H->1	I->1	L->1	M->1	O->1	P->1	R->2	S->6	V->2	W->2	X->1	a->666	b->223	c->9	d->309	e->289	f->534	g->128	h->140	i->539	j->34	k->170	l->105	m->343	n->128	o->429	p->282	q->2	r->200	s->515	t->246	u->240	v->197	y->21	ä->85	å->62	ö->59	
s!	 ->2	D->1	E->1	F->1	G->1	H->1	V->1	
s"	.->3	
s)	 ->2	
s,	 ->303	
s-	 ->43	,->1	C->1	J->2	b->3	d->1	f->1	i->2	n->2	p->1	s->1	
s.	 ->52	(->1	)->1	-->1	.->1	A->6	B->6	C->1	D->101	E->20	F->18	G->5	H->18	I->15	J->31	K->8	L->4	M->21	N->8	O->5	P->8	R->6	S->13	T->5	U->6	V->40	Y->2	k->4	Ä->5	Å->2	
s/	d->1	i->1	
s:	 ->7	
s;	 ->6	
s?	.->2	D->1	E->1	F->1	H->1	I->1	J->2	K->1	O->1	S->1	T->1	V->2	Ä->1	
sN	ä->1	
sa	 ->701	!->1	,->22	.->28	?->1	b->12	c->4	d->132	f->4	g->51	i->1	k->193	l->7	m->1167	n->116	r->131	s->36	t->304	u->1	v->26	
sb	a->9	e->78	i->11	o->11	r->20	u->6	y->44	å->1	ö->12	
sc	a->6	e->16	h->37	i->27	o->1	y->3	
sd	a->15	e->18	i->15	o->10	r->5	u->6	ö->2	
se	 ->362	"->1	,->19	-->2	.->28	;->1	?->1	a->1	b->2	d->111	e->60	f->18	g->22	h->1	i->3	k->203	l->143	m->12	n->691	o->1	p->16	r->1089	s->34	t->110	u->2	v->16	w->1	x->26	
sf	a->26	e->2	i->35	l->18	o->31	r->109	u->18	ä->2	å->1	ö->292	
sg	a->7	e->1	i->17	r->21	y->7	å->3	ö->1	
sh	 ->2	,->1	a->19	e->53	i->15	j->2	o->2	u->2	ä->3	å->1	
si	a->5	b->1	d->133	e->94	f->37	g->442	k->224	l->7	m->5	n->390	o->1299	s->195	t->328	v->45	ä->2	
sj	o->17	u->36	ä->192	ö->21	
sk	 ->363	,->7	-->4	.->13	a->3278	b->8	e->275	f->4	h->7	i->314	j->31	k->3	l->70	n->78	o->542	r->279	t->277	u->667	v->24	y->162	ä->78	å->12	ö->33	
sl	a->680	e->47	i->231	o->35	u->532	y->18	ä->74	å->110	ö->67	
sm	 ->38	,->11	.->20	?->1	a->40	e->155	i->29	o->10	u->6	y->31	ä->51	å->79	ö->7	
sn	a->173	e->13	i->158	o->7	y->2	ä->5	å->6	ö->4	
so	 ->6	,->1	-->1	c->208	d->1	e->1	f->8	l->186	m->3714	n->130	p->1	r->89	s->6	t->1	v->64	
sp	"->1	.->2	a->43	e->339	i->7	l->54	o->252	r->254	u->18	ä->14	å->14	ö->4	
sq	u->2	
sr	a->73	e->66	i->21	o->1	u->7	y->3	ä->62	å->23	ö->2	
ss	 ->486	"->1	)->1	,->24	.->34	:->1	?->3	a->607	b->15	c->1	e->360	f->7	g->7	h->6	i->1297	j->1	k->44	l->34	m->4	n->38	o->17	p->3	r->5	t->445	u->65	v->5	y->59	ä->84	
st	 ->654	!->2	,->26	-->6	.->23	:->1	?->2	a->1696	b->9	d->11	e->1782	f->18	g->6	h->6	i->538	j->9	k->5	l->9	m->7	n->183	o->553	p->5	r->903	s->81	t->3	u->39	v->7	y->61	ä->853	å->605	ê->1	ö->584	
su	a->1	b->38	c->5	d->1	e->2	g->1	l->127	m->85	n->12	p->7	r->53	s->5	t->96	v->17	
sv	.->6	a->515	e->15	i->78	u->4	ä->49	å->98	
sw	a->1	
sy	d->5	f->74	k->1	l->21	m->18	n->224	r->11	s->301	
sä	g->269	k->400	l->20	m->22	n->30	r->166	s->1	t->683	
så	 ->1115	,->18	.->9	:->1	d->163	g->23	h->1	l->46	n->3	r->4	s->32	t->15	v->43	
sí	 ->1	
sö	d->8	k->143	n->8	r->16	v->16	
t 	"->15	(->24	,->1	-->92	1->28	2->10	3->3	4->6	5->4	6->1	7->4	8->4	9->6	:->1	A->13	B->10	C->4	D->10	E->161	F->18	G->7	H->5	I->13	J->6	K->11	L->3	M->9	N->1	O->3	P->8	R->8	S->13	T->22	U->1	V->4	W->3	a->2059	b->872	c->18	d->1612	e->805	f->2245	g->841	h->766	i->1202	j->152	k->916	l->413	m->1334	n->438	o->1266	p->785	r->437	s->2495	t->802	u->667	v->1290	w->1	y->35	z->1	Ö->6	ä->1054	å->143	ö->189	
t!	 ->7	"->1	(->1	.->2	D->2	H->3	J->1	K->1	L->1	M->1	N->1	P->1	T->1	
t"	 ->5	,->4	.->2	
t)	 ->7	,->3	.->4	N->1	
t,	 ->1019	
t-	 ->3	E->1	a->5	b->5	f->1	s->2	
t.	 ->38	(->5	)->5	-->1	.->6	1->1	A->21	B->11	D->268	E->44	F->68	G->7	H->67	I->50	J->149	K->23	L->15	M->86	N->33	O->34	P->23	R->6	S->38	T->20	U->9	V->117	e->20	o->7	Ä->11	Å->6	Ö->3	
t:	 ->35	
t;	 ->13	
t?	 ->2	.->4	A->3	D->4	E->2	H->3	I->1	J->5	K->2	N->6	O->2	R->1	S->2	T->1	U->1	V->5	Ä->1	
tB	e->1	
tJ	a->1	
tN	ä->1	
ta	 ->2625	!->2	,->82	.->116	:->6	;->2	?->4	N->1	a->1	b->95	c->149	d->198	f->10	g->556	i->26	k->39	l->1189	m->12	n->842	p->9	r->615	s->309	t->903	u->5	v->10	x->4	
tb	a->11	e->15	i->65	l->1	o->54	r->6	u->5	y->20	
tc	.->5	?->1	h->2	
td	e->15	i->2	
te	 ->2690	!->2	,->38	-->2	.->51	:->2	?->5	a->4	b->16	c->47	d->7	e->9	f->10	g->181	i->3	k->59	l->80	m->290	n->1376	o->2	p->2	r->3536	s->81	t->1244	u->9	x->45	
tf	a->102	e->1	l->4	o->42	r->17	u->15	ä->30	å->1	ö->126	
tg	a->1	i->27	j->4	r->7	ä->245	å->47	ö->63	
th	 ->4	,->1	-->7	a->6	e->16	i->2	o->3	u->8	y->1	ä->5	å->11	ö->1	
ti	 ->61	!->3	"->1	,->14	-->3	.->16	a->84	b->11	c->11	d->608	e->96	f->188	g->759	h->1	i->1	k->479	l->2692	m->54	n->181	o->1282	p->3	q->2	r->1	s->640	t->222	v->707	ö->12	
tj	a->42	o->2	u->5	ä->184	
tk	a->17	l->1	o->41	r->5	u->3	v->1	ä->1	ö->3	
tl	a->22	e->12	i->608	o->3	ä->22	å->2	ö->5	
tm	a->26	e->3	i->28	o->1	y->4	ä->36	å->1	
tn	a->164	e->40	i->662	j->1	y->42	ä->9	
to	 ->16	-->2	.->2	/->1	a->2	b->12	c->3	d->45	g->68	k->26	l->154	m->140	n->132	p->35	r->642	s->14	t->34	w->3	x->1	
tp	a->9	e->12	l->6	o->13	r->8	u->3	
tr	a->606	e->446	i->216	o->620	u->272	y->155	ä->430	å->15	ö->30	
ts	 ->859	!->1	,->48	-->13	.->54	:->1	?->2	a->154	b->22	c->6	d->5	e->143	f->53	g->19	h->4	i->15	k->204	l->265	m->35	n->17	o->30	p->114	r->35	s->92	t->211	u->8	v->30	y->2	ä->170	å->68	
tt	 ->8485	,->85	.->119	:->6	?->5	B->1	a->1755	e->694	f->10	g->1	h->9	i->245	j->66	k->2	l->11	m->2	n->313	o->17	r->282	s->287	v->75	y->2	ä->1	é->59	ö->5	
tu	 ->21	a->130	d->15	e->58	f->2	g->98	l->43	m->88	n->43	r->495	s->27	t->172	
tv	a->6	e->304	i->406	u->11	ä->57	å->132	
ty	 ->13	-->1	c->94	d->257	g->120	m->3	n->11	p->42	r->64	s->28	v->30	
tz	 ->3	,->1	.->1	i->2	
tä	c->31	d->21	k->5	l->426	m->230	n->503	p->4	r->76	t->5	v->5	
tå	 ->65	,->3	.->2	:->1	d->2	e->46	g->5	l->47	n->226	r->193	s->6	t->34	
té	 ->10	e->4	f->2	n->41	s->2	
tê	t->3	
tó	n->1	
tö	d->434	k->12	l->1	m->6	r->171	t->19	v->37	
tü	r->1	
u 	-->1	3->1	A->3	B->1	E->2	F->1	L->1	M->2	P->2	R->3	S->4	T->1	W->1	a->21	b->13	c->1	d->13	e->25	f->31	g->15	h->29	i->56	k->59	l->8	m->50	n->10	o->18	p->11	r->7	s->41	t->96	u->5	v->12	ä->33	å->2	
u"	,->1	
u,	 ->18	
u-	l->1	
u.	.->1	D->1	E->1	J->1	K->2	L->1	V->2	
u:	 ->1	
u;	 ->1	
u?	J->1	
uM	e->1	
ua	 ->2	d->1	l->11	n->1	r->32	t->130	
ub	b->20	e->1	i->2	j->1	l->34	r->2	s->27	v->12	
uc	 ->1	c->5	e->35	h->12	k->7	t->1	
ud	 ->34	,->4	.->3	a->31	d->8	e->38	f->5	g->107	i->15	l->3	m->2	n->3	o->1	r->6	s->50	u->1	
ue	 ->1	,->2	c->1	i->1	l->68	n->1	r->15	s->6	
uf	f->2	m->1	t->16	ö->1	
ug	a->28	e->3	g->8	i->70	l->6	n->6	o->6	u->1	
uh	a->1	e->2	n->1	
ui	e->1	g->1	n->2	o->1	s->4	t->1	z->1	
uk	 ->10	!->1	,->9	.->1	a->26	d->1	e->20	f->1	h->7	i->1	n->3	s->23	t->266	v->3	
ul	 ->4	.->1	a->25	d->6	e->65	f->4	g->1	i->15	k->1	l->666	o->6	s->7	t->307	z->3	ä->4	
um	 ->139	!->2	,->12	.->18	a->8	b->5	e->188	g->1	h->3	l->1	m->26	p->12	r->1	t->4	u->2	ä->1	ö->2	
un	 ->1	.->1	a->6	c->3	d->1040	e->11	g->151	h->1	i->479	k->391	n->290	o->1	s->17	t->44	
uo	 ->1	,->1	
up	 ->3	a->15	e->8	g->7	n->5	p->1258	r->1	s->2	t->14	é->1	
uq	a->2	
ur	 ->343	,->21	-->4	.->14	?->1	a->38	b->2	d->1	e->141	f->65	g->16	h->5	i->76	k->59	l->110	m->2	n->6	o->1267	p->20	r->287	s->114	t->5	u->18	v->15	å->1	
us	 ->31	,->5	-->1	.->6	?->1	a->5	c->1	d->1	e->38	f->1	g->6	h->3	i->35	k->2	l->1	p->2	q->1	s->72	t->292	u->6	í->1	ö->1	
ut	 ->240	,->34	.->34	:->1	;->1	?->2	a->543	b->97	d->1	e->215	f->112	g->118	h->6	i->298	j->5	k->23	l->91	m->53	n->103	o->103	p->7	r->58	s->401	t->213	v->384	y->1	ä->5	å->1	ö->42	
uu	m->2	
uv	a->47	e->21	i->15	r->1	u->54	
ux	,->2	-->1	e->6	h->1	i->1	n->2	
uy	u->2	
v 	"->3	(->1	-->9	1->4	2->1	4->2	5->2	8->1	9->8	A->5	B->20	C->1	D->7	E->92	F->12	G->6	H->3	I->2	J->4	K->14	L->5	M->4	O->5	P->4	R->2	S->7	T->8	U->1	V->3	W->3	a->213	b->92	c->9	d->613	e->219	f->254	g->53	h->47	i->63	j->11	k->162	l->62	m->114	n->39	o->118	p->114	r->75	s->272	t->106	u->73	v->107	y->5	Ö->2	ä->17	å->26	ö->16	
v"	,->1	
v,	 ->49	
v.	 ->5	"->1	(->1	,->1	.->3	?->1	A->3	B->2	D->13	E->4	F->5	H->1	I->3	J->2	K->1	L->1	M->3	O->2	R->2	S->2	U->1	V->3	Y->1	
v:	 ->2	
v;	 ->1	
v?	F->1	N->1	V->1	
va	 ->305	,->9	.->8	?->1	c->9	d->251	g->49	k->53	l->243	n->165	p->28	r->1693	s->32	t->109	v->7	
vb	e->4	i->1	o->1	r->16	ä->1	
vd	a->27	e->16	v->1	
ve	 ->37	,->2	-->3	N->1	b->1	c->290	d->13	k->37	l->49	m->29	n->524	p->4	r->1540	s->20	t->497	u->1	
vf	a->25	o->1	ö->8	
vg	a->2	e->10	i->9	j->4	r->4	å->7	ö->61	
vh	e->1	j->4	ä->2	å->1	
vi	 ->1635	,->16	.->1	?->1	a->13	c->24	d->495	e->3	f->1	g->7	k->420	l->1213	n->228	r->16	s->817	t->146	v->43	
vj	a->1	e->1	u->3	
vk	a->1	l->21	o->2	r->4	u->1	
vl	a->22	e->2	i->14	o->1	ä->10	å->1	
vm	a->1	i->1	
vn	a->25	i->36	
vo	 ->26	,->11	.->12	?->2	N->1	f->1	k->7	l->18	n->18	r->34	s->7	t->20	å->1	
vp	l->1	r->1	
vr	a->15	e->3	i->82	u->1	ä->8	
vs	 ->100	,->10	.->57	?->1	a->11	c->3	d->2	e->95	f->2	i->41	k->38	l->89	m->98	n->4	o->1	p->5	s->2	t->49	u->1	v->2	ä->6	
vt	 ->130	,->7	.->7	a->90	i->3	r->1	s->3	v->1	
vu	d->54	l->2	n->23	x->3	
vv	a->6	e->10	i->23	ä->7	
vy	t->1	
vä	c->23	d->12	g->203	k->3	l->251	m->23	n->464	p->2	r->341	s->40	t->6	v->7	x->55	
vå	 ->170	,->13	.->22	:->2	;->1	?->1	d->1	e->14	g->14	h->1	l->13	n->38	r->503	
vö	,->1	.->1	n->1	r->1	
w 	Y->1	f->1	t->1	
w,	 ->1	
w-	h->1	
w.	M->1	
wa	g->1	l->2	n->1	r->1	
we	.->2	b->1	i->1	l->1	r->3	
wi	e->1	l->1	s->2	t->2	
wn	 ->2	,->1	
wo	b->3	o->3	r->1	
x 	a->7	e->2	f->1	i->1	m->11	o->1	p->2	s->1	t->2	ö->1	
x!	J->1	
x,	 ->5	
x-	a->1	f->3	
x.	 ->20	D->1	J->1	
xa	 ->3	,->1	.->2	k->18	l->5	m->16	n->9	s->7	t->1	
xb	e->1	
xc	e->6	
xe	l->4	m->124	n->1	r->8	
xf	i->1	
xh	a->1	
xi	b->27	d->5	k->1	l->2	m->9	n->2	s->29	t->1	
xk	l->3	
xl	a->3	i->2	
xm	å->1	
xn	a->2	i->1	
xo	n->3	r->1	
xp	a->6	e->47	l->3	o->6	
xt	 ->20	,->7	.->3	b->1	e->44	h->7	o->1	r->37	s->3	
xu	e->3	p->1	
xv	ä->1	
xx	o->3	
y 	-->1	C->3	E->1	F->1	b->1	d->4	e->3	f->8	g->1	h->3	i->4	k->8	l->3	m->1	n->2	o->4	p->4	r->2	s->7	t->1	u->2	v->8	ä->1	å->1	
y!	 ->1	
y,	 ->9	
y-	p->1	
y.	A->1	D->1	V->2	
yD	e->1	
ya	 ->167	,->1	;->1	b->3	g->4	l->1	n->6	r->2	s->2	v->1	
yb	a->39	e->2	i->3	
yc	k->794	l->1	
yd	 ->4	.->1	a->23	d->113	e->104	i->11	k->2	l->125	o->2	s->1	v->1	ö->1	
ye	 ->2	-->2	d->2	l->6	n->1	r->4	t->1	
yf	a->2	t->94	ö->2	
yg	 ->35	)->1	,->4	.->4	;->1	?->1	a->39	b->1	d->45	e->27	g->118	i->2	k->1	n->1	p->4	r->2	s->17	t->5	
yh	e->13	u->1	ö->1	
yi	s->2	
yk	.->1	a->31	e->10	l->4	o->1	s->2	t->29	
yl	 ->4	,->2	-->1	.->3	a->2	b->1	d->29	f->2	i->35	l->71	r->2	s->6	
ym	 ->4	.->1	a->2	b->9	d->2	e->2	i->1	m->18	p->14	r->10	s->1	t->2	
yn	 ->86	,->2	.->4	;->1	a->16	d->188	e->9	g->12	l->8	n->78	o->1	p->29	s->7	t->4	v->12	
yo	 ->1	l->2	n->3	s->1	t->7	
yp	 ->20	,->2	.->2	e->17	f->1	g->1	h->3	l->1	o->2	p->2	s->1	t->4	
yr	 ->5	.->1	a->53	d->1	e->17	i->33	k->39	n->9	s->2	t->6	å->36	
ys	 ->32	,->4	-->1	.->5	?->2	a->16	e->28	i->9	k->48	n->5	s->181	t->198	
yt	a->28	e->29	i->1	l->2	n->3	s->1	t->275	
yu	 ->2	
yv	a->1	e->2	ä->40	
yw	o->1	
yx	f->1	
yå	r->1	
z 	F->5	G->1	a->1	b->1	d->1	e->3	f->4	h->1	i->1	o->9	s->4	t->2	
z)	(->1	.->1	
z,	 ->9	
z-	k->3	
z.	 ->1	
zF	r->1	
za	 ->1	,->1	.->2	k->1	r->2	
zb	e->3	
ze	n->1	s->1	
zi	d->2	g->4	o->4	s->21	
zj	i->5	
zm	a->2	
zo	n->8	r->2	
zq	u->1	
zu	e->1	
zw	a->1	
zá	l->1	
º 	C->1	
Äm	n->1	
Än	 ->3	d->20	n->3	t->1	
Är	 ->27	a->6	
Äv	e->46	
Å 	E->1	P->1	a->10	e->2	k->1	s->1	
ÅD	S->1	
ÅG	O->1	
År	 ->5	e->1	l->1	
Åt	a->1	e->4	g->5	
Îl	e->1	
Ö 	(->2	f->1	h->1	i->1	m->1	o->4	s->1	v->1	ä->1	
Ö)	 ->1	.->1	
Ö-	l->1	m->1	
Ö:	s->4	
ÖS	T->2	
ÖV	P->6	
Ög	o->2	
Ök	a->1	
Öp	p->1	
Ös	t->88	
Öv	e->2	r->1	
ál	e->1	
án	,->1	c->1	
ão	 ->2	
ä 	u->1	ö->1	
äc	k->220	
äd	 ->5	,->1	.->1	a->80	d->31	e->111	j->24	r->1	s->17	
äe	r->1	
äf	f->117	t->32	
äg	 ->34	,->16	.->9	:->1	N->1	a->275	b->1	d->4	e->199	g->299	l->12	m->1	n->56	r->34	s->24	t->11	
äk	a->6	e->334	n->56	r->64	t->34	
äl	 ->138	,->5	.->9	a->3	b->1	d->32	e->16	f->12	g->3	h->1	i->1	j->30	k->54	l->1099	m->4	n->12	p->107	s->46	t->25	u->3	v->174	
äm	b->8	d->21	e->1	f->18	j->62	k->2	l->109	m->201	n->231	p->278	r->15	s->79	t->30	v->2	
än	 ->257	,->2	.->4	;->1	a->24	d->1263	f->1	g->272	h->47	i->14	k->423	l->15	n->417	s->451	t->193	v->35	
äp	a->1	n->3	p->24	r->1	
är	 ->3726	!->33	,->115	.->48	:->5	;->1	?->3	a->205	b->1	d->478	e->142	f->281	g->3	h->6	i->41	j->2	k->182	l->83	m->101	n->115	o->4	p->17	r->60	s->175	t->88	u->1	v->70	
äs	 ->3	a->3	b->2	c->2	d->1	e->42	f->1	k->2	n->2	o->1	s->31	t->161	
ät	 ->10	.->1	a->7	e->9	h->1	i->1	o->1	s->2	t->1677	v->11	
äv	 ->1	a->78	d->32	e->322	i->1	j->1	l->3	n->14	s->57	t->4	u->2	
äx	a->11	e->10	l->4	o->1	t->32	
å 	"->1	-->8	1->6	2->5	3->3	4->1	5->3	7->2	8->3	9->2	A->4	B->7	C->2	D->1	E->28	F->2	G->3	H->1	I->9	K->1	M->2	O->1	P->2	R->3	T->1	V->2	a->487	b->117	c->3	d->432	e->372	f->267	g->145	h->86	i->144	j->16	k->153	l->92	m->217	n->93	o->123	p->79	r->77	s->375	t->150	u->62	v->221	y->3	z->2	Ö->2	ä->60	å->22	ö->16	
å,	 ->59	
å.	 ->2	.->1	A->2	B->3	D->16	E->3	F->4	G->2	H->2	I->2	J->10	M->1	N->4	O->3	P->2	S->2	U->1	V->4	Ä->2	
å:	 ->7	
å;	 ->1	
å?	.->1	I->1	J->1	S->1	
åb	a->2	e->1	j->1	ö->11	
åd	 ->18	,->4	.->5	?->1	a->217	d->9	e->730	f->6	g->27	l->7	n->1	r->1	s->49	
åe	l->14	n->136	r->15	t->1	
åf	r->1	ö->10	
åg	 ->43	,->1	.->1	a->605	e->20	i->3	k->2	l->7	n->8	o->639	r->153	s->4	t->2	v->1	å->18	
åh	u->1	ä->7	ö->1	
åj	a->1	
åk	 ->5	.->1	a->10	e->4	i->3	l->40	o->2	r->30	t->2	
ål	 ->102	,->17	-->1	.->17	:->2	a->12	d->27	e->92	f->5	g->1	i->57	k->1	l->474	m->1	n->3	s->28	u->4	v->5	ä->6	
åm	i->30	
ån	 ->633	,->4	.->6	a->93	b->1	d->230	e->2	g->584	i->7	k->3	s->1	t->3	v->9	y->1	
åo	l->1	
åp	e->50	s->1	
år	 ->860	"->1	)->1	,->32	.->42	?->2	a->188	b->5	d->32	e->85	h->7	i->46	k->2	l->10	n->2	s->21	t->155	ö->1	
ås	 ->43	,->1	.->3	:->1	a->4	e->3	i->50	k->10	o->34	s->1	t->746	y->5	
åt	 ->180	"->1	,->5	.->9	a->122	e->287	f->12	g->241	i->4	l->5	m->27	n->7	r->3	s->12	t->155	v->4	
åv	a->2	e->37	i->7	o->2	ä->41	
åz	o->1	
ça	 ->5	
ço	i->1	
èr	e->1	
èt	e->1	
èv	e->3	
é 	-->3	a->3	e->1	f->3	h->1	j->1	k->1	m->1	o->4	p->1	s->5	u->1	ä->1	
é,	 ->1	
éa	v->1	
éb	e->1	é->1	
éc	h->1	
ée	,->1	r->21	
éf	é->1	ö->2	
ék	o->1	
én	 ->38	,->5	.->3	?->1	s->11	
ér	e->1	y->1	
és	 ->1	y->2	
ét	a->1	
éu	n->2	
êt	e->3	s->1	
í 	ä->1	
íe	z->1	
ín	c->1	
ón	 ->5	i->1	
ôn	e->1	
ö 	f->2	i->2	k->1	m->1	s->2	v->1	
ö!	D->1	
ö,	 ->12	
ö-	 ->2	
ö.	D->4	M->1	U->1	V->1	
öa	n->3	r->6	v->1	
öb	e->3	l->2	o->1	r->1	
öc	k->3	
öd	 ->166	,->14	.->44	;->1	?->1	a->19	b->1	d->4	e->151	f->1	g->1	i->15	j->72	m->2	n->2	o->3	p->1	r->9	s->18	v->125	å->5	
öe	n->1	r->4	
öf	a->10	r->4	t->11	ö->4	
ög	 ->21	,->1	a->20	e->34	h->3	l->1	n->4	o->19	r->20	s->29	t->17	
öi	n->1	
öj	a->30	d->24	e->15	l->309	n->2	o->1	s->3	t->4	
ök	 ->12	,->3	a->188	e->29	m->1	n->43	o->6	r->8	s->3	t->20	v->1	
öl	 ->2	,->1	a->2	d->4	j->174	l->25	n->2	
öm	 ->5	,->1	:->1	a->37	b->1	d->4	e->11	i->1	l->2	m->32	n->34	s->9	t->13	v->1	ä->13	å->3	
ön	 ->20	!->1	,->9	.->11	a->19	b->1	d->7	e->7	h->1	i->1	k->4	o->2	s->80	t->5	
öo	m->4	v->1	
öp	 ->2	a->13	e->15	k->1	o->8	p->99	r->4	s->2	t->9	å->1	
ör	 ->4373	"->1	,->32	.->24	:->3	;->1	?->5	a->972	b->229	d->350	e->897	f->136	g->20	h->195	i->43	j->131	k->95	l->161	m->70	n->84	o->83	p->27	r->144	s->1374	t->199	u->85	v->160	ä->74	å->4	ö->10	
ös	 ->12	,->1	.->1	a->67	e->6	g->1	h->44	i->1	k->18	n->52	r->1	s->5	t->294	y->6	
öt	 ->10	.->1	a->20	e->135	f->1	k->3	r->1	s->17	t->40	
öu	t->1	
öv	a->47	d->2	e->747	i->1	l->2	n->12	o->1	r->68	s->29	t->4	ä->10	
öw	 ->1	
öy	 ->1	
öö	w->1	
øn	,->2	
ør	g->2	
üh	r->1	
ün	c->1	
ür	k->1	
üs	s->4	
