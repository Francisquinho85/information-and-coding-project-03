 "A	m->1	t->1	
 "B	i->1	
 "D	e->4	
 "E	U->1	q->1	u->2	
 "J	a->1	
 "K	u->4	v->3	
 "L	o->1	
 "M	i->2	
 "O	l->1	m->1	
 "P	o->1	
 "T	i->2	y->1	
 "U	r->1	
 "a	f->1	l->3	n->3	v->1	
 "b	a->1	
 "c	o->1	
 "d	e->4	ö->1	
 "e	g->1	k->1	n->4	u->3	
 "f	o->1	ö->1	
 "g	e->2	
 "h	e->2	
 "i	n->2	r->1	
 "j	a->1	
 "k	o->2	r->1	u->1	
 "l	ä->3	
 "m	e->1	
 "n	a->1	e->1	o->1	å->1	
 "o	b->1	r->1	v->1	
 "p	a->1	å->1	
 "r	e->5	i->1	
 "s	e->1	h->1	k->1	p->1	v->1	
 "t	i->1	
 "u	t->2	
 "v	a->2	
 "å	t->1	
 "ö	p->1	v->1	
 'V	a->1	
 ("	d->1	
 (1	4->2	9->2	
 (5	7->1	
 (8	0->2	
 (9	6->1	
 (A	5->35	
 (B	5->4	e->1	r->2	
 (C	5->7	E->3	O->1	
 (D	E->1	
 (E	G->1	I->1	L->1	N->23	U->3	
 (F	I->2	P->1	R->12	U->1	
 (H	-->21	o->1	
 (I	C->1	F->1	M->1	n->1	
 (K	O->8	u->2	
 (P	P->1	T->15	
 (S	E->1	P->1	
 (U	t->2	
 (a	r->7	t->1	v->1	
 (d	e->2	
 (e	f->1	l->1	n->2	
 (f	i->4	o->1	ö->3	
 (h	ä->1	
 (i	 ->2	n->2	
 (k	o->4	r->2	
 (m	a->2	e->1	
 (o	c->1	
 (r	e->1	å->1	
 (s	e->1	å->1	
 (t	.->1	y->1	
 (u	n->1	
 (Ö	V->1	s->4	
 (å	t->1	
 , 	a->1	b->1	d->1	m->1	v->1	
 - 	"->1	'->1	,->1	1->26	2->1	3->1	6->1	8->1	A->2	C->21	D->1	E->1	H->1	K->2	P->1	R->3	S->2	a->44	b->4	c->1	d->58	e->26	f->23	g->5	h->15	i->28	j->16	k->12	l->5	m->23	n->14	o->73	p->8	r->6	s->53	t->10	u->11	v->23	Ö->2	ä->17	å->2	ö->5	
 -(	E->1	
 -,	 ->9	
 -e	r->1	
 -o	r->3	
 0 	p->1	
 00	0->25	8->2	
 01	1->1	
 05	5->1	
 06	5->1	
 1 	0->2	4->1	f->1	i->1	j->6	m->3	o->7	p->4	s->1	u->2	
 1,	 ->5	2->2	4->1	
 1-	2->1	o->4	r->5	s->2	
 1.	J->1	
 1/	3->1	
 10	 ->16	,->1	.->1	0->9	5->2	
 11	 ->6	,->4	.->6	0->1	5->1	
 12	 ->8	,->4	.->6	/->3	0->1	3->1	4->3	5->1	6->1	
 13	 ->13	,->2	.->2	0->1	3->1	8->1	
 14	 ->13	,->1	0->1	3->1	
 15	 ->12	,->2	.->2	0->2	8->4	
 16	 ->7	)->1	,->1	4->1	6->1	7->3	
 17	 ->5	,->2	.->2	0->1	4->1	6->2	
 18	 ->8	,->1	0->1	
 19	 ->5	.->1	1->1	2->1	3->2	4->3	5->3	6->7	7->2	8->6	9->192	
 2 	-->1	0->1	4->1	b->2	d->1	e->1	i->4	m->1	o->3	p->3	s->1	
 2,	 ->5	4->1	6->1	8->1	
 2-	o->2	s->1	
 2.	1->1	2->1	D->1	M->1	
 20	 ->16	,->1	.->1	0->97	1->2	
 21	 ->7	.->2	:->1	
 22	 ->2	,->4	.->1	6->1	
 23	 ->2	,->1	
 24	 ->5	5->1	8->1	
 25	 ->12	.->1	0->1	5->4	
 26	 ->6	2->1	
 27	 ->6	,->1	
 28	 ->4	,->2	0->5	:->1	
 29	 ->4	,->1	9->2	
 3 	0->2	f->1	j->1	m->1	o->2	p->2	
 3,	 ->1	8->2	
 3-	4->1	l->2	
 3.	1->1	8->1	I->1	
 30	 ->10	,->1	0->1	
 31	 ->6	4->1	
 32	 ->1	,->2	.->1	
 33	 ->7	2->1	
 34	 ->4	,->1	.->1	4->1	
 35	 ->6	.->1	0->1	
 36	 ->1	,->1	7->1	
 37	 ->3	,->2	.->1	/->1	0->1	
 38	 ->4	,->1	:->1	
 39	 ->3	,->1	
 3:	 ->1	
 4 	0->1	c->1	e->1	i->5	j->2	l->1	o->1	p->1	
 4,	 ->4	
 4.	2->1	I->2	J->1	
 40	 ->11	,->1	0->6	
 41	 ->4	0->1	
 42	 ->4	
 43	 ->1	.->1	
 44	 ->3	
 45	 ->4	,->1	.->4	
 46	 ->2	2->1	
 47	 ->1	
 48	 ->5	
 5 	0->5	f->1	g->1	m->3	o->1	v->1	å->1	
 5,	 ->3	5->1	8->1	
 5.	4->1	E->1	
 50	 ->7	,->1	-->3	0->1	
 51	9->1	
 52	 ->1	0->2	2->1	
 53	 ->1	
 54	0->1	
 55	 ->2	
 56	 ->1	,->1	
 57	,->1	
 5b	 ->1	-->1	.->1	
 6 	d->1	f->1	i->6	m->1	o->7	
 6,	 ->2	0->1	
 6.	S->1	
 60	 ->2	-->1	0->1	
 62	 ->1	
 67	 ->1	
 68	 ->1	5->1	
 7 	-->1	d->1	f->1	g->1	i->8	l->1	n->1	o->2	p->2	
 7)	.->1	
 7,	 ->5	2->1	4->1	
 7.	F->1	
 70	 ->2	0->4	
 73	,->1	
 75	 ->3	
 76	 ->1	
 77	 ->1	
 79	/->1	
 8 	4->1	b->1	f->1	o->3	r->1	t->1	ä->1	
 8,	 ->2	
 80	 ->14	
 81	 ->6	.->10	
 82	 ->2	)->1	,->4	.->1	
 83	 ->1	
 85	 ->4	
 86	 ->3	
 87	,->1	.->2	
 88	 ->3	/->2	
 89	 ->2	
 9 	d->1	f->3	i->1	m->3	
 9,	 ->2	
 9.	1->1	
 90	 ->5	-->1	
 91	 ->1	
 92	/->1	
 93	 ->1	/->1	
 94	 ->3	,->1	/->3	
 95	 ->4	/->1	
 96	/->5	
 97	.->1	/->1	
 98	 ->1	
 : 	P->1	
 A.	 ->1	
 AB	B->3	C->1	
 AD	R->1	
 AK	T->1	
 Ac	t->1	
 Ad	a->1	e->1	o->2	r->1	
 Af	r->4	
 Ag	r->1	u->1	
 Ah	e->7	
 Ai	d->1	
 Ak	k->3	
 Al	a->2	b->4	e->2	g->1	i->1	l->5	p->1	s->4	t->16	
 Am	e->1	o->7	s->36	
 An	g->1	k->1	l->1	m->1	n->1	t->1	v->1	
 Ap	a->1	
 Ar	a->2	b->1	i->4	t->1	
 As	i->2	s->2	t->1	
 At	a->2	l->3	t->3	
 Au	s->1	t->1	v->1	
 Av	 ->2	f->1	i->1	s->1	
 Az	o->2	
 B 	o->1	t->1	
 BN	I->7	P->9	
 BP	,->1	
 BR	Å->1	
 BS	E->6	
 Ba	l->8	n->1	r->29	s->3	
 Be	l->9	r->39	s->2	t->1	
 Bi	s->6	
 Bl	a->2	o->1	
 Bo	e->1	l->1	n->1	r->2	u->6	w->4	
 Br	a->4	e->8	i->1	o->9	u->1	y->16	
 Bu	d->1	l->1	s->2	
 By	r->3	
 C.	 ->2	
 C4	-->6	
 C5	-->15	
 CE	C->1	N->10	
 CS	U->2	
 Ca	d->6	m->2	n->5	s->2	u->1	v->1	
 Ce	n->11	r->1	y->1	
 Ch	a->1	i->1	
 Cl	i->1	
 Co	c->2	l->1	n->2	r->1	s->9	u->1	x->4	
 Cr	e->2	
 Cu	r->1	s->1	x->1	
 Cy	p->1	
 D 	k->1	
 DD	R->1	
 Da	 ->3	g->2	l->6	m->3	n->25	r->1	v->3	
 De	 ->19	l->3	m->2	n->28	r->1	s->4	t->88	u->1	
 Di	m->5	r->2	
 Do	m->1	r->1	
 Du	b->7	h->1	i->3	t->1	
 Dä	r->7	
 Då	 ->2	
 Dí	e->1	
 Dü	h->1	
 E-	k->1	
 EC	H->3	
 ED	D->3	
 EE	G->3	
 EG	 ->1	-->48	.->1	:->3	
 EI	F->1	
 EK	S->5	
 EL	D->3	
 EM	U->6	
 EU	 ->37	,->5	-->39	.->11	:->44	?->1	G->1	
 Ec	e->1	
 Ed	i->1	
 Ef	t->11	
 Eg	y->2	
 Eh	u->2	
 Ei	e->1	
 Ek	o->3	
 El	i->1	l->3	m->2	s->1	
 Em	i->1	
 En	 ->6	d->1	l->5	
 Eq	u->9	
 Er	a->1	i->25	k->2	t->1	
 Et	i->3	t->2	
 Eu	r->794	
 Ev	a->7	
 Ex	x->3	
 FB	I->1	
 FE	O->2	
 FM	I->1	
 FN	,->1	-->1	.->1	:->8	
 FP	Ö->14	
 FR	Å->1	
 Fa	c->1	r->1	
 Fe	i->2	
 Fi	n->7	r->1	s->4	
 Fl	a->2	o->16	é->1	
 Fo	U->2	g->1	l->3	n->1	r->2	
 Fr	a->48	i->2	u->11	ä->2	å->2	
 Fu	n->1	
 Fä	s->1	
 Få	r->2	
 Fö	l->1	r->70	
 GA	-->1	S->1	
 GU	E->2	S->1	
 Ga	l->3	m->3	r->5	z->6	
 Ge	m->2	n->13	
 Gi	l->2	n->1	
 Go	e->1	l->12	m->1	n->1	o->1	r->1	t->1	
 Gr	a->9	e->12	o->3	u->8	ö->2	
 Gu	a->1	i->1	l->1	s->1	t->2	
 Gö	t->1	
 Ha	a->1	d->1	g->1	i->36	m->1	n->3	r->4	t->2	v->1	
 He	b->1	d->2	i->1	l->21	n->1	r->30	
 Hi	c->1	l->1	m->1	t->7	
 Ho	l->3	n->1	
 Hu	h->1	l->24	r->1	
 Hä	n->2	r->3	
 Hå	l->1	
 I 	-->1	S->1	T->1	b->4	d->11	e->4	g->1	l->1	m->2	o->2	r->1	s->3	u->1	
 I-	p->1	
 IC	E->3	
 II	 ->3	,->1	-->2	I->2	
 IM	O->2	
 IN	T->4	
 IR	A->1	
 IS	P->1	
 IV	 ->3	
 IX	 ->1	,->1	
 Il	e->1	
 Im	b->3	
 In	d->5	g->6	i->1	t->22	
 Ir	l->21	
 Is	a->2	l->1	r->36	t->1	
 It	a->17	
 Iz	q->1	
 Ja	,->2	c->5	g->140	n->1	p->3	v->1	
 Je	a->1	r->2	
 Jo	n->15	r->3	s->1	
 Ju	g->1	n->1	
 Jä	m->1	
 Jö	r->14	
 Ka	l->3	n->5	r->11	s->1	u->4	z->1	
 Kf	o->1	
 Ki	n->31	r->5	
 Ko	c->14	m->12	n->2	r->2	s->60	u->12	
 Ku	l->11	m->1	n->1	
 Kv	i->1	ä->1	
 Ky	o->7	
 Kä	n->1	r->3	
 Kö	l->2	p->1	
 LT	C->1	
 La	 ->1	a->7	m->7	n->33	p->2	
 Le	a->5	d->1	i->8	o->1	
 Li	b->8	i->3	k->2	l->1	s->8	t->1	
 Ll	o->1	
 Lo	i->2	m->2	n->4	r->4	t->2	u->1	y->2	
 Lu	t->1	x->6	
 Ly	n->3	
 Lå	t->12	
 Lö	ö->1	
 MA	R->1	
 Ma	a->6	c->1	d->6	i->1	l->5	n->3	r->13	
 Mc	C->1	N->5	
 Me	d->5	l->17	n->15	x->1	
 Mi	c->1	d->2	n->7	s->1	t->4	
 Mo	n->19	r->9	s->1	u->9	
 Mu	l->1	
 Mü	n->1	
 Na	n->1	p->1	r->1	t->9	
 Ne	d->9	j->1	w->1	
 Ni	 ->6	e->5	k->2	
 No	g->1	i->1	r->3	
 Nu	 ->1	
 Ny	a->2	t->1	
 Nä	r->13	s->1	
 Nå	g->1	
 OC	H->1	
 OF	S->1	
 OL	A->15	F->1	
 OM	 ->1	
 OS	S->1	
 Ob	e->1	
 Oc	h->5	
 Of	f->2	
 Oi	l->1	
 Ol	i->1	j->1	y->1	
 Om	 ->5	a->1	
 On	e->1	
 Or	a->1	
 Os	l->3	m->1	
 Ou	v->1	
 Oz	 ->1	,->1	
 PP	E->12	
 PR	-->1	
 PS	E->4	
 PV	C->3	
 Pa	c->3	d->2	k->5	l->26	p->2	r->7	t->23	y->2	
 Pe	a->1	i->2	k->1	t->2	
 Pl	a->2	o->1	
 Po	e->5	h->1	l->2	m->1	n->1	o->1	r->24	w->3	
 Pr	e->1	i->1	o->29	í->1	
 Pu	r->1	
 På	 ->4	s->1	
 Pé	t->1	
 Qu	e->1	
 RE	P->2	
 RI	N->2	
 Ra	c->2	f->3	n->4	p->11	s->1	
 Re	a->1	d->8	g->1	p->1	v->2	
 Rh	ô->1	
 Ri	c->3	i->2	k->1	o->1	
 Ro	b->1	i->1	j->1	m->4	o->1	t->7	v->2	y->1	
 Ru	i->1	s->1	
 Ry	s->4	
 Rå	d->6	
 Ré	u->2	
 SE	K->3	M->1	
 SO	L->1	
 SP	Ö->1	
 SS	 ->1	
 Sa	g->1	i->1	l->1	m->15	n->4	v->7	
 Sc	h->35	
 Se	a->4	b->1	d->4	g->2	i->5	
 Sh	a->5	e->5	
 Si	m->1	
 Sj	u->1	ä->1	ö->4	
 Sk	o->5	u->1	ä->1	
 Sl	o->1	
 So	a->1	c->1	k->1	l->6	m->9	u->1	
 Sp	a->7	e->2	
 Sr	i->3	
 St	.->1	a->2	o->17	r->6	ö->1	
 Su	a->1	d->2	
 Sv	e->7	
 Sw	o->3	
 Sy	d->5	r->22	
 Sá	n->1	
 Sã	o->2	
 Så	 ->2	
 Sö	d->2	
 TV	 ->1	-->3	
 Ta	c->9	d->4	i->1	l->1	m->22	n->2	u->1	
 Te	r->3	s->1	x->2	
 Th	e->19	y->4	
 Ti	b->19	d->1	l->8	
 To	d->1	m->3	r->3	t->6	
 Tr	a->1	e->1	i->1	o->1	
 Ts	a->3	
 Tu	r->37	
 Ty	s->20	
 Tå	g->1	
 UC	K->1	L->1	
 UE	N->1	
 UN	I->1	M->3	
 US	A->10	D->1	
 Ul	s->1	
 Un	d->6	i->3	
 Up	p->1	
 Ur	b->1	q->1	s->1	
 Ut	n->1	s->2	v->1	
 Uz	b->2	
 V 	-->1	
 VD	 ->1	
 VI	 ->1	I->2	
 Va	d->9	l->6	n->3	p->1	r->5	t->3	
 Ve	l->1	m->3	n->4	r->3	
 Vi	 ->39	,->1	c->1	d->2	l->1	s->1	t->7	v->1	
 Vl	a->1	
 Vo	d->1	l->1	
 Vä	r->3	s->4	
 Vå	r->5	
 WT	O->1	
 Wa	f->2	l->15	s->3	
 We	b->1	s->1	
 Wi	d->1	e->9	l->1	
 Wo	g->18	
 Wu	l->2	r->3	
 Wy	e->3	n->1	
 X 	o->1	
 XX	V->2	
 Ya	s->1	
 Yo	r->1	
 Ze	e->2	
 Zi	m->1	
 [K	O->2	
 [S	E->1	
 a 	p->3	
 a)	 ->2	
 ab	s->45	
 ac	c->57	q->1	
 ad	 ->3	d->1	e->5	j->2	m->23	r->1	v->5	
 af	f->4	
 ag	e->43	g->1	i->1	r->2	
 ai	d->5	
 aj	o->1	
 ak	t->80	u->1	
 al	-->1	b->9	d->29	i->1	k->3	l->1028	t->12	
 am	b->28	e->11	
 an	 ->10	a->51	b->5	d->340	f->16	g->76	h->4	i->5	k->5	l->58	m->28	n->131	o->12	p->12	s->654	t->193	v->159	
 ap	p->8	r->4	
 ar	a->8	b->407	g->16	k->2	m->4	r->10	t->107	v->4	
 as	"->1	p->30	s->3	t->1	y->21	
 at	l->1	o->4	t->6142	
 au	c->1	k->6	t->9	
 av	 ->2672	,->5	.->7	a->2	b->11	d->8	e->2	f->26	g->85	h->5	i->4	k->3	l->16	m->1	p->1	r->5	s->275	t->56	u->1	v->40	
 ax	e->1	l->1	
 b)	 ->2	
 ba	c->2	d->5	g->2	i->1	k->57	l->25	n->20	r->247	s->24	x->1	
 be	 ->19	a->32	b->2	d->92	f->150	g->158	h->317	i->1	k->142	l->36	m->17	n->5	o->1	r->202	s->451	t->593	u->3	v->113	
 bi	b->13	d->109	e->2	f->3	g->1	l->215	n->14	o->9	s->20	t->5	
 bj	u->2	
 bl	.->27	a->57	e->15	i->264	o->13	u->4	y->8	å->1	
 bo	 ->2	e->1	g->1	j->1	k->5	l->5	m->10	n->2	r->127	s->14	t->13	v->2	
 br	a->87	e->26	i->80	o->59	u->12	y->14	ä->14	å->21	ö->4	
 bu	d->114	r->1	s->1	
 by	g->50	r->34	t->3	x->1	
 bä	r->30	s->42	t->75	
 bå	d->69	t->9	
 bé	b->1	
 bö	c->3	d->1	j->2	r->322	t->1	
 c 	i->1	
 c)	 ->1	
 ca	 ->1	.->1	l->1	n->3	p->10	s->1	
 ce	m->2	n->55	r->5	
 ch	a->15	e->6	o->5	
 ci	r->9	t->8	v->19	
 co	m->3	n->3	p->1	r->5	s->5	
 cr	i->1	
 d)	 ->1	
 da	 ->6	g->328	m->44	n->24	t->20	
 de	 ->1753	,->4	a->1	b->167	c->41	f->35	g->2	l->340	m->316	n->2284	p->5	r->92	s->491	t->3848	
 di	a->31	e->2	f->5	g->2	k->5	l->3	m->12	o->2	p->11	r->212	s->180	t->7	v->4	
 dj	u->44	ä->9	
 do	c->61	g->5	k->39	l->9	m->89	
 dr	a->100	i->28	o->7	u->5	y->4	å->1	ö->8	
 du	 ->6	b->15	g->1	k->1	m->8	n->1	s->1	
 dv	s->45	
 dy	k->7	l->3	n->5	r->7	s->1	
 dä	c->1	m->2	r->518	
 då	 ->148	,->2	.->1	?->1	l->19	v->1	
 dö	 ->1	d->20	e->1	l->10	m->11	p->4	r->11	t->3	
 e)	 ->1	
 e-	m->1	
 e.	d->1	
 ec	u->2	
 ed	 ->1	e->1	
 ef	f->129	t->358	
 eg	e->124	n->44	o->2	
 ej	 ->11	,->1	.->2	
 ek	o->260	v->1	
 el	-->6	e->20	i->3	l->323	m->1	o->2	v->2	
 em	b->3	e->64	i->2	o->55	
 en	 ->2427	,->2	.->1	a->49	b->30	d->122	e->98	g->28	h->85	i->10	k->47	l->122	o->32	s->61	t->11	v->6	
 ep	o->4	
 er	 ->136	,->25	.->8	:->2	a->37	b->19	f->31	h->10	i->13	k->39	s->22	t->38	ö->1	
 et	 ->1	a->16	c->6	i->2	n->11	t->1368	
 eu	r->391	
 ev	e->21	i->3	
 ex	 ->6	a->34	c->5	e->116	i->19	k->3	p->58	t->37	
 f.	d->2	
 fa	b->1	c->4	d->1	i->1	k->133	l->163	m->15	n->26	r->147	s->120	t->79	u->1	v->1	x->1	
 fe	b->16	d->8	l->35	m->55	n->3	
 fi	c->26	e->3	l->6	n->470	r->1	s->40	
 fj	o->12	ä->11	
 fl	a->17	e->150	i->3	o->7	y->38	ä->1	ö->1	
 fo	d->6	g->2	k->5	l->77	n->26	r->372	s->2	t->4	
 fr	a->692	e->69	i->138	o->6	u->86	y->2	ä->140	å->1253	
 fu	l->97	n->103	s->8	t->1	
 fy	l->7	r->28	s->9	
 fä	d->1	l->10	n->1	r->9	s->12	
 få	 ->206	,->3	.->3	g->9	n->5	r->186	s->1	t->58	
 fö	d->7	g->2	l->125	n->1	r->6369	t->3	
 ga	g->7	l->3	m->32	n->26	r->91	s->1	t->1	v->12	
 ge	 ->128	.->1	d->2	m->379	n->463	o->10	r->64	s->16	t->21	
 gi	c->8	f->2	g->5	l->16	s->1	v->48	
 gj	o->112	
 gl	a->26	e->1	o->12	u->1	ä->40	ö->19	
 gn	u->2	ä->1	
 go	d->236	l->1	t->19	
 gr	a->131	e->9	i->8	o->3	u->394	y->1	ä->60	å->2	ö->19	
 gu	d->2	l->2	m->1	v->1	
 gy	n->11	
 gä	c->1	l->404	r->33	
 gå	 ->71	.->2	n->132	r->92	t->20	
 gö	m->4	r->434	
 ha	 ->190	,->1	.->1	d->85	f->37	k->1	l->25	m->40	n->488	p->1	r->1706	s->1	t->4	v->44	
 he	b->1	d->6	j->2	k->2	l->389	m->38	n->27	r->209	s->1	t->8	
 hi	e->4	g->1	n->45	s->33	t->63	
 hj	ä->117	
 ho	b->2	c->2	m->4	n->57	p->100	r->6	s->50	t->39	
 hu	g->3	m->9	n->11	r->212	s->7	v->47	
 hy	c->5	g->2	l->2	p->2	r->1	s->9	
 hä	f->1	l->27	m->3	n->208	r->301	s->1	v->30	
 hå	l->149	n->2	r->28	v->1	
 hö	g->126	j->17	l->6	n->1	r->79	s->1	
 i 	"->1	-->1	1->1	2->3	A->29	B->30	C->9	D->14	E->201	F->30	G->13	H->15	I->21	J->1	K->45	L->21	M->26	N->6	O->2	P->12	R->4	S->40	T->41	U->5	V->3	W->5	Y->1	a->142	b->73	c->3	d->713	e->232	f->346	g->65	h->80	i->13	j->16	k->112	l->41	m->159	n->36	o->57	p->102	r->98	s->404	t->54	u->82	v->173	y->4	z->2	Ö->38	ä->14	å->17	ö->21	
 i,	 ->2	
 i.	A->1	D->2	N->1	S->2	
 ia	k->8	n->1	
 ib	e->1	l->19	
 ic	k->34	
 id	a->1	e->30	r->4	é->33	
 if	a->2	r->35	
 ig	e->46	n->4	å->7	
 ih	j->1	o->10	ä->1	å->16	
 ik	a->1	r->4	
 il	l->17	s->2	
 im	a->2	m->8	p->16	
 in	 ->91	,->4	b->34	c->8	d->72	e->3	f->279	g->194	h->8	i->69	k->39	l->98	n->259	o->283	p->1	r->185	s->352	t->1957	v->74	ö->1	
 ir	a->1	l->8	o->2	r->7	
 is	 ->2	c->1	o->7	r->19	t->1	ä->2	
 it	a->17	u->20	
 iv	e->2	ä->3	
 ja	 ->7	,->5	g->1088	k->3	n->16	p->1	
 je	t->1	
 jo	b->4	n->1	r->69	u->2	
 ju	 ->70	,->2	b->1	d->3	l->13	n->13	r->45	s->104	v->1	
 jä	m->55	r->17	t->1	
 ka	b->4	d->3	l->33	m->88	n->863	o->2	p->28	r->27	s->4	t->77	
 ke	d->4	l->1	m->6	
 ki	d->1	l->5	n->9	
 kl	.->21	a->173	i->14	o->10	y->5	
 km	 ->2	,->1	.->1	
 kn	a->16	i->1	o->1	u->8	y->8	ä->2	
 ko	a->12	d->5	f->1	h->1	k->1	l->209	m->2076	n->833	o->1	p->7	r->114	s->101	
 kr	a->142	e->9	i->123	o->5	y->4	ä->151	å->2	ö->1	
 ku	b->1	l->112	m->2	n->314	r->8	s->27	
 kv	a->84	e->3	i->62	o->11	ä->11	
 ky	l->3	
 kä	l->9	m->5	n->108	r->110	
 kö	k->1	l->5	n->4	p->6	r->8	t->2	
 l'	e->1	
 la	 ->1	b->3	d->17	g->219	n->170	p->3	r->5	s->7	w->2	
 le	 ->2	d->230	g->33	j->1	k->2	m->2	t->11	v->36	
 li	b->26	c->1	d->11	g->76	k->159	l->5	n->20	s->12	t->72	v->124	
 lj	u->13	
 lo	b->5	c->2	g->13	j->5	k->42	p->2	s->2	t->4	v->18	
 lu	c->5	d->2	f->2	g->6	k->1	n->1	r->2	t->2	
 ly	c->59	d->5	f->8	k->1	s->35	
 lä	c->4	g->163	k->5	m->102	n->216	r->20	s->19	t->42	x->2	
 lå	g->14	n->116	s->3	t->50	
 lö	f->11	j->3	k->1	n->12	p->20	r->1	s->93	v->1	
 m.	m->1	
 ma	g->2	i->5	j->46	k->45	l->3	n->665	r->207	s->17	t->31	x->8	
 me	d->2304	g->1	k->9	l->199	n->465	r->203	s->44	t->27	
 mi	d->1	g->235	k->4	l->282	n->498	r->1	s->80	t->70	x->1	
 mj	u->1	
 mo	b->7	d->65	g->2	m->1	n->29	r->56	t->338	
 mu	l->9	n->8	r->1	s->6	t->1	
 my	c->452	g->1	l->1	n->110	t->1	
 mä	k->3	n->166	r->23	t->4	
 må	 ->3	h->5	l->152	n->248	r->1	s->696	t->5	
 mö	b->1	d->2	j->281	r->7	t->31	
 na	c->6	i->2	k->1	m->16	r->6	t->300	z->8	
 ne	d->50	g->26	j->5	k->5	o->2	p->5	r->8	u->2	
 ni	 ->222	,->11	.->1	m->1	o->14	v->67	
 nj	u->1	
 no	g->41	l->3	m->3	n->2	r->53	t->29	v->11	
 nr	 ->29	
 nu	 ->206	,->6	.->4	:->1	?->1	l->2	m->7	n->1	v->45	
 ny	 ->39	a->169	b->2	c->7	d->1	e->2	f->2	h->12	k->3	l->30	n->6	p->1	s->14	t->77	v->1	å->1	
 nä	m->126	r->470	s->48	t->17	
 nå	 ->18	b->2	d->1	g->504	r->2	t->7	
 nö	d->127	j->26	t->6	
 oa	c->31	k->1	n->6	v->12	
 ob	a->6	e->64	j->1	l->14	s->2	
 oc	h->4559	k->590	
 od	d->1	e->1	i->1	j->2	u->1	
 oe	f->1	g->5	k->1	n->8	r->13	t->1	
 of	 ->1	a->2	e->1	f->110	r->4	t->54	u->2	ö->21	
 og	e->2	r->2	y->1	
 oh	j->1	ä->1	ö->1	
 oi	g->1	n->6	
 oj	ä->7	
 ok	l->14	o->2	r->2	t->8	u->3	ä->2	
 ol	a->4	i->120	j->40	o->1	y->46	ä->3	ö->2	
 om	 ->1775	"->1	)->1	,->21	.->26	I->1	b->19	d->4	e->21	f->90	g->5	h->1	i->1	k->15	l->3	m->1	o->3	p->9	r->258	s->65	t->1	v->17	ö->16	
 on	d->6	e->1	s->5	t->2	ö->11	
 op	a->2	e->12	i->4	p->7	r->3	t->8	
 or	d->309	e->4	g->69	i->15	k->3	m->2	o->87	s->29	t->2	w->1	ä->11	
 os	a->1	s->324	t->3	v->6	y->1	ä->8	å->1	
 ot	a->1	i->17	j->1	r->3	v->3	y->4	ä->1	å->1	
 ou	m->4	n->6	t->3	
 ov	a->7	e->1	i->4	ä->4	
 oä	n->4	
 oö	n->1	v->6	
 p.	g->1	
 pa	k->3	l->12	p->5	r->534	s->18	t->3	
 pe	a->1	d->2	k->19	l->8	n->72	r->218	s->6	t->1	
 ph	a->1	t->1	
 pi	l->3	o->1	r->1	
 pl	a->131	e->9	i->6	u->4	ä->2	å->1	ö->4	
 po	e->1	l->341	o->1	p->5	r->75	s->82	t->5	ä->12	
 pr	a->45	e->122	i->202	o->629	ä->4	ö->7	
 ps	y->1	
 pu	b->7	m->2	n->171	r->1	
 py	r->1	
 på	 ->1764	,->16	.->16	:->3	?->2	b->12	d->1	f->4	g->21	l->3	m->30	p->49	s->28	t->16	v->39	
 qu	a->2	o->2	
 ra	d->42	k->7	m->91	n->15	p->98	s->29	t->20	
 re	a->50	c->2	d->191	e->4	f->138	g->655	h->1	j->3	k->47	l->37	m->1	n->40	p->31	s->356	t->15	v->36	
 ri	d->1	g->5	k->179	m->19	n->6	s->86	
 ro	 ->1	,->2	c->1	l->65	m->5	p->3	s->4	t->2	
 ru	b->4	i->1	l->6	m->32	n->10	s->5	t->9	
 ry	c->1	g->4	k->8	m->1	s->3	
 rä	c->34	d->28	k->56	t->491	
 rå	d->380	g->1	k->1	o->1	t->1	
 ré	f->1	
 rö	d->3	r->96	s->120	t->5	v->1	
 s.	k->4	
 sa	 ->1	d->75	f->1	g->49	k->122	l->2	m->686	n->40	t->32	
 sc	e->6	h->1	i->1	o->1	
 se	 ->159	d->102	g->20	i->2	k->68	l->1	m->5	n->106	p->16	r->99	s->16	t->49	x->24	
 si	d->81	f->17	g->406	k->27	m->3	n->306	s->57	t->220	
 sj	u->32	ä->192	ö->20	
 sk	a->963	e->83	i->84	j->25	o->45	r->74	u->505	y->113	ä->62	å->2	ö->25	
 sl	a->40	i->4	o->4	u->182	ä->14	å->15	ö->4	
 sm	a->1	i->5	u->5	ä->4	å->67	
 sn	a->137	e->12	ä->2	å->1	ö->1	
 so	 ->1	c->203	f->1	l->34	m->3392	p->1	r->12	v->1	
 sp	a->20	e->153	i->1	l->3	o->7	r->24	ä->13	å->8	ö->4	
 sr	i->1	
 st	a->384	e->43	i->27	o->332	r->311	u->25	y->38	ä->245	å->284	ö->511	
 su	b->38	c->5	d->1	m->10	n->5	p->1	s->1	t->1	v->17	
 sv	a->96	e->6	ä->2	å->93	
 sy	d->4	f->68	m->18	n->120	r->8	s->222	
 sä	g->252	k->243	l->8	m->10	n->20	r->159	s->1	t->309	
 så	 ->478	,->6	.->4	:->1	d->163	g->7	h->1	l->44	n->3	r->2	s->31	t->1	v->43	
 sö	d->6	k->9	n->8	r->10	
 t.	e->19	o->7	
 ta	 ->220	.->1	?->1	b->1	c->144	g->77	k->10	l->608	n->82	p->3	r->65	s->33	x->4	
 te	a->1	c->11	k->45	l->6	m->8	n->12	o->2	r->32	x->35	
 th	e->3	
 ti	b->9	d->252	g->3	l->2539	m->9	n->3	o->16	s->2	t->23	
 tj	a->1	o->2	u->4	ä->119	
 to	b->2	g->29	l->39	m->4	n->23	p->12	r->19	t->34	x->1	
 tr	a->150	e->149	i->2	o->240	u->5	y->12	ä->46	å->8	ö->6	
 tu	f->2	l->2	m->3	n->22	r->39	s->9	
 tv	e->34	i->69	u->11	ä->18	å->132	
 ty	 ->12	c->77	d->110	g->1	n->11	p->41	s->25	v->29	
 tä	c->14	m->3	n->74	p->4	r->1	t->4	v->3	
 tå	g->5	l->3	
 tö	m->1	
 u-	l->1	
 ul	t->3	
 um	g->1	
 un	d->572	g->29	i->440	
 up	p->1011	
 ur	 ->42	a->11	b->1	h->4	m->1	s->38	v->13	
 ut	 ->95	,->20	.->18	:->1	?->2	a->360	b->73	d->1	e->30	f->102	g->109	h->2	i->16	j->5	k->22	l->19	m->53	n->44	o->16	p->5	r->44	s->215	t->201	v->364	ö->40	
 va	c->9	d->239	g->4	k->14	l->95	n->48	p->15	r->895	t->26	
 ve	c->40	d->13	k->4	l->7	m->18	n->1	r->353	t->209	
 vi	 ->1634	,->16	.->1	?->1	a->12	c->13	d->322	f->1	g->2	k->352	l->1093	n->23	r->4	s->343	t->55	
 vo	l->7	n->18	r->29	t->4	
 vr	a->4	e->1	i->1	ä->1	
 vu	n->3	x->3	
 vä	c->17	d->10	g->108	k->2	l->186	n->88	p->2	r->137	s->31	v->4	x->34	
 vå	g->9	l->13	n->2	r->398	
 vö	r->1	
 wa	l->1	
 we	b->1	
 wo	r->1	
 yn	g->2	
 yp	p->2	
 yr	k->20	
 yt	a->1	l->2	t->131	
 zi	g->4	
 zo	n->4	
 º 	C->1	
 Äm	n->1	
 Än	d->1	n->2	
 Är	 ->1	a->2	
 Äv	e->11	
 Å 	P->1	k->1	s->1	
 År	l->1	
 Åt	g->3	
 Îl	e->1	
 ÖV	P->4	
 Öp	p->1	
 Ös	t->82	
 äc	k->1	
 äg	a->36	d->1	e->5	g->1	n->28	t->9	
 äk	t->1	
 äl	d->7	s->2	
 äm	b->7	n->29	
 än	 ->186	,->1	.->1	d->363	g->1	n->77	t->20	
 är	 ->2566	,->13	.->9	:->5	?->1	a->26	e->18	l->8	o->1	
 ät	e->1	
 äv	e->275	
 å 	P->1	a->7	d->3	e->11	m->2	r->1	u->1	
 åb	e->1	
 åh	ö->1	
 åk	l->37	t->1	
 ål	a->3	d->9	i->5	ä->5	
 ån	y->1	
 år	 ->132	,->18	.->27	a->1	e->70	h->7	l->8	s->16	t->5	
 ås	a->4	i->50	k->2	t->25	y->5	
 åt	 ->80	,->2	.->2	a->54	e->250	f->12	g->218	m->27	n->1	s->5	t->6	
 åv	i->1	
 öa	r->6	
 öb	o->1	
 öd	e->13	
 ög	a->1	o->19	
 ök	a->106	n->18	
 öl	 ->1	
 öm	 ->1	m->1	s->5	t->1	
 ön	 ->1	s->63	
 öp	p->98	
 ör	e->8	o->3	
 ös	t->59	
 öv	a->1	e->602	n->5	r->65	
! 1	9->1	
! A	l->2	t->1	v->3	
! B	e->3	l->1	
! C	e->1	
! D	a->1	e->52	i->1	ä->1	í->1	
! E	U->1	f->4	n->1	r->2	t->1	u->7	
! F	r->3	å->1	ö->16	
! G	e->1	o->1	r->3	
! H	e->1	i->1	
! I	 ->18	n->2	
! J	a->110	o->1	ä->1	
! K	a->1	o->5	
! L	i->2	å->9	
! M	a->1	e->1	i->5	
! N	i->5	u->1	ä->7	å->1	
! O	l->1	m->2	
! P	P->1	a->1	r->1	å->3	
! R	e->1	o->1	å->2	
! S	c->1	e->3	k->1	o->7	t->1	
! T	a->3	h->1	i->7	o->1	r->1	
! U	n->4	p->1	r->1	t->2	
! V	a->5	i->23	å->3	
! Ä	n->1	v->9	
! Å	 ->3	r->1	
! Ö	s->1	
!".	D->1	
!"D	e->1	
!"J	a->1	
!"O	m->1	
!(P	a->1	
!. 	(->1	
!.(	N->1	
!.H	e->1	
!Al	l->2	
!Am	s->1	
!An	d->1	
!Av	 ->1	
!De	 ->3	n->3	t->14	
!Dä	r->1	
!Ef	t->2	
!En	 ->1	
!Er	i->1	
!Eu	r->1	
!Fr	u->3	
!Fö	r->2	
!Ge	n->1	
!Ha	n->1	
!He	r->9	
!Hä	r->1	
!I 	d->1	
!Ja	g->18	
!Ku	l->1	
!Le	d->1	
!Lå	t->1	
!Me	d->1	n->4	
!Mi	n->2	
!My	c->1	
!Mä	n->1	
!Ni	 ->1	
!Nä	r->3	
!Om	 ->2	
!Pr	e->1	
!Rö	s->1	
!Sa	n->1	
!Sk	a->1	
!Ta	c->1	
!Ti	l->3	
!Tr	o->1	
!Tv	ä->1	
!Un	d->1	
!Vi	 ->5	
!Äv	e->2	
" (	s->1	
" -	 ->1	
" a	l->1	t->1	v->1	
" b	i->1	
" e	t->1	
" f	r->1	ö->1	
" g	e->1	ö->1	
" h	a->1	
" i	 ->1	
" m	e->2	å->2	
" o	c->6	
" p	å->1	
" s	k->1	o->8	
" t	i->2	
" v	a->1	
" Ä	r->1	
" ä	r->1	
"!I	 ->1	
"),	 ->1	
", 	"->1	a->1	b->1	d->4	e->1	f->1	i->1	m->1	o->4	s->5	v->3	
"..	 ->1	
".B	a->1	å->1	
".D	e->10	
".E	n->1	u->1	
".H	i->1	
".I	 ->1	
".J	a->4	u->1	
".K	a->1	i->1	
".N	ä->1	
".O	m->1	r->1	
".R	å->1	
".V	i->1	
"; 	ö->1	
"Am	s->1	
"At	t->1	
"Bi	g->1	
"De	t->6	
"EU	-->1	
"Eq	u->1	
"Eu	r->2	
"I 	d->1	
"Ja	 ->1	,->1	g->2	
"Ku	l->4	
"Kv	i->3	
"Lo	t->1	
"Me	d->1	
"Mi	n->1	s->1	
"Ol	j->1	
"Om	 ->2	
"Po	r->1	
"Ti	b->2	
"Ty	 ->1	
"Ur	b->1	
"af	f->1	
"al	d->2	l->1	
"an	g->3	
"av	g->1	
"ba	n->1	
"co	u->1	
"de	n->3	t->1	
"di	e->1	
"dö	d->1	
"eg	e->1	
"ek	o->1	
"en	 ->3	t->1	
"eu	r->3	
"fo	r->1	
"fö	r->1	
"ge	m->1	n->1	
"he	l->1	r->1	
"in	 ->1	d->1	l->1	
"ir	r->1	
"ja	 ->1	
"ko	l->2	
"kr	o->1	
"ku	l->1	
"lä	n->1	s->2	
"me	l->1	
"na	t->1	
"ne	 ->1	
"no	r->1	
"nå	g->1	
"ob	e->1	
"or	m->1	
"ov	i->1	
"pa	r->1	
"på	p->1	
"re	f->1	s->4	
"ri	k->1	
"se	 ->1	
"sh	a->1	
"sk	a->1	
"sp	e->1	
"sv	a->1	
"ti	l->1	
"ut	v->1	å->1	
"va	l->1	r->1	
"åt	e->1	
"öp	p->1	
"öv	e->1	
'Va	d->1	
'ea	u->1	
("d	i->1	
(14	0->2	
(19	9->13	
(57	1->1	
(80	9->2	
(96	1->1	
(98	)->1	
(99	)->2	
(A5	-->36	
(Ap	p->5	
(Ar	b->1	
(B5	-->4	
(Be	n->1	
(Br	y->2	
(C5	-->7	
(CE	N->2	R->1	
(CN	S->9	
(CO	D->13	S->2	
(DA	)->2	
(DE	)->3	
(EG	,->1	
(EI	F->1	
(EL	)->3	
(EN	)->34	
(ES	)->1	
(EU	-->1	G->2	
(FI	)->1	P->1	
(FP	Ö->1	
(FR	)->18	
(FU	F->1	
(Ge	n->1	
(H-	0->21	
(Ho	w->1	
(IC	E->1	
(IF	O->1	
(IM	O->1	
(IT	)->3	
(Ih	å->1	
(In	t->1	
(KO	M->8	
(Ku	l->2	
(Li	v->2	
(NL	)->4	
(PP	E->1	
(PT	)->16	
(Pa	r->16	
(Pr	o->1	
(SE	K->1	
(SP	Ö->1	
(SY	N->1	
(Sa	m->4	
(Ta	l->8	
(Ut	s->2	
(ar	t->7	
(at	t->1	
(av	s->1	
(de	 ->1	t->1	
(ef	t->1	
(el	l->1	
(en	 ->2	
(fi	s->4	
(fo	r->1	
(fö	r->3	
(hä	l->1	
(i 	d->1	s->1	
(in	f->1	r->1	
(ko	d->2	m->1	n->1	
(kr	i->2	
(ma	i->2	
(me	r->1	
(oc	h->1	
(re	c->1	
(rå	d->1	
(se	 ->1	
(så	s->1	
(t.	e->1	
(ty	v->1	
(un	g->1	
(ÖV	P->1	
(Ös	t->4	
(åt	e->1	
) "	T->1	
) (	C->1	K->2	S->1	U->2	f->1	
) -	 ->3	
) 0	1->1	5->1	6->1	
) 1	5->1	
) 3	4->1	
) 5	1->1	2->2	
) A	t->1	
) B	o->1	
) C	5->1	
) D	e->8	
) E	f->2	
) F	P->1	r->6	å->1	ö->1	
) H	e->23	
) I	 ->5	
) J	a->15	ö->1	
) K	o->1	
) L	e->1	å->2	
) M	i->1	
) N	e->1	ä->3	
) O	m->1	
) S	e->1	
) T	a->4	h->1	i->1	
) U	n->1	
) V	a->2	e->1	i->2	
) a	d->1	v->32	
) b	ä->1	
) e	f->1	
) f	i->1	r->3	ö->5	
) h	a->3	
) i	 ->4	n->5	
) l	i->1	
) m	i->1	
) o	c->12	m->1	
) p	å->1	
) s	a->1	i->1	o->2	
) t	ä->1	
) z	o->1	
) Ä	r->1	
) ä	r->2	
)(G	e->1	
)(P	a->9	
)(T	a->1	
)) 	(->3	i->2	
))(	G->1	P->7	
)).	 ->1	.->3	F->1	J->1	
))F	r->1	
))H	e->1	
))o	c->1	
), 	b->1	d->1	m->1	o->2	r->1	s->2	t->2	v->1	ä->1	
). 	V->1	
).(	E->1	
).)	B->1	
)..	 ->2	(->2	
).D	e->5	
).F	r->2	ö->1	
).H	e->5	
).J	a->3	
).K	a->1	o->1	
).L	i->1	
).V	i->2	
)00	0->2	6->1	
)05	9->2	
)06	6->1	
):A	n->19	
); 	a->1	e->1	
)? 	H->1	
)An	d->2	g->2	s->1	
)Be	t->8	
)De	t->1	
)Fr	u->8	
)Fö	r->2	
)Ge	m->1	
)He	a->1	r->2	
)Ja	g->3	
)Ju	s->1	
)Ko	n->1	
)Nä	s->3	
)Ol	j->1	
)Re	f->1	
)Sä	k->1	
)Ta	c->1	
)Ut	t->1	
)].	)->1	H->2	
)oc	h->1	
)Åt	e->1	
, "	a->1	e->1	n->1	o->1	s->1	
, (	B->1	
, ,	 ->1	
, 1	 ->1	0->1	1->3	2->4	3->1	5->3	6->4	8->1	9->3	
, 2	 ->1	0->1	2->1	4->3	7->1	8->2	
, 3	0->1	1->1	2->2	4->1	6->1	7->2	8->1	
, 4	,->1	0->1	2->2	4->1	6->1	
, 5	0->2	6->1	
, 6	,->1	
, 7	,->2	
, 8	,->1	8->1	
, 9	,->2	5->1	
, A	l->1	m->2	n->1	r->3	s->1	
, B	N->1	e->4	r->3	u->1	
, C	o->1	u->1	
, D	a->4	i->1	u->1	
, E	C->1	D->1	E->2	G->1	f->1	r->2	u->8	v->2	
, F	i->1	r->1	ö->1	
, G	a->1	i->2	r->1	
, H	a->3	e->1	
, I	I->2	V->1	l->1	n->1	r->1	t->2	
, J	a->1	o->3	
, K	a->3	o->2	u->1	v->1	
, L	a->5	e->1	i->1	o->2	u->1	
, M	a->1	i->2	
, N	e->1	o->1	
, O	L->1	b->1	l->1	
, P	V->1	a->4	e->1	
, R	a->2	e->2	o->1	
, S	E->2	a->2	c->2	h->1	l->1	o->1	p->3	t->1	v->1	
, T	a->1	h->1	o->2	y->3	
, U	z->1	
, V	 ->1	l->1	
, W	a->1	e->1	i->1	u->1	y->1	
, Z	i->1	
, a	c->2	d->2	k->1	l->25	m->1	n->32	r->7	t->174	v->29	
, b	a->6	e->27	i->5	l->30	o->9	r->5	y->2	ä->7	å->13	ö->19	
, c	i->1	o->1	
, d	e->238	i->4	j->4	r->1	u->1	v->43	ä->66	å->28	ö->3	
, e	f->122	k->3	l->31	m->1	n->106	r->3	t->42	u->3	x->8	
, f	a->11	i->12	l->1	o->15	r->122	u->2	å->11	ö->255	
, g	a->4	e->29	i->3	j->2	l->1	o->1	r->6	u->1	y->1	ä->1	å->7	ö->9	
, h	a->94	e->153	j->2	o->4	u->18	y->3	ä->10	å->2	ö->5	
, i	 ->146	b->2	c->1	d->1	g->1	n->142	r->1	
, j	a->39	o->2	u->16	ä->10	
, k	a->45	i->1	l->2	o->90	r->13	u->8	v->3	ä->50	
, l	a->4	e->9	i->37	j->1	o->1	ä->10	å->11	ö->1	
, m	a->9	e->422	i->49	o->13	u->2	y->7	ä->9	å->27	
, n	a->13	e->6	i->4	o->2	u->6	y->5	ä->106	å->29	ö->1	
, o	a->6	b->4	c->676	f->2	l->2	m->104	p->1	r->9	s->3	t->1	
, p	a->7	e->4	l->3	o->2	r->27	u->1	å->57	
, r	a->6	e->18	i->3	o->1	ä->13	å->11	ö->5	
, s	a->38	e->12	i->7	j->4	k->51	l->4	m->2	n->7	o->388	p->11	t->22	v->3	y->1	ä->68	å->149	ö->2	
, t	.->8	a->16	e->1	i->60	j->6	o->7	r->47	u->2	v->9	y->17	ä->2	å->2	ö->1	
, u	n->26	p->14	r->3	t->166	
, v	a->67	e->10	i->248	o->4	ä->13	å->8	
, y	t->1	
, Î	l->1	
, ä	g->2	n->12	r->111	v->60	
, å	 ->1	n->1	r->1	t->29	
, ö	k->2	p->3	v->6	
,07	 ->1	
,2 	m->1	o->1	p->1	
,3 	p->1	
,4 	t->1	
,42	 ->1	
,48	7->1	
,5 	m->1	p->2	
,6 	p->1	
,7 	p->1	
,8 	m->3	t->1	
,9 	p->1	
- "	d->1	
- '	V->1	
- (	D->1	P->14	
- ,	 ->1	
- 1	9->26	
- 2	,->1	
- 3	1->1	
- 6	 ->1	
- 8	0->1	
- A	l->2	
- C	4->6	5->14	a->1	
- D	e->1	o->1	
- E	U->1	
- F	r->1	
- H	e->3	
- K	a->1	o->1	
- P	a->1	
- R	e->1	i->1	å->1	
- S	a->2	
- a	l->5	n->2	r->1	t->27	v->9	
- b	e->1	i->1	l->1	ö->1	
- c	e->1	
- d	e->51	o->1	v->2	ä->2	å->2	
- e	f->2	k->1	l->6	n->12	t->3	v->1	x->2	
- f	a->1	i->1	r->3	å->3	ö->16	
- g	e->2	ä->1	ö->2	
- h	a->10	o->1	u->3	ä->1	
- i	 ->11	d->1	n->16	
- j	a->15	u->1	
- k	a->1	n->1	o->9	r->1	
- l	i->2	y->1	å->2	
- m	a->3	e->14	i->2	o->2	å->2	
- n	a->1	y->1	ä->6	å->6	
- o	c->160	f->1	m->9	r->1	
- p	a->1	r->3	å->5	
- r	a->1	e->2	i->1	å->1	ö->1	
- s	a->5	e->3	i->1	k->3	n->2	o->26	t->3	y->2	ä->2	å->6	ö->1	
- t	a->1	e->1	i->3	r->3	v->1	ä->1	
- u	n->1	t->10	
- v	a->2	e->2	i->18	ä->1	
- Ö	s->2	
- ä	r->7	v->10	
- å	t->2	
- ö	p->1	v->4	
-(E	N->1	
-, 	S->1	a->1	d->1	f->1	i->2	m->1	s->1	t->1	u->2	ä->1	
-00	0->17	1->9	2->3	4->4	5->1	6->1	7->2	8->1	9->1	
-01	0->9	2->2	6->1	8->2	
-02	0->2	1->1	
-03	0->1	2->2	3->4	4->2	5->3	
-07	1->1	7->1	8->6	9->5	
-08	0->4	1->3	2->1	
-19	9->4	
-2 	d->1	
-2-	o->1	
-20	0->22	
-4 	p->1	
-98	/->1	
-Al	p->1	s->2	
-Ar	d->1	
-At	l->1	
-Be	h->7	
-Ca	r->1	
-Cl	a->1	
-DE	)->1	-->7	
-De	l->1	
-Ex	u->1	
-Fi	n->3	
-Fr	a->2	
-Ha	r->1	
-He	i->1	
-I)	;->1	
-II	)->1	
-Is	r->1	
-Jø	r->2	
-Ke	e->1	
-Le	 ->1	
-Lo	i->1	
-Ma	n->1	t->2	
-No	r->1	
-PM	 ->1	
-Pl	a->4	
-Ro	b->1	m->1	
-SS	:->1	
-Sh	a->1	e->5	
-Sy	r->1	
-af	f->3	
-al	b->1	
-an	a->6	p->1	
-av	t->3	v->1	
-be	l->1	n->5	s->1	
-bi	l->3	s->1	
-br	i->1	
-bu	d->1	g->1	
-da	m->1	n->1	
-de	-->3	
-di	r->3	s->2	
-do	m->22	
-ef	f->1	
-el	-->1	
-en	h->1	
-er	 ->1	
-fa	l->1	
-fo	n->1	s->1	
-fr	a->1	e->3	å->1	
-fö	r->23	
-ge	m->1	n->1	
-gr	u->20	
-ho	w->1	
-in	i->2	s->5	t->2	
-ir	l->1	
-is	r->1	
-ka	n->1	t->3	
-ko	l->1	m->3	r->20	s->1	
-kr	i->4	
-la	g->1	n->1	
-le	d->2	k->1	
-li	t->2	
-lo	b->1	
-lä	n->5	
-ma	i->1	n->1	
-me	d->6	t->1	
-na	t->1	
-ni	v->1	
-no	t->1	
-ny	t->1	
-ol	y->1	
-om	r->8	
-or	d->1	g->3	
-po	s->1	
-pr	o->27	
-ra	m->1	s->1	
-re	g->7	
-rä	t->4	
-rå	d->4	
-sh	o->1	
-si	t->1	
-sk	a->1	
-so	c->2	
-sp	r->3	
-st	a->13	i->1	o->1	r->1	ö->2	
-sy	s->1	
-sä	n->3	
-ta	l->9	
-te	s->1	x->1	
-tr	a->1	
-up	p->1	
-ut	v->1	
-va	n->1	
-vä	r->1	
-zo	n->3	
. (	E->24	F->13	P->1	
. -	(->1	
. 1	1->8	2->7	3->1	5->2	7->1	9->1	
. 2	0->1	1->2	
. 7	 ->1	)->1	
. A	l->1	v->1	
. D	e->54	ä->6	å->2	
. E	f->2	n->6	q->1	t->1	u->4	
. F	o->1	r->4	ö->3	
. G	u->1	
. H	a->1	e->3	o->1	u->1	ä->3	å->1	
. I	 ->2	n->3	
. J	a->10	
. K	o->2	ä->1	
. L	å->1	
. M	a->2	e->15	
. N	e->1	i->1	ä->1	
. O	c->4	f->1	m->1	
. P	a->1	r->1	å->1	
. R	å->1	
. S	k->2	o->2	y->1	å->2	
. T	a->1	i->1	
. U	S->1	
. V	a->3	i->12	å->2	
. W	a->1	
. a	i->1	n->1	r->2	t->12	v->3	
. b	e->1	
. d	e->8	
. e	n->2	r->1	t->3	
. f	o->1	å->1	ö->8	
. g	e->1	r->1	ö->1	
. h	o->1	u->1	
. i	 ->4	d->1	n->6	
. j	a->1	
. k	r->1	u->1	ä->1	
. m	a->2	e->3	i->3	
. n	ä->6	
. o	c->2	l->2	m->3	
. p	å->3	
. s	k->3	o->1	p->1	t->1	ä->1	
. t	r->1	
. u	n->1	t->1	
. v	a->3	i->1	
. Ä	m->1	n->2	v->1	
. Å	t->1	
. Ö	s->1	
. ä	n->1	r->1	
. ö	s->1	
." 	Ä->1	
."D	e->1	
."I	 ->1	
."J	a->1	
."M	e->1	
.(A	p->5	r->1	
.(D	A->2	E->2	
.(E	L->2	N->10	S->1	
.(F	R->6	
.(I	T->3	h->1	
.(L	i->2	
.(N	L->4	
.(P	T->1	a->5	r->1	
.(S	a->4	
.(T	a->7	
.) 	H->3	T->1	
.).	D->1	H->1	
.)A	n->3	
.)B	e->8	
.)F	r->5	ö->2	
.)G	e->1	
.)H	e->2	
.)J	u->1	
.)O	l->1	
.)R	e->1	
.)S	ä->1	
.)Å	t->1	
., 	d->1	f->1	ä->1	
.- 	(->11	D->1	F->1	H->2	
.. 	(->26	-->1	D->1	F->2	H->1	P->1	T->1	V->1	
..(	D->4	E->7	F->5	I->1	N->3	T->5	
..)	.->1	
...	(->5	)->1	.->1	F->1	H->1	L->1	
..F	r->1	
..H	e->5	
..L	å->1	
..T	a->1	
..V	i->1	
.00	.->13	
.05	 ->1	
.1 	d->1	i->3	o->2	v->1	ö->1	
.1)	 ->1	
.1.	1->1	F->1	V->1	
.12	.->1	
.14	 ->1	
.15	 ->1	
.18	 ->1	
.19	9->1	
.2 	i->5	o->1	
.2)	.->1	
.25	.->1	
.3 	E->1	b->1	i->1	
.3,	 ->1	
.30	,->1	
.3;	 ->1	
.4 	i->1	
.4.	D->1	F->1	
.50	 ->1	
.55	)->1	
.8 	i->1	
.90	 ->1	
.?A	n->1	
.Ac	c->1	
.Ah	e->1	
.Ak	t->1	
.Al	d->1	l->44	t->2	
.Am	e->1	s->1	
.An	d->4	g->1	h->1	l->1	n->4	s->4	t->2	v->1	
.Ar	a->1	b->2	t->2	
.At	t->23	
.Av	 ->26	b->1	g->1	s->15	
.Ba	k->2	r->4	
.Be	d->4	f->1	k->1	r->3	s->3	t->22	v->1	
.Bi	l->5	s->1	
.Bl	a->7	
.Bo	r->2	s->1	
.Br	e->1	i->4	y->1	
.Bu	d->1	
.By	g->1	
.Bä	s->1	
.Bå	d->5	
.CS	U->1	
.Ce	n->2	
.Co	r->1	
.Cu	n->1	
.DE	B->1	
.Da	g->5	l->1	n->1	
.De	 ->127	l->2	n->228	r->1	s->56	t->988	
.Di	r->7	s->1	
.Do	c->2	k->1	m->2	
.Dä	r->121	
.Då	 ->23	
.EG	-->3	
.EK	S->1	
.EU	 ->2	-->3	
.Ef	f->5	t->36	
.Ek	o->2	
.Em	e->8	
.En	 ->59	b->1	d->9	k->1	l->31	
.Er	 ->1	f->2	i->4	t->1	
.Et	t->43	
.Eu	r->51	
.Ev	e->1	
.Ex	c->1	e->1	p->2	
.FE	O->1	
.FP	Ö->4	
.Fa	c->3	k->4	r->1	s->1	
.Fe	l->1	m->1	
.Fi	n->4	
.Fl	e->4	o->3	
.Fo	l->2	r->2	
.Fr	a->10	e->1	i->1	u->55	å->36	
.Fy	r->1	
.Få	r->1	
.Fö	l->5	r->229	
.Ge	m->3	n->26	r->1	
.Gi	v->2	
.Go	l->1	
.Gr	a->1	e->2	u->3	
.Gä	l->1	
.Gå	 ->1	
.Gö	r->2	
.Ha	d->2	i->1	n->21	r->3	
.He	l->5	r->268	
.Hi	s->2	t->5	
.Ho	n->3	p->1	
.Hu	l->1	r->25	v->7	
.Hy	c->1	
.Hä	n->2	r->30	
.Hö	g->1	
.I 	A->1	E->4	F->1	H->1	I->3	N->1	R->1	T->2	a->11	b->4	d->69	e->16	f->14	g->2	j->1	k->4	l->6	m->7	n->4	o->4	p->3	r->11	s->26	t->1	u->2	v->18	ä->1	ö->3	
.Ib	l->3	
.Id	é->1	
.Il	l->1	
.Im	m->1	
.In	d->1	f->4	g->12	i->1	n->2	o->10	r->3	s->2	t->12	
.Ir	l->1	
.Is	r->1	
.It	a->1	
.Ja	 ->2	,->3	c->2	g->765	
.Jo	n->1	r->1	
.Ju	 ->1	s->9	
.Jä	m->2	
.Ka	f->1	n->16	r->1	t->1	
.Ki	n->3	
.Kn	a->1	
.Ko	c->1	d->1	m->104	n->19	r->2	s->4	
.Kr	a->3	
.Ku	l->7	
.Kv	a->1	i->1	
.Kä	r->6	
.La	 ->1	n->2	
.Le	d->3	
.Li	k->11	t->1	v->3	
.Ly	c->2	n->1	
.Lä	g->2	n->1	
.Lå	n->2	t->48	
.Ma	j->1	l->2	n->53	r->5	x->2	
.Me	d->46	l->3	n->192	r->3	
.Mi	l->1	n->45	t->2	
.Mo	r->1	t->8	
.My	l->1	n->3	
.Mä	n->4	r->1	
.Må	h->1	l->2	n->10	
.Mö	j->2	
.Na	t->17	
.Ne	j->1	
.Ni	 ->35	e->1	v->1	
.No	r->1	
.Nu	 ->26	m->1	v->1	
.Ny	a->1	l->1	
.Nä	r->64	s->1	
.Nå	g->4	j->1	
.Nö	d->1	
.OK	,->1	
.OL	A->2	
.OM	R->2	
.Oa	v->2	
.Ob	e->2	
.Oc	h->60	k->2	
.Of	f->2	t->1	
.Om	 ->93	r->15	
.On	ö->1	
.Or	d->11	k->2	o->2	s->2	
.Oz	 ->1	
.PP	E->2	
.Pa	r->22	
.Pe	r->4	
.Pl	a->3	ä->1	
.Po	r->2	
.Pr	e->6	o->18	
.Pu	n->2	
.På	 ->42	
.Ra	p->3	s->1	
.Re	a->1	d->3	f->6	g->5	n->2	s->7	t->1	v->2	
.Ri	k->4	s->1	
.Ro	p->1	t->2	
.Ru	m->1	
.Rä	k->1	t->2	
.Rå	d->16	
.Sa	m->24	n->5	v->2	
.Sc	h->3	
.Se	d->15	t->1	
.Si	s->2	t->3	
.Sj	u->1	ä->2	
.Sk	a->4	o->1	u->4	y->1	
.Sl	u->38	
.Sm	å->2	
.Sn	a->2	
.So	c->3	m->45	
.St	a->9	o->4	r->3	ä->1	å->1	ö->10	
.Su	b->2	
.Sv	e->1	
.Sy	f->6	r->1	
.Sä	g->1	k->1	r->2	
.Så	 ->32	d->2	l->4	n->1	s->2	v->1	
.TV	-->1	
.Ta	 ->1	c->28	d->1	l->1	n->3	
.Te	r->1	
.Th	e->2	y->1	
.Ti	d->1	l->37	t->1	
.To	n->1	p->2	r->2	
.Tr	a->2	e->1	o->18	ä->1	
.Tu	s->1	
.Tv	ä->3	å->2	
.Ty	 ->7	d->1	v->9	
.Tä	n->1	
.Un	d->30	g->3	i->5	
.Up	p->6	
.Ur	 ->4	
.Ut	a->3	b->2	d->1	e->1	f->3	g->1	i->1	m->2	n->1	s->2	v->2	
.Va	d->59	l->3	n->2	r->25	
.Ve	m->4	r->1	t->2	
.Vi	 ->503	a->1	d->19	k->1	l->16	n->1	s->13	t->3	
.Vo	n->1	
.Vä	r->1	s->2	
.Vå	r->26	
.Wo	r->1	
.Yt	t->3	
.a.	 ->28	
.d.	 ->2	,->1	
.ex	.->20	
.g.	a->1	
.k.	 ->4	
.ko	m->1	
.m.	 ->6	,->1	O->1	
.o.	m->7	
.Än	 ->3	d->19	n->1	t->1	
.Är	 ->15	a->3	
.Äv	e->31	
.Å 	E->1	a->10	e->2	
.År	 ->5	e->1	
.Åt	a->1	e->2	g->2	
.ÖV	P->1	
.Ög	o->2	
.Ök	a->1	
.Ös	t->2	
.Öv	e->2	r->1	
/00	 ->1	)->2	1->2	8->1	9->1	
/01	0->2	6->2	9->2	
/02	2->1	4->2	
/03	1->1	5->1	7->4	
/08	0->2	2->2	
/1/	1->2	
/19	9->41	
/20	0->26	
/21	2->2	
/3 	a->1	
/35	/->4	
/40	9->1	
/43	.->1	
/55	/->2	
/59	1->2	
/60	/->1	
/71	 ->1	/->1	
/72	8->1	
/75	 ->1	
/92	 ->1	
/95	.->1	
/98	 ->1	-->1	
/99	 ->5	)->22	.->1	
/EG	 ->5	,->3	
/EK	S->2	
/Eu	r->1	
/NG	L->2	
/No	r->2	
/Oi	l->1	
/de	n->1	
/el	l->1	
/ha	l->1	
/in	t->1	
/ri	k->1	
/sa	m->1	
/år	)->1	,->1	
0 -	 ->6	
0 0	0->11	
0 E	n->1	
0 a	n->1	r->3	t->1	
0 b	a->1	i->1	
0 d	e->1	o->2	ö->1	
0 e	l->2	n->1	u->1	
0 f	r->5	å->2	ö->1	
0 g	u->1	å->1	
0 h	a->3	e->1	
0 i	 ->7	n->3	
0 j	a->1	u->2	
0 k	a->1	i->4	m->4	
0 l	ä->1	
0 m	e->2	i->19	o->1	
0 n	y->1	ä->1	
0 o	c->7	l->1	
0 p	r->37	å->1	
0 r	i->1	
0 s	k->2	o->2	t->1	
0 t	i->1	o->10	
0 u	t->2	
0 v	a->1	
0 º	 ->1	
0 ä	n->7	r->5	
0 å	r->10	t->1	
0" 	s->1	t->2	
0".	D->1	V->1	
0(C	N->2	O->3	
0) 	a->20	f->2	o->1	
0).	F->1	J->1	
0):	A->1	
0, 	1->1	2->1	3->1	4->1	d->1	f->1	i->1	m->2	o->1	s->2	ä->1	
0- 	o->1	
0-2	0->17	
0-b	u->1	
0-p	r->4	
0-t	a->9	
0.(	S->2	
0.)	A->1	O->1	
0.2	5->1	
0.4	.->1	
0.D	e->6	
0.F	a->1	r->1	ö->2	
0.J	a->2	
0.K	o->1	
0.M	a->1	e->1	
0.O	M->1	
0.S	a->1	t->2	
0.T	i->1	r->1	
0.V	i->1	
0/1	9->4	
0/2	0->3	
0/9	2->1	9->4	
00 	-->4	0->6	E->1	a->4	b->2	d->1	f->3	h->4	i->2	k->8	l->1	m->6	n->1	o->5	p->2	s->4	t->11	u->1	v->1	ä->8	å->1	
00"	 ->3	.->2	
00)	 ->23	.->2	:->1	
00,	 ->7	
00-	2->17	b->1	p->4	t->4	
00.	(->2	)->2	D->5	F->4	J->2	M->2	O->1	S->3	T->2	V->1	
000	 ->48	"->5	)->24	,->7	-->26	.->11	1->1	2->1	3->6	4->2	6->4	7->3	9->2	N->1	
001	 ->1	,->1	/->1	0->2	1->2	2->3	3->1	8->3	
002	 ->2	)->2	,->2	.->5	/->1	0->1	2->2	
003	 ->2	/->4	?->1	
004	 ->1	.->2	/->2	0->1	1->1	5->2	
005	0->1	
006	 ->11	,->5	.->9	/->4	6->1	9->1	
007	,->1	/->3	3->1	8->1	
008	 ->2	3->1	7->1	
009	/->2	0->1	5->1	
00N	ä->1	
01 	ä->1	
01,	 ->1	
01/	2->1	9->1	
010	 ->1	/->2	4->2	5->2	6->3	7->2	8->2	
011	/->2	3->1	
012	 ->1	(->1	/->2	0->1	2->1	
013	(->1	
016	7->1	9->2	
018	/->3	0->2	
019	4->2	
02 	(->1	f->1	
02)	 ->2	
02,	 ->2	
02.	 ->1	H->1	M->1	P->1	V->1	
02/	2->1	
020	/->1	8->2	
021	2->1	
022	/->2	8->1	
024	0->2	
03 	-->2	
03(	C->1	
03/	2->4	
030	5->1	
031	8->1	
032	7->2	
033	3->2	4->2	
034	1->2	
035	0->1	1->1	2->2	
037	0->2	1->2	
03?	H->1	
04 	i->1	
04.	D->1	K->1	
04/	1->3	2->1	
040	/->1	
041	/->1	
045	/->2	
05 	i->1	o->1	t->1	
05(	C->1	
05/	1->3	9->1	
050	/->1	
055	0->1	
059	8->2	
06 	[->1	f->2	g->1	k->1	l->1	o->1	s->1	t->2	å->1	
06(	C->2	
06,	 ->5	
06.	D->2	E->1	F->1	H->1	J->2	M->1	T->1	
06/	0->2	1->1	2->2	
065	2->1	
066	 ->1	2->1	
069	/->1	
07 	m->1	
07,	 ->1	
07/	1->2	2->3	9->1	
071	5->1	
073	/->1	
077	8->1	
078	/->1	0->1	1->1	2->1	5->1	6->1	8->1	
079	1->1	3->1	5->1	6->1	8->1	
08 	t->2	
08/	1->4	9->1	
080	1->1	3->1	5->2	7->1	8->1	
081	3->1	7->1	9->1	
082	5->2	9->1	
083	 ->1	
087	/->1	
09 	o->1	
09/	2->2	
090	(->1	
094	/->2	
095	/->3	
0Nä	s->1	
1 0	0->2	
1 4	0->1	
1 a	n->1	
1 d	å->1	
1 e	f->1	
1 f	r->3	
1 g	e->1	
1 i	 ->5	
1 j	a->9	u->2	
1 m	a->4	e->1	i->1	
1 o	c->19	m->1	
1 p	r->7	
1 r	i->1	
1 s	e->1	t->2	
1 u	r->2	t->1	
1 v	i->1	
1 ä	n->1	r->1	
1 å	r->1	
1 ö	v->1	
1(C	O->2	
1) 	e->1	
1, 	1->2	2->1	4->1	a->1	f->1	m->1	o->1	s->1	
1,2	 ->2	
1,3	 ->1	
1,4	 ->1	
1-2	 ->1	
1-o	m->4	
1-r	e->5	
1-s	t->2	
1.0	0->4	
1.1	 ->4	.->2	
1.3	 ->3	,->1	;->1	
1.5	5->1	
1.A	l->1	
1.E	x->1	
1.F	ö->1	
1.J	a->1	
1.K	u->1	
1.V	i->1	
1/1	9->5	
1/2	0->3	
1/3	 ->1	
1/9	9->4	
1/E	G->1	K->2	
10 	0->2	e->2	f->1	i->1	j->1	k->1	m->2	p->4	r->1	s->1	ä->2	å->1	
10,	 ->1	
10.	K->1	
10/	2->2	
100	 ->9	
104	/->2	
105	 ->2	/->2	
106	(->2	/->1	
107	/->2	
108	/->2	
11 	i->1	j->2	m->1	o->1	s->1	
11,	 ->3	3->1	
11.	0->3	A->1	E->1	K->1	
11/	2->2	
110	 ->1	
113	 ->1	
115	 ->1	
12 	e->1	f->1	i->1	j->1	m->2	o->1	p->1	s->1	
12(	C->1	
12,	 ->4	
12.	0->7	
12/	1->1	2->2	9->3	
120	 ->1	/->1	
122	/->1	
123	 ->1	(->1	
124	4->3	
125	 ->1	
126	0->1	
127	(->1	
13 	(->1	-->1	0->1	A->1	f->1	i->2	j->1	n->1	o->1	p->2	s->1	ä->1	
13(	C->1	
13,	 ->2	
13.	0->1	F->1	
13/	1->1	9->1	
130	 ->1	
133	.->1	
138	.->1	
14 	e->1	f->5	l->1	m->5	o->1	s->1	t->1	
14,	 ->1	
14/	1->1	
140	 ->1	9->2	
143	 ->1	
15 	a->1	m->3	o->3	p->3	r->1	s->2	å->1	
15,	 ->2	
15.	0->2	
15/	9->1	
150	 ->2	
158	 ->2	)->1	.->1	
16 	0->1	o->3	p->2	r->1	
16)	 ->1	
16,	 ->1	
164	 ->1	
166	 ->1	
167	 ->3	/->1	
169	(->2	
17 	d->2	m->1	o->2	s->1	
17,	 ->2	
17.	3->1	S->1	
17/	9->1	
170	 ->1	
174	 ->1	
176	2->2	
18 	d->1	h->1	i->1	m->3	n->3	
18(	S->1	
18,	 ->1	
18/	2->2	9->1	
180	 ->1	/->2	
19 	-->1	d->1	m->1	p->1	s->1	ä->1	
19.	5->1	
19/	9->1	
191	7->1	
192	3->1	
193	 ->1	0->1	
194	(->2	.->1	5->1	8->1	
195	 ->1	7->2	
196	7->6	9->1	
197	6->1	7->1	
198	2->2	6->3	9->1	
199	0->2	1->3	2->4	3->8	4->6	5->9	6->18	7->42	8->33	9->126	
1:a	 ->1	
2 (	K->1	
2 -	 ->4	
2 0	0->1	
2 4	0->1	
2 a	v->1	
2 b	l->2	
2 d	a->1	e->1	
2 e	l->1	n->1	u->1	
2 f	a->1	r->2	
2 h	a->1	
2 i	 ->12	n->2	
2 j	a->1	
2 m	i->5	å->1	
2 o	c->9	
2 p	r->4	u->1	
2 r	i->1	
2 s	k->1	o->2	t->1	
2 u	n->1	p->1	
2 å	r->1	
2(C	N->1	O->1	
2) 	-->2	f->1	
2).	K->1	
2, 	1->3	2->2	3->2	d->2	e->2	f->1	i->2	k->1	l->1	s->3	t->2	v->2	
2,4	8->1	
2,5	 ->1	
2,6	 ->1	
2,8	 ->1	
2-o	m->3	
2-s	t->1	
2. 	J->1	
2.0	0->7	
2.1	 ->1	
2.2	 ->1	
2.D	e->1	
2.H	e->1	
2.I	 ->1	s->1	
2.J	a->1	
2.M	a->1	e->1	i->1	
2.P	å->1	
2.V	i->1	
2.Ä	v->1	
2/1	9->3	
2/2	0->5	
2/4	3->1	
2/9	9->4	
20 	-->1	0->1	e->1	f->1	g->1	m->3	n->1	p->3	º->1	ä->1	å->5	
20,	 ->1	
20.	2->1	
20/	1->1	9->1	
200	 ->5	0->97	1->2	2->11	3->1	4->3	6->25	7->1	
201	0->1	2->1	
208	/->2	
21 	j->2	o->2	s->1	ä->1	å->1	
21.	0->1	5->1	
212	/->1	3->1	7->1	
21:	a->1	
22 	-->1	a->1	r->1	
22,	 ->3	5->1	
22.	Ä->1	
22/	1->1	2->2	
226	 ->1	
228	(->1	
23 	d->1	i->1	p->1	
23(	C->1	
23,	 ->1	7->1	
24 	n->2	o->2	p->1	
240	(->2	
244	 ->1	.->2	
245	 ->1	
248	,->1	
25 	g->1	m->3	o->1	p->7	t->1	
25(	C->2	
25.	)->1	D->1	
250	 ->1	
255	 ->4	
26 	"->1	i->2	m->1	n->1	o->1	p->1	
260	/->1	
262	 ->1	
27 	d->1	f->1	l->1	o->1	p->2	
27(	C->1	
27,	 ->1	
27/	1->2	
28 	f->1	j->1	n->1	p->1	
28(	C->1	
28,	 ->2	
28/	E->1	
280	 ->4	.->1	
28:	e->1	
29 	d->1	f->1	l->1	m->1	
29,	 ->1	
29/	9->1	
299	.->2	
3 (	C->1	E->1	
3 -	 ->3	
3 0	0->5	
3 A	m->1	
3 E	G->1	
3 a	v->2	
3 b	l->1	
3 d	e->1	
3 f	e->2	r->1	ö->1	
3 h	a->1	ö->1	
3 i	 ->3	n->2	
3 j	a->2	
3 m	a->1	
3 n	y->1	
3 o	c->4	k->2	m->1	
3 p	e->2	r->6	u->1	
3 s	a->1	
3 u	t->1	
3 ä	r->1	
3(C	N->2	O->1	
3, 	1->1	2->2	7->1	e->1	n->1	
3,7	 ->1	
3,8	 ->2	
3,9	 ->1	
3-1	9->2	
3-4	 ->1	
3-l	i->2	
3.0	5->1	
3.1	)->1	
3.2	 ->1	
3.8	 ->1	
3.F	r->1	ö->1	
3.I	 ->1	
3.O	m->1	
3.T	y->1	
3/1	9->4	
3/2	0->4	
3/7	5->1	
3/9	9->2	
30 	d->1	f->1	i->2	j->1	m->2	o->1	p->3	
30,	 ->2	
30-	t->1	
300	 ->1	
305	/->1	
31 	f->1	j->1	m->2	o->2	
314	 ->1	
318	(->1	
32 	m->1	
32,	 ->3	
32.	J->1	
327	/->2	
33 	0->2	a->1	f->2	i->1	o->1	
33.	2->1	
33/	1->2	
332	,->1	
333	/->2	
334	/->2	
34 	i->1	s->1	t->1	å->1	
34,	 ->1	
34.	1->1	
34/	1->2	
341	/->2	
344	 ->1	
35 	f->1	m->5	
35.	S->1	
35/	E->4	
350	 ->1	/->1	
351	/->1	
352	(->1	/->1	
36 	f->1	
36,	 ->1	
367	 ->1	
37 	f->1	i->1	p->1	
37,	 ->2	
37.	2->1	
37/	6->1	
370	 ->1	(->2	
371	(->2	
38 	f->2	o->2	
38,	 ->1	
38.	4->1	
38:	 ->1	
39 	f->1	i->1	p->1	
39,	 ->1	
3: 	f->1	
3; 	d->1	
3?F	r->1	
3?H	e->1	
4 -	 ->1	
4 0	0->1	
4 c	 ->1	
4 e	n->1	t->1	u->1	
4 f	e->5	r->1	
4 h	a->1	
4 i	 ->6	n->2	
4 j	u->2	
4 l	e->1	i->1	
4 m	e->5	
4 n	y->2	ä->1	
4 o	c->8	k->1	
4 p	r->5	
4 r	ö->1	
4 s	e->1	k->1	
4 t	i->2	r->1	u->1	
4 å	r->1	
4(C	O->2	
4, 	1->2	3->1	6->1	e->1	f->1	k->1	o->1	
4-0	0->1	2->1	3->3	7->1	
4-1	9->1	
4.1	.->1	
4.2	)->1	
4.D	e->3	
4.F	ö->1	
4.I	 ->3	
4.J	a->2	
4.K	o->1	
4/1	9->8	
4/2	0->1	
4/5	5->2	
4/7	2->1	
40 	f->1	j->1	m->2	p->6	å->3	
40(	C->2	
40,	 ->1	
40/	9->1	
400	 ->6	
409	 ->1	4->2	
41 	f->1	p->1	r->1	u->1	
41/	1->2	9->1	
410	 ->1	
42 	f->1	i->1	m->1	o->2	
43 	h->1	o->1	
43.	F->1	T->1	
44 	-->1	f->1	o->3	
44.	I->1	J->1	
45 	a->1	c->1	f->1	g->1	o->1	
45,	 ->1	
45.	 ->1	"->1	F->1	H->1	V->1	
45/	0->1	2->1	
46 	o->2	
462	 ->1	
47 	g->1	
48 	g->1	i->3	ä->1	
48,	 ->1	
48.	D->1	
487	 ->1	
5 (	e->1	
5 -	 ->1	
5 0	0->5	
5 a	v->2	
5 c	e->1	
5 f	r->3	
5 g	r->1	ä->2	
5 h	a->1	
5 i	 ->5	n->1	
5 k	o->1	
5 m	a->2	e->1	i->17	o->1	
5 o	c->4	k->1	l->2	m->3	
5 p	r->14	
5 r	i->1	ä->1	
5 s	e->1	l->1	t->1	
5 t	i->4	
5 v	i->1	
5 å	r->3	
5(C	N->3	
5)U	t->1	
5, 	1->2	d->2	n->1	o->2	u->1	
5,5	 ->1	
5,8	 ->1	
5-0	0->37	1->14	2->2	3->9	
5-1	9->1	
5. 	D->1	
5."	I->1	
5.)	J->1	
5.0	0->2	
5.4	 ->1	
5.D	e->1	
5.E	m->1	
5.F	r->2	
5.H	e->1	
5.S	å->1	
5.V	i->1	
5/0	0->1	
5/1	/->2	9->4	
5/2	0->1	
5/3	5->1	
5/9	5->1	8->1	9->3	
5/E	G->6	
50 	-->1	0->1	g->1	i->1	m->4	o->2	p->3	
50,	 ->1	
50-	 ->1	t->2	
50/	1->1	2->1	
500	 ->1	
51/	1->1	
519	 ->1	
52 	-->1	i->1	
52(	C->1	
52/	1->1	
520	 ->2	
522	 ->1	
53 	p->1	
540	 ->1	
55 	i->4	m->1	p->1	
55)	U->1	
55/	E->2	
550	 ->1	
56 	p->1	
56,	 ->1	
57 	(->1	
57,	5->1	
57.	E->1	
571	3->1	
58 	-->1	i->1	
58)	.->1	
58.	1->1	
591	/->2	
598	 ->2	
5b 	k->1	
5b-	o->1	
5b.	D->1	
6 "	p->1	
6 -	 ->2	
6 0	0->1	
6 [	K->1	
6 d	e->1	
6 e	f->1	l->1	m->1	
6 f	r->2	ö->2	
6 g	ä->1	
6 h	a->2	
6 i	 ->10	n->1	
6 k	o->1	
6 l	i->1	å->1	
6 m	e->1	i->1	
6 n	o->1	
6 o	c->15	m->1	
6 p	e->1	r->6	
6 r	a->1	
6 s	å->1	
6 t	a->1	o->1	
6 v	a->1	i->1	
6 ä	r->1	
6 å	r->2	t->1	
6(C	O->2	
6) 	s->1	
6, 	2->1	3->1	7->1	f->1	h->1	m->1	n->1	s->3	t->1	v->1	
6,0	7->1	
6.D	e->3	
6.E	n->2	
6.F	r->1	
6.H	e->1	
6.J	a->3	
6.M	a->1	e->1	
6.O	c->1	
6.S	å->1	
6.T	a->1	
6.Å	r->1	
6/0	0->2	
6/1	9->1	
6/2	0->2	
6/3	5->3	
6/7	1->2	
6/9	9->2	
60 	0->1	f->1	
60-	t->1	
60/	9->2	
600	 ->1	
614	/->1	
62 	-->1	e->1	i->1	u->2	
62.	M->1	
64 	r->1	
652	 ->1	
66 	-->1	e->1	
662	 ->1	
67 	0->1	h->1	i->2	m->4	o->2	
67,	 ->1	
67/	1->1	
68 	a->1	
685	/->1	
69 	o->1	
69(	C->2	
69/	1->1	
7 (	a->1	m->1	
7 -	 ->3	
7 0	0->1	
7 d	e->4	ä->1	
7 f	a->1	r->1	ö->2	
7 g	r->1	ä->1	
7 h	a->2	ä->1	
7 i	 ->12	
7 l	e->1	y->1	ä->1	
7 m	e->1	i->7	
7 n	ä->1	
7 o	c->11	k->1	m->1	
7 p	r->5	å->2	
7 s	å->1	
7 t	r->2	
7 u	p->1	
7 ä	r->1	
7 å	r->1	
7(C	O->1	
7) 	0->1	
7).	.->1	
7, 	1->1	3->1	4->2	8->1	9->1	d->1	m->1	o->3	r->1	s->2	v->1	
7,2	 ->1	
7,4	2->1	
7,5	 ->1	
7.-	 ->1	
7..	 ->1	
7.1	 ->1	
7.2	 ->2	
7.3	0->1	
7.B	e->1	
7.D	e->2	
7.E	u->1	
7.F	r->1	
7.I	 ->1	
7.M	a->1	
7.N	u->1	
7.S	e->1	l->1	
7.V	i->2	
7/0	1->2	3->5	
7/1	9->6	
7/2	0->3	
7/6	0->1	
7/9	9->3	
70 	a->1	m->2	p->1	
70(	C->2	
700	 ->4	
71 	a->1	
71(	C->2	
71/	E->1	
713	/->1	
715	/->1	
728	/->1	
73,	9->1	
73/	1->1	
74 	t->1	
75 	-->1	m->2	o->1	
76 	e->1	p->1	
762	 ->1	.->1	
77 	-->1	m->1	
778	/->1	
78/	1->1	9->1	
780	/->1	
781	/->1	
782	/->1	
785	/->1	
786	/->1	
788	/->1	
79/	4->1	
791	/->1	
793	/->1	
795	/->1	
796	/->1	
798	/->1	
7?D	e->1	
7Nä	s->1	
8 -	 ->4	
8 4	6->1	
8 a	t->1	
8 b	e->1	
8 d	e->1	
8 f	r->3	ö->1	
8 g	o->1	ä->1	
8 h	a->1	ä->1	
8 i	 ->6	n->1	
8 j	u->1	
8 k	o->1	
8 m	i->6	å->1	
8 n	o->3	y->1	
8 o	c->12	
8 p	r->1	
8 r	e->2	
8 s	k->1	
8 t	i->2	o->2	
8 u	n->1	t->2	
8 v	a->2	
8 ä	n->1	r->4	
8(C	N->1	
8(S	Y->1	
8) 	5->3	
8).	D->1	
8)0	6->1	
8, 	2->2	3->2	4->1	9->1	S->2	d->1	s->1	
8-2	0->2	
8-9	8->1	
8. 	D->1	
8.1	 ->1	
8.4	.->1	
8.D	e->1	
8.P	r->1	
8.S	t->1	
8/0	1->4	3->1	
8/1	9->5	
8/2	0->2	
8/5	9->2	
8/9	8->1	9->4	
8/E	G->1	
80 	e->1	i->4	m->1	p->11	ä->1	å->1	
80.	4->1	
80/	1->2	9->1	
801	/->1	
803	(->1	
805	(->1	/->1	
807	/->1	
808	/->1	
809	5->2	
81 	o->5	p->1	
81.	1->5	3->5	
81/	9->1	
813	/->1	
817	/->1	
819	/->1	
82 	h->1	i->1	
82)	 ->1	
82,	 ->5	
82.	I->2	
82/	9->1	
825	(->2	
829	/->1	
83 	(->1	p->1	
85 	o->2	p->1	t->1	
85/	9->2	
86 	h->1	i->2	o->1	p->1	
86.	Å->1	
86/	9->1	
87 	m->1	
87,	 ->1	
87.	1->1	2->1	
87/	1->1	
88 	i->1	o->1	ä->1	
88/	5->2	9->1	
89 	i->1	t->1	
89,	 ->1	
8: 	f->1	
8:e	 ->1	
9 (	H->1	
9 -	 ->28	
9 a	n->3	v->1	
9 b	e->1	
9 d	e->2	ä->1	ö->1	
9 e	r->1	
9 f	a->1	e->1	r->5	
9 g	o->1	
9 h	a->5	
9 i	 ->5	n->2	
9 j	ä->1	
9 k	a->1	o->2	u->1	
9 l	ä->1	
9 m	a->1	i->4	
9 n	ä->1	
9 o	c->7	m->1	
9 p	r->4	
9 r	a->1	
9 s	k->1	o->1	
9 t	i->2	
9 u	p->2	t->1	
9 v	a->2	i->1	
9 ä	r->1	v->1	
9 å	r->1	
9 ö	v->1	
9".	B->1	
9(C	O->2	
9) 	0->2	1->1	3->1	a->12	f->2	o->1	
9).	K->1	
9)0	0->3	5->2	
9):	A->18	
9)A	n->2	
9, 	1->1	3->1	4->1	a->2	b->1	d->1	f->1	h->1	n->1	o->2	
9-2	0->2	
9. 	V->1	
9..	(->1	
9.1	 ->1	
9.2	 ->2	
9.5	0->1	
9.D	e->3	
9.E	n->1	u->1	
9.F	r->1	ö->2	
9.J	a->2	
9.K	o->1	
9.U	n->1	
9.V	i->1	
9/0	0->4	2->3	8->4	
9/1	9->1	
9/2	0->2	1->2	
9/4	0->1	
9/9	9->2	
90 	d->2	p->4	u->1	
90(	C->1	
90-	t->1	
90.	D->1	
91 	e->1	g->1	o->1	p->1	
91/	9->1	E->2	
917	 ->1	
92 	o->1	s->2	å->1	
92,	 ->1	
92/	4->1	
923	,->1	
93 	h->1	o->2	p->1	u->1	
93,	 ->1	
93-	1->2	
93.	O->1	
93/	7->1	9->1	
930	-->1	
93?	F->1	
94 	e->1	h->1	n->1	o->2	p->2	
94(	C->2	
94,	 ->2	
94-	1->1	
94.	D->1	
94/	1->2	5->2	7->1	
945	.->1	
948	.->1	
95 	(->1	h->1	i->1	k->1	m->3	r->1	s->1	t->1	å->1	
95,	 ->2	
95-	1->1	
95.	F->1	
95/	1->3	3->1	9->1	
957	 ->1	.->1	
96 	-->1	e->1	h->1	i->1	l->1	o->1	v->2	ä->1	å->2	
96,	 ->2	
96.	D->1	E->1	J->1	M->1	O->1	
96/	3->3	7->2	9->1	
961	4->1	
967	 ->5	,->1	
969	 ->1	
97 	(->1	-->1	d->1	f->1	h->2	i->1	l->1	o->6	p->1	t->2	u->1	ä->1	å->1	
97)	 ->1	
97,	 ->2	
97.	-->1	.->1	B->1	D->2	I->1	M->1	N->1	S->1	V->2	
97/	0->7	9->1	
976	 ->1	
977	 ->1	
97?	D->1	
97N	ä->1	
98 	-->3	g->1	h->1	k->1	m->1	o->6	r->1	s->1	u->3	v->2	ä->2	
98)	 ->3	0->1	
98,	 ->3	
98-	2->2	9->1	
98.	 ->1	P->1	S->1	
98/	0->5	9->1	
982	,->1	.->1	
986	 ->2	.->1	
989	,->1	
99 	(->1	-->27	a->4	b->1	d->1	e->1	f->2	g->1	h->5	i->4	j->1	k->4	n->1	o->6	p->1	r->1	s->1	t->1	u->3	v->3	ä->1	å->1	ö->1	
99"	.->1	
99)	 ->19	.->1	0->5	:->18	A->2	
99,	 ->7	
99-	2->2	
99.	 ->1	.->1	2->2	D->3	E->2	F->3	J->2	K->1	U->1	V->1	
99/	0->11	2->2	
990	 ->1	.->1	
991	 ->3	
992	 ->3	,->1	
993	 ->3	,->1	-->2	.->1	?->1	
994	 ->4	,->1	-->1	
995	 ->6	,->2	-->1	
996	 ->11	,->2	.->5	
997	 ->20	)->1	,->2	.->10	/->7	?->1	N->1	
998	 ->18	)->3	,->3	-->2	.->3	/->4	
999	 ->67	"->1	)->21	,->7	-->2	.->14	/->13	:->1	
99:	 ->1	
9: 	"->1	
: "	A->1	D->4	J->1	M->1	O->1	a->1	d->1	h->1	i->1	j->1	v->1	
: A	n->2	r->2	s->1	t->1	
: D	e->9	
: E	f->1	r->1	u->1	
: F	i->2	l->1	r->3	ö->5	
: G	e->2	r->1	
: H	a->2	o->1	
: I	 ->3	n->1	
: J	a->7	o->1	
: K	o->6	ä->2	
: M	a->1	
: N	a->1	y->1	ä->3	
: O	m->1	s->1	
: P	a->1	o->1	å->1	
: R	e->1	
: S	t->2	
: T	u->1	å->1	
: U	n->2	t->2	
: V	a->4	e->3	i->7	
: a	n->4	t->8	
: b	a->1	e->1	
: d	e->25	i->1	u->1	ä->1	
: e	n->8	t->2	
: f	o->2	r->2	ö->12	
: g	e->2	ö->1	
: h	a->2	u->4	ö->1	
: i	 ->3	n->3	
: j	a->5	
: k	a->1	o->3	
: m	a->1	e->2	i->1	
: n	u->1	ä->2	
: o	m->4	p->1	
: p	a->1	r->1	
: r	ä->1	
: s	k->1	y->1	
: t	a->1	i->1	o->1	
: u	n->1	p->1	t->4	
: v	a->5	e->3	i->12	å->2	
: Ä	r->1	v->1	
: Å	t->2	
: Ö	p->1	
: å	 ->1	
: ö	n->1	
:An	g->19	
:De	n->1	t->1	
:Fö	r->2	
:a 	å->1	
:e 	r->2	å->1	
:s 	(->1	B->1	E->1	a->4	b->8	d->3	e->3	f->4	g->3	h->2	i->6	k->2	l->3	m->5	n->2	o->6	p->4	r->2	s->8	t->2	u->3	v->1	
:s.	L->1	
; D	a->1	
; J	a->1	
; a	l->1	n->2	r->1	t->3	v->1	
; b	)->1	
; d	e->31	ä->1	å->1	
; e	n->7	
; f	i->1	o->1	r->1	ö->7	
; h	ä->1	
; i	 ->3	n->4	
; j	a->4	
; k	o->1	
; l	o->1	
; m	a->1	e->2	i->2	
; o	c->5	
; p	u->3	
; s	a->1	k->1	l->1	
; u	n->1	
; v	i->6	
; ä	n->1	
; å	 ->1	
; ö	v->1	
? 2	1->1	
? D	e->2	
? H	a->2	
? I	n->1	
? M	e->1	
? O	c->1	
? R	å->1	
?"J	a->1	
?, 	r->2	
?- 	(->3	
?. 	(->9	
?.(	E->2	
?.H	e->2	
?An	s->4	
?At	t->2	
?Av	 ->1	s->1	
?Bo	r->1	
?Da	g->1	
?De	 ->3	n->8	s->1	t->19	
?Dä	r->3	
?Ef	t->1	
?El	l->1	
?En	d->1	l->1	
?Et	t->3	
?Eu	r->2	
?Fi	n->1	
?Fo	l->1	
?Fr	u->6	å->3	
?Fö	r->8	
?Ha	r->4	
?He	m->1	r->15	
?Hu	r->10	
?Hä	r->2	
?I 	F->1	d->2	e->1	f->1	m->1	s->1	v->1	
?In	i->1	t->1	
?Ja	,->2	g->21	
?Jo	 ->1	,->3	
?Ka	n->5	
?Ko	l->1	m->6	
?Kä	r->1	
?Ma	n->1	
?Me	n->3	
?Na	t->1	
?Ne	j->6	
?Ni	 ->3	
?Nä	r->3	s->1	
?Oc	h->3	
?Ol	i->1	
?Om	 ->2	
?Pa	r->1	
?Pr	o->1	
?På	 ->2	
?RI	N->1	
?Re	g->1	
?Se	d->1	r->1	
?Sk	u->3	
?So	m->2	
?Sv	a->1	
?Ta	c->1	
?Ti	l->1	
?Ty	c->1	
?Tä	n->1	
?Ut	g->1	
?Va	d->7	
?Ve	m->2	t->1	
?Vi	 ->11	l->13	s->2	
?Är	 ->11	
?Äv	e->2	
A -	 ->1	
A O	C->1	
A a	t->1	
A e	l->1	
A h	a->3	
A p	å->1	
A v	a->1	
A) 	D->1	V->1	
A, 	K->1	e->1	s->1	
A-i	n->1	
A-s	t->1	
A. 	G->1	
A.J	a->1	
A.V	i->1	
A5-	0->36	
A:s	.->1	
ABB	 ->1	-->2	
ABC	 ->1	
ADR	)->1	
AF 	g->1	i->2	k->2	s->1	
AF,	 ->8	
AF.	A->1	F->1	H->1	M->1	
AF:	s->2	
AKT	U->1	
AND	E->1	
ARP	O->1	
AS 	(->1	
ASP	 ->1	
ATT	 ->1	
Acc	e->1	
Act	.->1	
Ada	n->1	
Ade	n->1	
Ado	l->2	
Adr	i->1	
Afr	i->4	
Agr	i->1	
Agu	s->1	
Ahe	r->8	
Aid	s->1	
Akk	u->2	ö->1	
Akt	i->1	
Ala	v->2	
Alb	a->2	e->1	r->1	
Ald	r->1	
Ale	x->2	
Alg	e->1	
Ali	c->1	
All	a->25	d->1	m->4	t->21	
Alp	e->2	
Als	a->3	t->3	
Alt	e->18	
Ame	r->2	
Amo	c->1	k->5	s->1	
Ams	t->39	
And	r->7	
Ang	e->1	å->22	
Anh	å->1	
Ank	a->1	
Anl	e->1	ä->1	
Anm	ä->1	
Ann	a->5	
Ans	e->4	l->1	v->4	
Ant	a->2	ó->1	
Anv	e->1	ä->1	
Apa	r->1	
App	l->5	
Ara	b->2	f->1	
Arb	e->4	
Ard	e->1	
Ari	 ->1	a->3	
Art	i->3	
Asi	e->2	
Ass	a->2	
Ast	u->1	
Ata	t->2	
Atl	a->4	
Att	 ->28	a->1	
Aus	c->1	
Aut	o->1	
Auv	e->1	
Av 	4->1	a->5	b->2	d->15	e->1	o->1	s->2	t->1	v->2	
Avb	r->1	
Avf	a->1	
Avg	å->1	
Avi	a->1	
Avs	a->1	e->2	l->14	
Azo	r->2	
B A	l->1	
B o	c->1	
B t	a->1	
B-A	l->2	
B5-	0->4	
BAT	T->1	
BB 	A->1	
BB-	A->2	
BC 	d->1	
BI 	-->1	
BNI	 ->6	,->1	
BNP	 ->7	,->2	
BP,	 ->1	
BRÅ	D->1	
BSE	 ->2	-->4	
Bak	o->2	
Bal	f->1	k->7	
Ban	k->1	
Bar	a->13	c->2	e->1	n->15	ó->2	
Bas	k->2	s->1	
Bed	r->2	ö->2	
Bef	o->1	
Beh	r->7	
Bek	v->1	
Bel	g->9	
Ben	e->1	
Ber	e->14	g->13	l->7	n->5	o->1	t->2	
Bes	l->4	q->1	
Bet	r->7	ä->25	
Bev	i->1	
Big	 ->1	
Bil	i->1	l->2	t->2	
Bis	c->6	t->1	
Bla	k->1	n->8	
Blo	k->1	
Boe	t->1	
Bol	k->1	
Bon	d->1	
Bor	d->4	t->1	
Bos	ä->1	
Bou	r->6	
Bow	e->2	i->2	
Bra	n->2	s->1	v->1	
Bre	m->1	t->8	
Bri	s->3	t->2	
Bro	k->9	
Bru	n->1	
Bry	s->19	
Bud	a->1	g->1	
Bul	g->1	
Bus	h->1	q->1	
Byg	g->1	
Byr	n->2	å->1	
Bäs	t->1	
Båd	a->5	
C d	e->1	
C, 	a->1	
C-l	e->1	
C. 	D->1	E->1	
C.V	i->1	
C4-	0->6	
C5-	0->22	
CAF	:->1	
CEC	A->1	
CEN	 ->4	)->2	,->2	:->4	
CER	N->1	
CES	)->1	-->3	
CH 	B->1	
CHO	 ->1	,->1	.->1	
CK 	n->1	
CLA	F->1	
CM.	A->1	
CNS	)->9	
COD	)->13	
COS	)->2	
CSU	-->1	:->2	
Cad	i->5	o->1	
Cam	r->1	u->1	
Can	a->1	d->1	y->3	
Car	p->1	t->1	
Cas	a->2	
Cau	d->1	
Cav	a->1	
Cen	t->13	
Cer	m->1	
Cey	h->1	
Cha	m->1	
Chi	q->1	
Cla	u->1	
Cli	n->1	
Coc	a->1	i->1	
Col	a->1	
Con	a->1	s->1	
Cor	b->1	p->1	
Cos	t->9	
Cou	n->1	
Cox	 ->2	!->1	,->1	
Cre	s->2	
Cun	h->1	
Cur	i->1	
Cus	í->1	
Cux	h->1	
Cyp	e->1	
D b	ö->1	
D f	ö->1	
D k	r->1	
D))	 ->4	(->4	.->3	H->1	
D)]	.->1	
D, 	o->1	
D-g	r->2	
DA)	 ->2	
DD,	 ->1	
DD-	g->2	
DDR	.->1	
DE 	F->1	
DE)	 ->3	.->1	
DE-	 ->2	g->4	l->1	
DEB	A->1	
DR 	a->1	
DR)	 ->1	
DR-	g->1	
DR.	S->1	
DR:	s->1	
DSK	A->1	
Da 	C->3	
Dag	e->5	l->2	m->1	
Dal	a->7	
Dam	 ->2	a->1	
Dan	m->26	
Dar	m->1	
Dav	i->3	
De 	1->2	G->1	P->1	R->1	a->8	b->5	d->5	e->2	f->22	g->10	h->12	i->1	k->12	l->2	m->7	n->8	o->3	p->4	r->1	s->26	t->7	u->4	v->3	ä->4	å->2	
Del	g->1	o->3	s->1	v->1	
Dem	i->1	o->1	
Den	 ->211	n->57	
Der	a->2	
Des	s->61	
Det	 ->903	,->1	a->1	s->1	t->211	
Deu	t->1	
Dim	i->5	
Dir	e->9	
Dis	k->1	
Doc	k->2	
Dok	u->1	
Dom	s->3	
Dor	i->1	
Dub	l->7	
Duh	a->1	
Dui	s->3	
Dut	r->1	
Där	 ->15	a->2	e->10	f->96	i->3	m->4	u->1	v->1	
Då 	b->1	d->1	f->3	g->1	h->2	k->7	m->1	o->1	s->2	t->1	v->2	ä->2	ö->1	
Díe	z->1	
Düh	r->1	
E F	R->1	
E h	a->2	
E o	c->2	
E t	i->1	
E ä	r->1	
E) 	H->1	J->1	Ä->1	
E).	(->1	
E)J	a->1	
E- 	o->2	
E-D	E->8	
E-g	r->12	
E-k	o->1	r->3	
E-l	e->1	
E-t	e->1	
E/N	G->2	
EBA	T->1	
ECA	F->1	
ECH	O->3	
EDD	,->1	-->2	
EEG	 ->1	,->2	
EG 	a->1	o->2	s->1	t->2	u->1	
EG,	 ->7	
EG-	d->24	f->8	i->1	k->16	r->3	
EG.	V->1	
EG:	s->3	
EG?	,->1	
EIF	 ->1	)->1	
EK 	(->1	
EK(	1->3	9->1	
EKS	G->8	
EL)	 ->3	
ELD	R->3	
ELL	A->1	
EM-	2->1	
EMU	,->1	-->2	:->3	
EN 	e->1	h->1	k->1	o->1	
EN)	 ->36	
EN,	 ->2	
EN-	g->1	
EN:	s->4	
EO 	b->2	ä->1	
EP 	(->1	r->1	
ERN	)->1	
ERR	E->3	
ES)	 ->2	
ES-	z->3	
EU 	"->1	I->1	a->3	b->2	d->1	f->1	g->2	h->2	i->4	k->3	m->3	o->4	p->1	r->1	s->6	u->2	ä->2	
EU,	 ->5	
EU-	b->2	e->1	f->6	g->1	i->5	k->6	l->5	m->6	n->1	o->1	p->2	r->2	s->3	t->1	u->1	v->1	
EU.	.->1	A->1	D->3	F->1	N->1	R->1	V->3	
EU:	s->44	
EU?	H->1	
EUG	F->3	
Ece	m->1	
Edi	n->1	
Eff	e->5	
Eft	a->2	e->48	
Egy	p->2	
Ehu	d->2	
Eie	c->1	
Eko	f->2	n->3	
Eli	s->1	
Ell	e->4	
Elm	a->2	
Els	t->1	
Eme	l->8	
Emi	l->1	
En 	a->16	b->4	d->7	f->4	g->1	k->5	m->2	p->2	r->4	s->9	u->1	v->10	ö->2	
Enb	a->1	
End	a->11	
Enk	e->1	
Enl	i->37	
Equ	a->8	q->2	
Er 	a->1	
Era	 ->1	
Erf	a->2	
Eri	k->29	t->1	
Erk	k->2	
Ert	 ->2	
Eti	o->3	
Ett	 ->48	
Eur	a->4	o->847	
Eva	n->7	
Eve	n->1	
Exc	e->1	
Exe	m->1	
Exp	e->2	
Exu	p->1	
Exx	o->3	
F g	ö->1	
F h	a->1	
F i	 ->2	
F k	a->1	o->1	
F s	k->1	
F) 	ä->1	
F),	 ->1	
F, 	E->1	d->1	e->1	k->1	s->2	v->1	ö->1	
F.A	l->1	
F.F	ö->1	
F.H	e->1	
F.M	e->1	
F:s	 ->2	
FAF	,->1	
FBI	 ->1	
FEO	 ->3	
FI)	 ->1	
FIL	,->1	
FIP	O->1	
FJ)	 ->1	,->1	
FJ:	s->1	
FMI	 ->1	
FN,	 ->1	
FN-	u->1	
FN.	H->1	
FN:	s->8	
FOP	)->1	
FPÖ	 ->12	)->1	-->2	:->4	
FR)	 ->18	
FRÅ	G->1	
FSR	 ->1	
FUF	)->1	
Fac	k->3	t->1	
Fak	t->4	
Far	l->1	o->1	
Fas	c->1	
Fei	r->2	
Fel	a->1	
Fem	 ->1	
Fin	a->6	l->6	n->4	
Fir	m->1	
Fis	c->4	
Fla	u->2	
Fle	r->4	
Flo	r->19	
Flé	c->1	
FoU	,->1	-->1	
Fog	 ->1	
Fol	k->6	
Fon	t->1	
For	d->1	e->1	s->2	
Fra	g->1	m->9	n->49	s->1	
Fre	d->1	
Fri	h->3	
Fru	 ->82	t->3	
Frä	m->2	
Frå	g->42	n->2	
Fun	d->1	
Fyr	t->1	
Fäs	t->1	
Får	 ->3	
Föl	j->6	
För	 ->186	b->5	d->3	e->55	f->1	h->4	i->2	l->1	m->1	o->1	p->1	s->39	t->2	u->7	v->4	ä->1	
G a	t->1	
G o	m->2	
G s	k->1	
G t	i->2	
G u	p->1	
G(P	a->1	
G, 	E->6	f->1	o->1	v->1	
G-d	i->2	o->22	
G-f	ö->14	
G-i	n->1	
G-k	o->16	
G-r	ä->3	
G.(	E->1	
G.V	i->1	
G:s	 ->3	
G?,	 ->1	
GA-	s->1	
GAS	P->1	
GFJ	)->2	:->1	
GL-	g->2	
GOR	N->1	
GUE	/->2	
GUS	P->1	
Gal	e->1	i->2	
Gam	a->3	
Gar	g->5	
Gaz	a->6	
Gem	e->6	
Gen	e->10	o->28	è->3	
Ger	 ->1	
Gil	-->2	
Gin	o->1	
Giv	e->2	
Goe	b->1	
Gol	a->9	f->3	l->1	
Gom	e->1	
Gon	z->1	
Goo	d->1	
Gor	s->1	
Got	t->1	
Gra	c->4	t->1	ç->5	
Gre	k->14	
Gro	s->3	
Gru	n->1	p->10	
Grö	n->2	
Gua	t->1	
Gui	g->1	
Gul	f->1	
Gus	p->1	
Gut	e->2	
Gäl	l->1	
Gå 	h->1	
Gör	 ->2	
Göt	e->1	
H B	R->1	
H-0	0->1	7->12	8->8	
HO 	i->1	
HO,	 ->1	
HO.	D->1	
Haa	r->1	
Had	e->3	
Hag	u->1	
Hai	d->37	
Ham	b->1	
Han	 ->18	d->4	s->3	
Har	 ->11	r->1	
Hat	z->2	
Hav	e->1	
Hea	t->1	
Heb	r->1	
Hed	g->1	k->1	
Hei	n->2	
Hel	a->3	i->1	s->20	t->2	
Hem	l->1	
Hen	r->1	
Her	r->329	
Hic	k->1	
Hil	t->1	
Him	a->1	
His	t->2	
Hit	 ->3	l->6	t->3	
Hol	l->1	z->2	
Hon	 ->4	
Hop	p->1	
How	i->1	
Huh	n->1	
Hul	t->25	
Hur	 ->35	u->1	
Huv	u->7	
Hyc	k->1	
Hän	d->2	s->2	
Här	 ->33	m->2	o->1	
Hål	l->1	
Hög	e->1	
I -	 ->4	
I A	m->1	
I E	u->4	
I F	r->2	
I H	e->1	
I I	r->2	t->1	
I N	e->1	
I R	a->1	
I S	c->1	
I T	i->1	u->1	y->1	
I a	l->3	n->3	p->1	r->1	v->3	
I b	e->6	u->1	ö->2	
I d	a->24	e->60	i->1	ä->1	
I e	g->7	n->11	r->1	t->2	
I f	j->1	l->1	o->1	r->6	ö->6	
I g	å->3	
I h	a->2	
I i	 ->3	
I j	u->1	
I k	l->1	o->3	r->1	
I l	i->7	
I m	e->1	i->2	o->6	å->1	
I n	o->2	ä->2	
I o	c->8	k->1	
I p	a->1	e->2	r->2	
I r	a->2	e->8	ä->1	å->1	
I s	a->3	i->3	j->4	k->1	l->3	t->11	y->2	å->4	
I t	j->1	
I u	p->1	t->2	
I v	a->2	e->1	i->7	o->1	ä->2	å->6	
I ä	n->1	
I ö	v->3	
I) 	J->1	o->1	
I);	 ->1	
I, 	e->1	h->1	
I-p	r->3	
I. 	f->2	
I:e	 ->2	
ICE	S->4	
IF 	h->1	
IF)	,->1	
IFI	L->1	
IFO	P->1	
II 	-->2	h->2	i->1	k->1	s->1	
II)	 ->1	
II,	 ->1	
II-	p->2	
II.	 ->1	
II:	e->2	
III	 ->4	:->1	
IK,	 ->1	
IK.	D->2	
IL,	 ->1	
IMO	)->1	.->1	:->1	
INA	 ->2	,->1	
ING	(->1	.->1	
INT	E->4	
IPO	L->1	
IRA	 ->1	
ISP	A->1	
IT)	 ->3	
IV 	-->1	i->2	
IX 	o->1	
IX,	 ->1	
Ibl	a->3	
Idé	n->1	
Ihå	l->1	
Ile	-->1	
Ill	e->1	
Imb	e->3	
Imm	i->1	
Ind	i->5	u->1	
Inf	ö->4	
Ing	a->2	e->14	l->2	
Ini	t->3	
Inn	e->2	
Ino	m->10	
Inr	e->2	ä->1	
Ins	a->2	
Int	e->36	
Irl	a->22	
Isa	b->2	
Isl	a->1	
Isr	a->38	
Ist	a->1	
Ita	l->18	
Izq	u->1	
J) 	f->1	
J),	 ->1	
J:s	 ->1	
Ja 	E->1	e->1	t->1	
Ja,	 ->8	
Jac	k->2	o->2	q->3	
Jag	 ->953	
Jan	-->1	
Jap	a->3	
Jav	e->1	
Jea	n->1	
Jer	u->2	
Jo 	d->1	
Jo,	 ->3	
Jon	a->2	c->14	
Jor	d->4	
Jos	p->1	
Ju 	m->1	
Jug	o->1	
Jun	k->1	
Jus	t->10	
Jäm	f->2	s->1	
Jör	g->14	
Jør	g->2	
K (	d->1	
K n	u->1	
K(1	9->3	
K(9	9->1	
K, 	d->1	v->1	
K.D	e->2	
KAN	D->1	
KOM	(->10	
KSG	,->2	-->6	
KTU	E->1	
Kaf	o->1	
Kal	e->3	
Kan	 ->13	a->1	s->9	t->3	
Kar	a->3	l->7	t->2	
Kas	p->1	
Kat	a->1	
Kau	f->1	k->3	
Kaz	a->1	
Kee	s->1	
Kfo	r->1	
Kin	a->10	n->24	
Kir	g->5	
Kna	p->1	
Koc	h->15	
Kod	e->1	
Kol	l->1	
Kom	 ->1	m->120	p->1	
Kon	k->14	r->1	s->5	v->2	
Kor	e->2	t->2	
Kos	o->60	t->4	
Kou	c->12	
Kra	v->3	
Kul	t->25	
Kum	a->1	
Kun	g->1	
Kva	n->1	
Kvi	n->5	
Kvä	k->1	
Kyo	t->7	
Kän	n->1	
Kär	a->6	n->4	
Köl	n->2	
Köp	e->1	
L (	e->1	
L) 	A->1	F->1	H->4	J->1	
L),	 ->1	
L, 	f->1	
L-g	r->2	
LA 	O->1	
LAF	 ->6	,->7	.->4	:->1	
LAS	 ->1	
LDR	 ->1	-->1	:->1	
LFA	F->1	
LLA	 ->1	
LTC	M->1	
La 	R->2	
Laa	n->7	
Lam	a->7	
Lan	d->2	g->30	k->3	
Lap	p->2	
Le 	B->1	
Lea	d->5	
Led	a->4	n->1	
Lei	n->8	
Leo	n->1	
Lib	a->5	e->2	y->1	
Lii	k->3	
Lik	a->3	r->1	s->8	v->1	
Lil	l->1	
Lis	s->8	
Lit	a->1	t->1	
Liv	l->2	s->3	
Llo	y->1	
Loi	r->3	
Lom	é->2	
Lon	d->4	
Lor	d->2	r->2	
Lot	h->3	
Lou	s->1	
Loy	o->2	
Lut	t->1	
Lux	e->6	
Lyc	k->2	
Lyn	n->4	
Läg	g->2	
Län	d->1	
Lån	 ->1	g->1	
Låt	 ->61	
Löö	w->1	
M A	K->1	
M s	o->1	
M(1	9->8	
M(9	8->1	9->1	
M-2	0->1	
M.A	t->1	
MAR	P->1	
MI 	d->1	
MIK	,->1	.->2	
MO)	.->1	
MO.	D->1	
MO:	s->1	
MRÖ	S->2	
MU,	 ->1	
MU-	a->1	k->1	
MU:	s->3	
Maa	s->6	
Mac	a->1	
Mad	a->1	e->2	r->3	
Mai	n->1	
Maj	o->1	
Mal	t->7	
Man	 ->56	n->2	
Mar	g->2	i->8	k->5	p->1	s->1	t->1	
Mat	h->2	
Max	i->2	
McC	a->1	
McN	a->5	
Med	 ->35	a->4	b->3	e->3	g->1	l->9	
Mel	l->20	
Men	 ->209	,->3	a->1	t->1	
Mer	 ->3	
Mex	i->1	
Mic	h->1	
Mid	d->1	l->1	
Mil	j->1	
Min	 ->32	a->18	d->1	i->1	n->1	s->1	u->1	
Mis	t->2	
Mit	r->1	t->5	
Mon	t->19	
Mor	a->5	b->1	g->4	
Mos	k->1	
Mot	 ->8	
Mou	r->8	s->1	
Mul	d->1	
Myc	k->1	
Myl	l->1	
Myn	d->3	
Män	n->5	
Mär	k->1	
Måh	ä->1	
Mål	e->2	
Mån	g->10	
Möj	l->2	
Mün	c->1	
N e	l->1	
N h	a->1	
N k	o->1	
N o	c->1	
N) 	D->2	F->6	H->4	I->3	J->7	K->1	L->2	M->1	S->1	T->4	U->1	V->2	i->2	s->1	
N))	.->1	
N, 	a->1	s->2	
N-g	r->1	
N-u	p->1	
N.H	e->1	
N:s	 ->12	
NA 	h->1	v->1	
NA,	 ->1	
NDE	 ->1	
NG(	P->1	
NG.	(->1	
NGL	-->2	
NI 	b->1	i->1	o->2	p->2	
NI,	 ->1	
NIF	I->1	
NIN	G->2	
NL)	 ->4	
NMI	K->3	
NP 	j->1	m->1	p->4	å->1	
NP,	 ->2	
NS)	)->9	
NTE	 ->1	R->3	
Nal	l->5	
Nan	a->1	
Nap	o->1	
Nar	k->1	
Nat	i->7	o->5	u->15	
Ned	e->9	
Nej	,->7	.->1	
New	 ->1	
Ni 	a->1	b->4	f->3	h->11	k->9	l->1	m->4	n->1	s->6	t->2	v->3	
Nie	l->6	
Nik	i->2	
Niv	å->1	
Nog	u->1	
Noi	r->1	
Nor	d->3	g->2	m->2	
Nu 	a->2	b->1	f->3	h->7	k->2	m->1	t->1	v->2	ä->7	å->1	
Num	e->1	
Nuv	a->1	
Nya	 ->3	
Nyl	i->1	
Nyt	t->1	
När	 ->83	
Näs	t->26	
Någ	o->3	r->2	
Nåj	a->1	
Nöd	v->1	
O b	e->2	
O i	 ->1	
O ä	r->1	
O).	F->1	
O, 	a->1	
O.D	e->2	
O:s	 ->1	
O?E	n->1	
OCH	 ->1	
OD)	)->12	]->1	
OFS	R->1	
OK,	 ->1	
OL 	(->1	
OL)	,->1	
OLA	F->17	S->1	
OLF	A->1	
OM 	A->1	
OM(	1->8	9->2	
OMR	Ö->2	
OP)	.->1	
ORN	ä->1	
OS)	]->2	
OSS	E->1	
Oav	s->2	
Obe	r->3	
Och	 ->67	:->1	
Ock	s->2	
Off	e->3	i->1	
Oft	a->1	
Oil	 ->1	-->1	
Oli	k->1	v->1	
Olj	e->3	
Oly	m->1	
Om 	5->1	E->2	S->2	a->3	b->1	d->23	e->5	f->1	g->2	i->4	j->2	k->5	l->1	m->11	n->8	o->1	p->2	r->2	s->2	t->2	u->1	v->23	
Oma	g->1	
Omr	ö->15	
One	s->1	
Onö	d->1	
Ora	n->1	
Ord	 ->1	e->3	f->7	
Ork	a->2	
Oro	n->1	v->1	
Ors	a->2	
Osl	o->3	
Osm	a->1	
Ouv	r->1	
Oz 	d->1	h->1	
Oz,	 ->1	
P (	"->1	Ö->2	
P a	t->2	
P j	ä->1	
P m	i->2	å->1	
P o	c->1	
P p	e->3	å->1	
P r	e->1	
P å	r->1	
P) 	o->1	
P).	V->1	
P, 	e->1	i->1	m->1	
PA-	i->1	
PE 	h->1	ä->1	
PE-	D->8	g->5	
PM 	s->1	
POL	 ->1	)->1	
PPE	 ->2	-->13	
PR-	e->1	
PSE	)->1	-->3	
PT)	 ->16	
PVC	,->1	-->1	.->1	
Pac	k->3	
Pad	d->2	
Pak	i->5	
Pal	a->15	e->11	
Pap	a->2	
Par	a->1	i->3	l->42	
Pat	t->23	
Pay	s->2	
Pea	k->1	
Pei	j->2	
Pek	i->1	
Per	s->4	
Pet	e->1	r->1	
Pla	n->2	s->2	t->5	
Plo	o->1	
Plä	d->1	
Poe	t->5	
Poh	j->1	
Pol	e->1	l->1	
Pom	é->1	
Pon	n->1	
Poo	s->1	
Por	t->27	
Pow	e->3	
Pre	c->6	s->1	u->1	
Pri	o->1	
Pro	b->9	c->3	d->30	g->1	j->2	t->2	v->3	
Prí	n->1	
Pun	k->2	
Pur	v->1	
PÖ 	(->2	f->1	h->1	i->1	m->1	o->4	s->1	v->1	ä->1	
PÖ)	 ->1	.->1	
PÖ-	l->1	m->1	
PÖ:	s->4	
På 	a->1	d->22	e->1	g->2	l->1	m->3	o->2	p->1	s->11	u->1	v->3	
Pås	t->1	
Pét	a->1	
Que	c->1	
R -	 ->1	
R a	n->1	
R) 	"->1	D->4	E->1	F->1	H->1	I->2	J->4	N->3	T->1	o->1	
R-e	f->1	
R-g	r->1	
R.S	e->1	
R:s	 ->1	
RA 	h->1	
REG	,->1	-->1	?->1	
REP	 ->2	
RIN	A->3	
RN)	 ->1	
RNä	s->1	
RPO	L->1	
RRE	G->3	
Rac	k->2	
Raf	a->3	
Ran	d->4	
Rap	k->11	p->3	
Ras	c->1	i->1	
Rea	d->1	k->1	
Red	a->3	i->8	
Ref	o->7	
Reg	e->6	i->1	
Ren	t->2	
Rep	u->1	
Res	t->2	u->5	
Ret	r->1	
Rev	i->4	
Rhô	n->1	
Ric	h->3	
Rii	s->2	
Rik	a->1	t->4	
Rio	f->1	
Ris	k->1	
Rob	e->1	l->1	
Roi	s->1	
Roj	o->1	
Rom	-->1	a->3	á->1	
Roo	 ->1	
Rop	e->1	
Rot	h->7	t->2	
Rov	e->2	
Roy	a->1	
Rui	z->1	
Rum	ä->1	
Rus	h->1	
Rys	s->4	
RÅD	S->1	
RÅG	O->1	
RÖS	T->2	
Räk	n->1	
Rät	t->2	
Råd	e->21	s->1	
Réu	n->2	
Rös	t->1	
S (	I->1	
S o	c->1	
S) 	-->1	ä->1	
S))	 ->1	(->4	.->2	F->1	o->1	
S)]	.->2	
S-z	o->3	
S:s	 ->1	
SA 	-->1	a->1	e->1	h->1	p->1	
SA,	 ->2	
SA.	J->1	V->1	
SA:	s->1	
SD 	f->1	
SE 	o->2	t->1	
SE)	J->1	
SE-	g->3	k->3	t->1	
SEK	 ->1	(->4	
SEM	-->1	
SG,	 ->2	
SG-	f->6	
SKA	N->1	
SOL	A->1	
SP 	m->1	o->1	
SPA	-->1	
SPÖ	 ->1	)->1	
SR 	-->1	
SS 	o->1	
SS:	s->1	
SSE	 ->1	
STN	I->2	
SU-	g->1	
SU:	s->2	
SYN	)->1	
Sag	e->1	
Sai	n->1	
Sal	a->1	
Sam	h->2	m->26	o->1	t->14	
San	 ->1	n->6	t->3	
Sav	e->9	
Sch	e->10	r->18	u->3	w->2	ö->1	ü->4	
Sea	t->4	
Seb	a->1	
Sed	a->20	
Seg	n->1	u->1	
Sei	x->5	
Ser	i->1	
Set	t->1	
Sha	r->6	
She	i->5	l->2	p->3	
Sim	p->1	
Sis	t->2	
Sit	u->3	
Sju	 ->1	k->1	
Sjä	l->2	t->1	
Sjö	s->4	
Ska	d->1	l->4	
Sko	g->1	t->5	
Sku	l->8	
Sky	d->1	
Skä	l->1	
Slo	v->1	
Slu	t->38	
Små	 ->1	f->1	
Sna	b->1	r->1	
Soa	r->1	
Soc	i->4	
Sok	r->1	
Sol	a->4	b->2	
Som	 ->53	l->3	
Sou	l->1	
Spa	n->7	
Spe	n->1	r->1	
Sri	 ->3	
St.	V->1	
Sta	b->1	d->1	t->9	
Sto	c->3	r->18	
Str	a->7	u->1	ä->1	
Stä	m->1	
Stå	l->1	
Stö	d->7	r->4	
Sua	n->1	
Sub	v->2	
Sud	r->2	
Sva	r->1	
Sve	p->1	r->7	
Swo	b->3	
Syd	a->2	k->1	o->2	
Syf	t->6	
Syr	i->24	
Sán	c->1	
São	 ->2	
Säg	 ->1	
Säk	e->2	
Sär	s->2	
Så 	b->1	d->3	e->2	f->1	h->1	j->3	k->2	l->5	n->1	r->1	s->4	t->1	v->6	ä->3	
Såd	a->2	
Sål	e->4	
Sån	g->1	
Sås	o->2	
Såv	ä->1	
Söd	e->2	
T O	M->1	
T) 	D->1	E->1	F->1	H->10	J->2	L->1	N->1	O->1	V->1	
TCM	.->1	
TE 	h->1	
TER	R->3	
TNI	N->2	
TO?	E->1	
TT 	O->1	
TUE	L->1	
TV 	a->1	
TV-	b->1	k->1	p->1	s->1	
Ta 	d->1	
Tac	i->2	k->38	
Tad	z->5	
Tai	w->1	
Tal	a->1	m->9	
Tam	m->22	
Tan	g->1	i->1	k->3	
Tau	e->1	
Ter	r->4	
Tes	a->1	
Tex	a->2	
The	a->21	
Thy	s->5	
Tib	e->21	
Tid	i->1	n->1	
Til	l->49	
Tit	t->1	
Tod	i->1	
Tom	 ->1	é->2	
Ton	g->1	
Top	p->2	
Tor	r->3	v->2	
Tot	a->6	
Tra	n->3	
Tre	 ->1	d->1	
Tri	t->1	
Tro	r->2	t->17	v->1	
Trä	d->1	
Tsa	t->3	
Tur	k->37	
Tus	e->1	
Tvä	r->4	
Två	 ->2	
Ty 	e->1	h->1	i->1	s->1	u->1	v->3	
Tyc	k->1	
Tyd	l->1	
Tys	k->20	
Tyv	ä->9	
Tän	k->2	
Tåg	k->1	
U "	c->1	
U I	 ->1	
U a	g->1	t->2	
U b	l->1	ö->1	
U d	ä->1	
U f	r->1	
U g	e->1	ö->1	
U h	a->2	
U i	 ->1	n->3	
U k	a->3	
U m	e->1	y->1	å->1	
U o	c->4	
U p	å->1	
U r	e->1	
U s	k->1	o->4	y->1	
U u	t->2	
U ä	r->2	
U, 	f->1	l->1	m->1	n->1	p->1	t->1	v->1	
U-a	n->1	
U-b	i->1	u->1	
U-e	n->1	
U-f	o->1	ö->5	
U-g	e->1	r->1	
U-i	n->5	
U-k	o->6	r->1	
U-l	a->2	ä->3	
U-m	a->1	e->5	
U-n	i->1	
U-o	r->1	
U-p	r->2	
U-r	a->1	e->1	ä->1	
U-s	t->1	ä->2	
U-t	e->1	
U-u	t->1	
U-v	ä->1	
U..	 ->1	
U.A	l->1	
U.D	a->1	e->2	
U.F	r->1	
U.N	u->1	
U.R	o->1	
U.V	i->3	
U:s	 ->49	
U?H	e->1	
UCK	 ->1	
UCL	A->1	
UE/	N->2	
UEL	L->1	
UEN	-->1	
UF)	 ->1	
UGF	J->3	
UNI	F->1	
UNM	I->3	
USA	 ->5	,->2	.->2	:->1	
USD	 ->1	
USP	 ->1	
Uls	t->1	
Und	a->3	e->34	
Ung	d->1	e->2	
Uni	o->8	
Upp	d->1	e->1	f->1	g->3	r->1	
Ur 	d->2	e->1	p->1	
Urb	a->2	
Urq	u->1	
Urs	ä->1	
Uta	n->3	
Utb	i->2	
Utd	e->1	
Ute	s->1	
Utf	o->2	ö->1	
Utg	i->2	
Uti	f->1	
Utm	a->2	
Utn	ä->2	
Uts	k->6	
Utt	j->1	
Utv	e->1	i->1	ä->1	
Uzb	e->2	
V -	 ->2	
V a	n->1	
V i	 ->2	
V-b	i->1	
V-k	a->1	
V-p	r->1	
V-s	ä->1	
VC,	 ->1	
VC-	l->1	
VC.	V->1	
VD 	b->1	
VI 	i->1	
VII	:->1	I->3	
VP 	(->2	a->2	m->1	
VP)	 ->1	
Vad	 ->75	a->1	
Val	d->3	e->3	l->3	
Van	 ->3	d->1	l->1	
Vap	e->1	
Var	 ->7	e->3	f->12	j->7	k->1	
Vat	a->3	
Vel	z->1	
Vem	 ->7	s->2	
Ven	d->1	e->1	s->2	
Ver	h->2	k->1	s->1	
Vet	e->2	s->1	
Vi 	a->25	b->40	d->8	e->2	f->34	g->8	h->102	i->13	j->1	k->60	l->4	m->83	o->1	p->2	r->6	s->46	t->18	u->9	v->60	ä->35	ö->1	
Vi,	 ->1	
Via	 ->1	
Vic	h->1	
Vid	 ->14	a->7	
Vik	t->1	
Vil	j->1	k->24	l->5	
Vin	d->1	
Vis	s->16	
Vit	b->3	o->7	
Viv	i->1	
Vla	a->1	
Vod	a->1	
Vol	k->1	
Von	 ->1	
Vär	d->1	l->3	
Väs	t->6	
Vår	 ->16	a->8	t->7	
WTO	?->1	
Waf	f->2	
Wal	e->11	l->4	
Was	h->3	
Web	,->1	
Wes	t->1	
Wid	e->1	
Wie	b->1	l->4	n->4	
Wil	h->1	
Wog	a->18	
Wor	l->1	
Wul	f->2	
Wur	t->3	
Wye	 ->1	-->2	
Wyn	n->1	
X o	c->2	
X, 	f->1	
XVI	I->2	
XXV	I->2	
YN)	)->1	
Yas	s->1	
Yor	k->1	
Ytt	e->3	
Zee	l->2	
Zim	e->1	
[KO	M->2	
[SE	K->1	
].)	 ->1	
].H	e->2	
a "	A->1	b->1	i->1	l->1	s->1	u->1	
a (	K->1	a->1	
a -	 ->62	,->1	
a 1	 ->3	0->3	2->2	3->1	5->1	6->3	7->1	
a 2	 ->2	0->1	5->5	
a 3	0->1	3->1	5->1	7->1	
a 4	0->1	
a 5	 ->1	5->1	
a 6	 ->1	0->1	
a 7	0->1	
a 8	1->5	5->3	7->1	
a 9	0->1	
a A	h->1	l->3	m->1	t->1	z->1	
a B	 ->1	a->3	e->2	o->1	r->2	
a C	o->9	
a D	a->2	
a E	E->1	G->5	U->15	l->2	r->2	u->56	v->1	
a F	N->2	P->2	e->1	i->1	l->4	r->4	ö->1	
a G	o->1	r->2	
a H	a->6	i->1	u->1	
a I	X->1	n->1	s->2	z->1	
a J	a->1	e->2	o->1	ö->2	
a K	a->1	o->4	u->1	
a L	a->1	i->4	o->2	
a M	a->3	e->1	o->9	u->1	
a N	a->2	i->1	
a O	L->1	
a P	P->1	V->1	a->4	o->2	r->1	
a R	a->1	i->1	o->3	y->1	é->2	
a S	a->2	c->1	h->1	t->1	u->1	v->1	
a T	V->1	e->2	u->2	y->2	
a U	C->1	
a W	a->1	
a Z	e->2	
a a	b->3	d->5	f->3	g->6	k->13	l->73	m->8	n->176	p->2	r->102	s->19	t->481	u->2	v->242	
a b	a->30	e->366	i->92	j->1	l->29	o->27	r->31	u->24	y->11	ä->13	å->9	ö->26	
a c	a->1	e->14	h->5	i->2	
a d	a->64	e->909	i->99	j->7	o->32	r->20	u->4	y->4	ä->20	å->6	ö->6	
a e	f->49	g->28	k->35	l->54	m->17	n->434	r->71	t->186	u->35	v->3	x->25	
a f	a->126	e->11	i->31	l->20	o->119	r->437	u->20	y->1	ä->2	å->38	ö->899	
a g	a->21	e->131	i->18	j->6	l->6	n->1	o->15	r->133	ä->30	å->47	ö->35	
a h	a->218	e->46	i->26	j->6	o->27	u->44	y->3	ä->71	å->23	ö->28	
a i	 ->419	.->3	a->2	b->1	c->2	d->16	f->5	g->13	h->18	k->1	l->2	m->5	n->428	r->1	s->3	t->14	v->1	
a j	a->6	o->17	u->9	ä->9	
a k	a->118	e->2	i->2	l->33	n->5	o->566	r->77	u->42	v->37	y->1	ä->33	ö->2	
a l	a->52	e->39	i->73	j->2	o->12	u->3	y->5	ä->103	å->5	ö->30	
a m	a->64	e->500	i->147	o->58	u->4	y->102	ä->30	å->143	ö->66	
a n	a->47	e->13	i->21	o->15	r->26	u->5	y->46	ä->62	å->81	ö->13	
a o	a->1	b->14	c->559	d->2	e->3	f->19	g->1	i->1	j->2	k->4	l->34	m->430	n->3	p->9	r->176	s->65	t->1	
a p	a->134	e->50	h->1	i->1	l->29	o->90	r->253	u->80	å->228	
a r	a->68	e->377	i->60	o->8	u->27	y->1	ä->98	å->46	ö->33	
a s	.->1	a->168	c->4	e->67	i->304	j->26	k->214	l->46	m->13	n->13	o->261	p->42	t->386	u->16	v->31	y->82	ä->131	å->53	ö->2	
a t	.->2	a->82	e->51	i->366	j->27	o->24	r->66	u->6	v->34	y->39	ä->6	å->2	
a u	l->1	m->1	n->338	p->198	r->16	t->228	
a v	a->142	e->107	i->198	o->6	r->2	ä->96	å->52	
a y	r->3	t->16	
a Ö	s->6	
a ä	g->10	m->20	n->109	r->307	v->10	
a å	 ->2	k->8	r->60	s->9	t->147	
a ö	a->3	d->2	g->6	k->10	n->7	p->6	r->2	s->6	v->82	
a! 	D->1	V->1	
a!A	v->1	
a!D	e->4	
a!F	r->3	ö->1	
a!H	e->2	
a!J	a->1	
a!L	å->1	
a!M	ä->1	
a!O	m->1	
a!Ä	v->1	
a" 	b->1	s->1	v->1	
a",	 ->1	
a".	.->1	B->1	D->2	H->1	J->1	K->1	
a";	 ->1	
a"i	n->1	
a) 	a->1	b->1	
a, 	1->1	5->1	B->1	E->1	J->1	K->1	S->2	a->36	b->11	c->1	d->54	e->36	f->55	g->5	h->36	i->39	j->6	k->16	l->11	m->57	n->18	o->106	p->10	r->12	s->89	t->23	u->26	v->47	ä->13	å->4	ö->2	
a-,	 ->1	
a-I	s->1	
a-R	o->1	
a-o	l->1	
a. 	1->1	D->4	E->1	F->1	H->1	J->1	K->2	M->3	S->1	V->2	a->2	b->1	d->1	e->2	f->5	g->2	i->2	k->1	m->1	n->3	o->2	p->1	s->3	u->1	v->1	Å->1	
a.(	I->1	P->1	T->2	
a.)	B->1	F->1	
a.-	 ->4	
a..	 ->2	(->3	.->2	
a.1	8->1	
a.A	l->10	m->1	n->3	v->5	
a.B	a->2	e->5	i->1	l->1	o->1	
a.C	o->1	
a.D	e->155	o->1	ä->14	å->2	
a.E	G->1	f->8	m->3	n->13	t->8	u->4	
a.F	a->2	r->8	ö->26	
a.G	e->2	i->1	
a.H	a->2	e->34	u->4	ä->4	
a.I	 ->33	b->2	n->7	
a.J	a->98	u->2	
a.K	a->2	o->12	ä->2	
a.L	i->2	ä->1	å->6	
a.M	a->4	e->38	i->10	å->2	
a.N	a->2	i->6	u->3	ä->10	
a.O	c->9	m->11	r->2	
a.P	a->1	e->1	r->4	å->11	
a.R	e->2	u->1	å->2	
a.S	a->1	e->2	i->2	j->1	k->1	l->3	m->1	o->6	t->3	y->1	ä->1	å->4	
a.T	a->3	i->2	o->1	r->5	y->1	
a.U	n->4	p->2	r->1	t->5	
a.V	a->13	e->2	i->81	ä->2	å->3	
a.Ä	n->3	r->3	v->5	
a.Å	 ->2	r->1	
a.Ö	v->1	
a/E	u->1	
a/h	a->1	
a/s	a->1	
a: 	"->2	D->1	F->2	I->2	J->2	N->1	V->2	a->2	d->1	g->1	h->2	m->1	o->1	r->1	s->1	u->3	v->5	Ä->1	
a:F	ö->1	
a; 	d->1	e->1	f->2	j->2	k->1	l->1	o->1	p->1	v->2	
a?"	J->1	
a?.	 ->1	
a?A	n->1	v->1	
a?D	e->8	
a?E	t->1	
a?F	r->1	ö->1	
a?H	a->1	e->1	u->1	
a?I	 ->2	n->1	
a?J	a->3	o->1	
a?M	a->1	
a?N	e->1	ä->1	
a?P	r->1	å->1	
a?S	v->1	
a?V	a->3	i->4	
a?Ä	r->1	
aHe	r->1	
aNä	s->2	
aaf	f->1	
aam	s->1	
aan	 ->1	.->1	s->5	
aar	d->1	
aas	t->6	
ab 	s->1	
aba	r->1	s->1	
abb	 ->4	a->74	t->43	v->1	
abe	h->7	k->1	l->40	r->1	t->2	
abi	l->25	n->3	s->7	
abl	a->15	e->13	o->1	
abo	c->2	n->8	r->3	
abr	e->1	i->4	
abs	o->41	t->3	u->3	
abu	 ->1	k->2	l->1	
abv	ä->1	
ac 	b->2	o->1	
ac"	,->1	
ac-	s->1	
aca	 ->4	o->1	
acc	e->88	
ace	 ->1	.->2	r->17	u->1	
aci	l->1	o->15	s->2	t->5	
ack	 ->56	,->15	-->1	.->3	a->108	d->8	e->3	f->7	l->2	n->6	o->1	r->6	s->12	
aco	-->1	b->2	
acq	u->4	
act	o->1	
acè	t->1	
ad 	-->1	A->1	B->1	E->1	F->1	G->1	K->2	S->1	a->47	b->37	d->39	e->17	f->33	g->66	h->10	i->28	j->14	k->34	l->1	m->32	n->7	o->36	p->19	r->11	s->103	t->19	u->7	v->38	y->1	ä->14	ö->19	
ad,	 ->20	
ad-	k->1	
ad.	"->1	(->1	D->7	E->1	F->1	H->6	J->4	K->2	M->6	O->14	P->1	R->1	S->1	U->1	V->3	
ad:	 ->1	
ad;	 ->1	
ad?	D->1	H->1	V->1	
ada	 ->13	!->1	,->3	.->1	d->2	g->1	k->1	n->4	r->6	t->4	
add	a->1	e->3	i->3	
ade	 ->747	,->27	.->32	:->1	?->1	e->2	f->1	i->2	k->5	l->2	m->4	n->167	r->184	s->119	t->3	
adg	a->28	o->1	
adi	e->4	k->16	n->2	o->2	t->19	u->4	z->5	
adj	e->2	
adk	o->24	
adl	i->11	
adm	i->28	
ado	,->1	r->26	u->1	x->6	
adr	a->3	i->4	
ads	 ->1	-->4	/->1	a->5	b->5	c->1	d->1	e->18	f->5	i->3	k->1	l->2	m->2	n->1	o->2	p->6	s->3	t->1	u->1	v->3	
adt	,->1	
adv	i->3	o->5	
adz	j->5	
adö	r->1	
ael	 ->24	,->4	-->1	.->4	?->1	e->5	i->15	k->1	s->6	
af 	o->1	
afa	e->3	t->1	
afe	t->1	
aff	 ->2	,->1	-->2	a->29	b->1	e->3	l->1	p->2	r->28	ä->12	
afi	 ->1	.->2	k->9	n->1	s->10	
afl	y->1	
afo	n->1	r->1	
afr	a->1	i->2	y->2	å->12	
aft	 ->72	,->11	.->6	?->2	e->26	f->12	i->34	o->1	s->10	t->5	v->8	
ag 	-->11	1->19	2->7	3->5	4->8	5->2	6->2	G->1	I->1	a->209	b->81	c->2	d->31	e->37	f->184	g->49	h->218	i->139	j->4	k->126	l->25	m->84	n->34	o->84	p->32	r->44	s->358	t->322	u->68	v->342	Ö->1	ä->122	å->7	ö->13	
ag,	 ->109	
ag.	 ->3	(->1	)->3	.->1	A->3	B->2	D->23	E->3	F->8	G->1	H->8	I->7	J->14	K->4	L->2	M->3	O->2	P->1	R->2	S->3	T->2	U->1	V->9	
ag:	 ->2	D->1	
ag;	 ->1	
ag?	D->1	F->3	
aga	 ->18	!->1	,->2	.->3	d->5	n->229	r->168	s->8	t->5	v->3	
agb	a->15	
agd	 ->4	,->1	a->7	
age	 ->2	d->4	l->6	m->9	n->224	r->73	s->1	t->215	
agf	ö->5	
agg	 ->6	,->7	.->5	;->1	a->5	e->2	n->1	o->1	r->1	
agh	 ->1	e->12	
agi	n->1	s->6	t->129	v->3	
agl	i->35	
agm	a->2	
agn	 ->3	a->36	e->12	i->71	
ago	g->5	l->4	m->4	r->57	s->1	
agr	a->6	e->1	o->1	u->1	
ags	 ->35	,->2	.->1	a->6	b->2	d->1	e->5	f->5	g->10	i->1	j->2	k->2	l->3	m->2	n->2	r->7	s->4	t->134	ä->3	
agt	 ->74	,->9	.->2	e->2	s->38	
agu	e->1	
agå	n->10	
aha	n->1	
ahu	s->1	
ahå	l->43	
ai 	L->7	
aid	e->37	s->5	
ail	 ->1	l->1	u->1	
ain	"->1	,->1	e->3	s->32	t->1	
air	e->1	
aiv	a->1	i->1	
aiw	a->1	
aj 	1->3	2->1	f->1	
aj,	 ->1	
aj.	J->1	T->1	
ajo	r->42	u->1	
ak 	a->4	b->2	f->1	g->3	h->5	i->2	j->1	k->2	l->1	m->5	n->1	s->12	t->3	u->1	v->6	ä->2	ö->1	
ak,	 ->6	
ak.	A->1	D->3	E->1	N->1	T->2	
ak:	 ->1	
ak?	N->1	
aka	 ->57	.->5	?->1	d->7	g->4	m->1	r->9	s->5	t->9	v->4	
akd	ö->1	
ake	,->1	l->3	n->15	r->45	t->10	
akf	ö->1	
akg	r->31	
aki	e->1	s->11	
akk	u->2	
akl	a->1	i->11	u->1	
akn	a->40	i->14	
ako	l->1	m->25	n->1	p->5	
akp	r->1	
akr	e->1	o->6	y->2	
aks	 ->4	a->9	o->1	t->1	
akt	 ->54	,->3	.->9	:->1	a->92	b->4	d->2	e->33	f->2	h->3	i->177	k->1	l->17	m->3	o->24	t->8	u->100	ä->9	ö->13	
aku	l->1	t->1	u->2	
akä	m->1	
akå	t->3	
al 	-->2	C->1	D->1	I->2	K->1	U->1	a->27	b->11	c->1	d->6	e->4	f->20	g->1	h->3	i->20	k->6	l->3	m->24	n->5	o->34	p->13	r->10	s->53	t->11	u->13	v->4	ä->7	å->3	ö->3	
al!	H->1	
al"	 ->2	
al,	 ->24	
al-	 ->7	F->3	S->1	s->2	
al.	 ->1	D->5	E->1	F->5	H->3	I->2	J->2	K->2	M->1	P->1	S->4	V->3	
al:	 ->2	
al;	 ->1	
alF	i->1	
ala	 ->332	"->1	,->5	.->8	?->3	c->15	d->35	f->1	g->5	i->7	m->1	n->93	r->122	s->17	t->33	y->1	
alb	a->19	e->3	l->1	
ald	 ->11	,->6	.->1	a->16	e->32	i->20	j->1	o->1	r->31	
ale	i->2	j->1	k->4	m->2	n->30	o->1	r->21	s->39	t->72	u->1	
alf	a->1	o->18	r->10	å->4	ö->11	
ali	b->2	c->2	e->41	f->15	g->5	n->4	s->146	t->72	
alj	 ->2	,->2	.->1	a->1	e->26	f->1	k->2	
alk	a->7	e->1	o->2	r->4	
all	 ->801	"->1	,->12	.->16	a->401	d->23	e->131	f->1	i->15	k->2	m->123	o->1	p->1	r->10	s->30	t->376	v->74	y->5	
alm	a->427	e->1	
aln	a->1	i->15	
alo	g->33	
alp	a->2	o->44	r->2	
alr	e->4	i->4	ä->1	
als	 ->27	.->1	e->2	f->1	k->9	l->1	o->1	p->7	r->1	s->1	t->5	u->1	y->1	
alt	 ->61	,->5	.->6	a->11	e->16	i->1	n->47	s->5	
alu	f->1	n->3	t->25	
alv	 ->4	a->4	e->1	h->1	i->1	m->1	o->2	t->5	v->2	å->5	ö->3	
aly	d->3	s->60	
alö	s->1	
am 	"->1	-->5	1->1	8->1	D->1	a->10	b->7	c->1	d->24	e->59	f->48	g->4	h->10	i->18	k->4	l->6	m->19	n->7	o->15	p->12	r->11	s->39	t->51	u->4	v->11	ä->5	å->3	ö->4	
am!	D->1	
am,	 ->36	
am.	.->1	D->5	F->4	G->2	H->2	I->1	J->2	K->2	M->2	N->2	O->1	R->1	S->3	T->1	V->2	
am?	J->1	V->1	
ama	 ->6	.->2	f->1	n->1	r->91	s->3	t->6	v->3	
amb	a->49	i->26	u->3	
ame	-->1	l->1	n->675	r->58	t->2	x->2	
amf	a->1	i->1	u->5	ö->179	
amg	i->1	å->52	
amh	e->97	ä->54	å->17	ö->2	
ami	d->1	k->1	l->15	n->21	s->4	
amk	a->4	o->10	
aml	a->61	e->1	i->27	ä->8	
amm	 ->1	a->590	e->133	
amn	 ->11	,->2	.->3	a->28	b->1	e->4	i->3	k->2	u->4	
amo	,->1	d->2	r->38	t->74	
amp	 ->11	a->7	e->19	l->8	o->1	r->12	å->1	
amr	a->1	e->2	u->1	ä->1	å->9	
ams	 ->1	k->6	t->52	y->3	
amt	 ->101	,->2	.->3	a->21	i->174	l->25	r->2	v->2	y->6	
amu	s->1	t->1	
amv	e->6	i->3	
amå	l->13	t->22	
amö	t->84	v->2	
an 	"->1	-->6	1->26	4->1	8->2	A->2	B->2	C->2	D->4	E->18	F->2	G->2	H->25	I->13	J->1	K->2	L->1	N->1	P->5	R->1	S->6	V->1	W->3	a->213	b->117	c->3	d->187	e->88	f->208	g->110	h->168	i->246	j->51	k->146	l->63	m->146	n->65	o->249	p->79	r->67	s->249	t->154	u->93	v->177	y->2	Ö->1	ä->103	å->23	ö->23	
an!	 ->224	A->1	D->2	E->2	J->6	M->1	S->1	T->2	U->1	V->2	
an"	 ->2	,->1	.->1	
an,	 ->247	
an-	 ->1	C->1	K->1	
an.	 ->1	(->3	)->1	A->2	D->19	E->2	F->5	H->5	I->4	J->14	K->3	L->1	M->3	N->2	O->1	S->8	T->2	U->3	V->9	
an:	 ->7	
an;	 ->3	
an?	 ->1	F->1	H->2	J->1	O->1	S->1	V->1	Ä->1	
anN	ä->1	
ana	 ->76	,->2	d->6	l->69	m->4	n->2	r->32	s->4	t->5	
anb	e->2	i->9	l->3	o->1	r->2	u->6	
anc	,->1	a->2	e->5	i->1	
and	 ->297	)->1	,->35	.->33	?->1	a->144	e->2524	f->1	i->24	l->360	m->1	n->10	o->14	r->344	s->88	u->3	v->2	z->4	
ane	 ->2	,->1	l->1	n->35	r->108	s->1	t->7	
anf	a->14	l->1	ö->50	
ang	 ->32	,->8	.->12	a->1	e->92	i->5	r->14	å->28	
anh	a->47	e->2	ä->5	å->54	ö->4	
ani	 ->1	,->4	e->9	f->2	k->1	n->35	o->1	s->74	t->2	u->2	v->1	
anj	 ->3	.->1	e->2	o->1	ä->1	
ank	 ->2	"->1	-->1	a->29	e->87	f->9	i->1	l->4	n->1	o->5	r->50	s->2	t->9	
anl	a->1	e->50	i->16	ä->15	ö->4	
anm	a->27	ä->29	
ann	 ->5	,->1	-->1	a->148	e->30	h->1	i->25	l->3	o->13	s->16	ä->2	
ano	 ->4	i->1	n->10	r->13	s->2	
anp	a->14	å->1	
anr	ö->6	
ans	 ->169	,->18	.->5	;->1	?->1	a->10	c->7	d->1	e->250	i->89	j->17	k->252	l->60	m->7	p->116	r->22	t->95	v->317	ä->5	å->13	ö->11	
ant	 ->99	!->1	,->7	.->5	:->1	a->202	e->128	i->81	k->1	l->3	n->1	o->24	r->38	v->2	y->2	ö->3	
anu	a->16	t->1	
anv	a->4	i->1	ä->184	
any	o->3	
anz	 ->3	e->1	
anç	o->1	
anö	s->19	v->1	
ao 	t->1	
aor	d->1	
aos	 ->2	
ap 	-->1	a->22	b->2	d->3	e->1	f->3	g->1	h->1	i->7	k->1	m->2	n->1	o->15	s->11	t->1	u->2	v->1	ä->1	
ap"	 ->1	!->1	,->1	
ap,	 ->16	
ap.	 ->1	D->7	E->1	I->2	J->2	S->1	T->1	V->2	
ap:	 ->1	
apa	 ->100	c->5	d->5	n->28	r->195	s->13	t->10	y->2	
ape	a->1	n->152	r->23	s->1	t->97	
api	t->35	
apk	a->11	
apl	a->1	i->37	
apn	e->2	
apo	l->2	
app	 ->3	,->1	.->1	a->19	e->10	h->3	j->1	l->8	n->1	o->112	s->1	t->5	v->2	y->1	
apr	i->3	o->6	
aps	 ->1	-->1	a->2	b->3	d->1	f->1	i->14	k->3	l->3	m->20	n->11	o->1	p->7	r->18	s->4	å->2	
apt	e->2	
ar 	"->1	(->3	-->13	1->9	2->1	3->1	4->1	9->1	A->2	B->3	C->1	E->15	F->2	G->1	I->1	K->1	L->4	P->3	R->4	S->3	T->1	W->1	a->305	b->134	c->2	d->370	e->244	f->343	g->116	h->125	i->318	j->102	k->131	l->107	m->246	n->118	o->344	p->155	r->93	s->384	t->189	u->120	v->264	y->2	Ö->1	ä->67	å->14	ö->40	
ar!	 ->19	D->1	J->1	M->2	T->1	
ar"	 ->2	
ar)	.->1	
ar,	 ->215	
ar-	 ->1	
ar.	 ->4	)->1	-->1	.->3	A->2	B->4	D->64	E->7	F->16	G->3	H->9	I->14	J->32	K->4	L->3	M->11	N->3	O->9	P->2	R->4	S->7	T->5	U->2	V->30	Ä->2	
ar:	 ->13	
ar;	 ->4	
ar?	I->1	J->1	K->2	N->2	
ara	 ->723	"->1	,->7	.->10	:->2	?->1	b->9	d->23	g->3	k->24	l->5	m->2	n->391	r->94	s->24	t->14	v->4	
arb	a->3	e->564	
arc	e->2	o->1	
ard	 ->9	,->3	-->1	.->1	;->1	a->4	e->24	i->9	
are	 ->602	!->1	"->3	,->77	.->67	:->1	?->3	b->3	f->1	l->3	m->2	n->153	p->1	r->25	s->20	t->72	u->5	
arf	o->1	ä->1	ö->52	
arg	a->8	i->6	o->2	u->17	ö->17	
arh	e->21	u->1	ä->1	å->4	
ari	 ->20	!->1	,->10	.->2	a->3	c->1	e->6	g->62	k->24	n->35	o->4	s->32	t->129	u->2	
arj	e->91	
ark	 ->38	,->4	.->4	a->31	b->1	e->32	i->6	l->1	n->191	o->13	s->2	t->23	
arl	 ->4	-->1	a->606	e->1	i->135	s->2	ä->10	ø->2	
arm	 ->4	-->1	a->16	o->19	r->2	s->3	t->12	y->14	é->3	
arn	 ->8	,->3	a->537	b->1	h->1	i->21	p->2	s->1	
aro	 ->4	,->1	n->3	r->6	u->1	
arp	a->1	e->1	o->1	t->2	
arr	 ->1	a->6	e->2	i->5	o->2	
ars	 ->61	,->4	.->3	a->7	b->3	c->1	e->1	f->55	k->13	l->1	m->3	o->8	p->5	t->11	y->1	
art	 ->203	!->1	,->8	.->16	:->1	a->19	e->64	h->1	i->199	l->1	n->28	o->1	p->1	r->2	s->8	y->69	
arv	 ->1	,->3	.->3	a->9	e->6	i->3	l->1	s->3	ä->1	
ary	 ->1	
arz	w->1	
arä	m->1	
arå	d->2	
aré	b->1	
aró	n->2	
as 	-->2	4->1	E->8	S->2	a->216	b->27	c->5	d->43	e->69	f->116	g->22	h->20	i->144	j->15	k->44	l->22	m->86	n->39	o->106	p->78	r->31	s->109	t->66	u->59	v->49	y->4	ä->13	å->10	ö->14	
as!	D->1	E->1	G->1	H->1	
as"	.->1	
as,	 ->90	
as.	 ->4	-->1	A->2	B->4	C->1	D->31	E->5	F->6	G->3	H->8	I->10	J->10	K->4	M->9	N->3	O->1	P->7	R->1	S->3	T->2	U->1	V->20	Y->1	Ä->1	Å->2	
as:	 ->2	
as;	 ->1	
as?	H->1	S->1	
asa	b->1	c->1	d->2	r->2	s->1	t->2	
asb	o->5	
asc	h->4	i->12	
ase	.->1	b->1	n->9	r->14	
ash	a->1	i->3	u->1	
asi	a->2	e->5	f->1	l->1	n->1	s->31	
ask	 ->1	a->4	e->2	i->12	r->1	u->1	
asm	 ->3	a->1	u->1	
asn	i->3	
aso	c->1	r->1	
asp	e->36	i->1	
ass	 ->6	a->25	e->9	i->23	l->1	m->3	n->4	o->4	p->1	t->1	u->1	
ast	 ->163	!->1	,->5	-->1	.->5	?->1	a->31	e->163	i->17	k->1	l->5	n->8	o->1	r->112	s->72	u->1	ä->1	å->2	
asu	n->1	s->3	
asy	l->21	
asä	k->1	t->19	
aså	 ->4	
at 	"->2	-->11	3->1	9->1	A->1	B->1	E->6	F->2	I->1	K->1	S->1	a->71	b->20	d->42	e->45	f->70	g->12	h->27	i->44	j->2	k->20	l->11	m->36	n->11	o->56	p->30	r->8	s->95	t->26	u->28	v->22	y->1	ä->16	å->5	ö->2	
at,	 ->55	
at.	 ->4	.->1	B->2	D->22	E->3	F->3	G->2	H->8	I->5	J->10	K->4	L->1	M->1	N->1	O->2	P->1	T->3	V->4	Ä->1	Å->1	Ö->1	
at:	 ->3	
at;	 ->1	
at?	.->1	J->1	
ata	 ->24	,->1	b->1	l->10	n->3	r->1	s->90	
atc	h->2	
ate	 ->2	g->71	k->1	l->3	m->2	n->46	r->417	s->1	t->55	
atf	ö->4	
ath	 ->3	,->1	i->2	
ati	 ->18	"->1	,->4	.->9	e->8	f->14	k->5	n->25	o->722	r->1	s->152	v->186	
atj	ä->1	
atl	a->3	i->102	ä->10	
atn	y->1	
ato	 ->10	.->1	a->1	b->2	g->2	l->7	m->8	n->2	r->31	s->13	
atp	e->10	r->1	
atr	i->1	
ats	 ->203	,->28	-->5	.->27	?->2	a->13	b->2	e->104	f->1	k->1	m->4	n->8	o->3	p->1	s->22	
att	 ->6200	,->22	.->26	:->2	?->1	B->1	a->231	e->187	i->36	k->1	l->4	n->82	r->2	s->3	
atu	e->2	l->37	m->14	r->152	s->11	
atz	i->2	
atä	c->1	
atö	r->4	v->6	
atü	r->1	
au 	d->1	f->4	o->1	s->3	
au"	,->1	
au,	 ->7	
au.	E->1	
auM	e->1	
aub	e->1	
auc	t->1	
aud	e->1	r->1	
aue	n->1	r->2	
auf	m->1	
auk	a->3	t->6	
aum	a->1	
aun	a->1	i->3	
aur	e->1	o->1	
aus	 ->3	s->1	u->6	
aut	o->9	r->2	
aux	,->1	
av 	"->3	-->6	1->4	2->1	4->1	5->2	8->1	A->5	B->20	C->1	D->7	E->91	F->12	G->6	H->3	I->2	J->4	K->14	L->5	M->4	O->5	P->4	R->2	S->7	T->8	U->1	V->3	W->3	a->177	b->85	c->9	d->589	e->211	f->223	g->51	h->36	i->41	j->11	k->147	l->54	m->105	n->37	o->69	p->97	r->71	s->210	t->74	u->66	v->97	y->5	Ö->2	ä->8	å->23	ö->15	
av,	 ->11	
av.	(->1	.->1	D->5	E->2	J->1	M->1	O->1	R->1	
av?	V->1	
ava	 ->1	l->5	n->5	r->7	
avb	r->14	
avd	e->8	
ave	 ->4	,->1	-->3	N->1	c->1	n->32	r->13	t->33	u->1	
avf	a->22	o->1	ö->3	
avg	a->2	e->10	i->9	j->4	r->4	å->6	ö->61	
avh	j->2	ä->2	å->1	
avi	 ->1	d->3	e->1	s->9	
avk	l->1	r->1	u->1	
avl	a->9	e->2	i->2	o->1	ä->10	
avm	a->1	
avo	r->1	
avp	r->1	
avr	a->1	e->2	u->1	ä->1	
avs	 ->9	,->4	.->4	?->1	a->7	e->93	f->2	i->39	k->29	l->75	m->2	n->4	o->1	p->5	t->32	v->1	ä->5	
avt	 ->1	a->90	v->1	
avu	n->1	
avv	a->6	e->10	i->23	ä->3	
aw,	 ->1	
aw.	M->1	
ax 	a->1	e->1	i->1	
ax-	f->3	
axa	 ->2	
axb	e->1	
axe	l->1	r->1	
axi	m->9	s->8	
axl	a->1	
ay 	f->2	h->1	
ay,	 ->4	
ay.	V->1	
ayD	e->1	
aya	b->3	g->4	n->2	
ayb	e->1	
aye	d->2	r->1	
ays	 ->3	-->1	
aza	 ->1	,->1	.->2	k->1	r->2	
azi	s->16	
aça	 ->5	
b S	ö->2	
b e	f->1	
b h	a->1	j->1	
b k	a->1	
b o	c->3	
b s	k->1	
b v	a->1	
b) 	i->1	m->1	
b, 	e->1	s->2	v->1	
b-o	m->1	
b.A	n->1	
b.D	e->1	
ba 	a->1	b->2	f->1	o->2	p->1	r->1	t->1	u->1	v->1	å->1	
ba-	,->1	
bac	i->1	k->2	è->1	
bad	 ->4	a->1	e->27	s->1	
bag	a->2	
bai	n->1	
bak	 ->1	,->1	a->51	d->1	g->31	o->21	s->2	t->1	å->3	
bal	 ->1	a->39	i->5	l->1	t->2	
ban	 ->1	"->1	a->6	b->1	d->53	e->6	i->2	k->20	n->1	o->8	s->4	t->2	
bar	 ->42	,->1	.->4	a->287	b->2	d->1	e->11	g->1	h->9	i->2	k->1	l->12	m->1	n->13	r->2	t->98	é->1	
bas	 ->10	,->1	.->1	a->2	e->14	i->4	k->5	s->1	t->6	u->1	
bat	 ->3	s->9	t->172	
bax	a->1	
bay	e->1	
bb 	e->1	h->1	o->3	v->1	
bb,	 ->2	
bba	 ->12	d->27	r->15	s->11	t->12	
bbe	l->7	
bbi	g->1	
bbl	a->11	
bbp	l->1	
bbt	 ->34	,->3	.->6	
bbv	a->1	
bby	,->1	a->1	b->1	g->2	i->2	m->1	n->3	v->1	
be 	P->1	e->5	f->1	h->2	k->6	o->2	p->1	s->1	
bea	k->30	r->2	
beb	o->1	y->1	å->1	
bed	d->1	r->51	s->1	ö->51	
bef	a->11	i->41	l->1	o->82	r->20	ä->12	
beg	a->4	r->105	ä->60	å->11	
beh	a->87	o->67	ä->1	å->29	ö->166	
bei	v->1	
bek	a->3	i->2	l->42	o->2	r->30	v->15	y->16	ä->42	
bel	 ->9	!->1	,->4	.->5	a->14	g->8	l->6	o->16	s->3	t->29	v->1	y->4	ä->7	ö->2	
bem	a->2	y->1	ä->5	ö->10	
ben	 ->1	e->6	g->1	h->1	i->3	s->1	ä->1	å->1	
beo	r->1	
ber	 ->81	,->13	.->6	a->32	b->1	e->65	g->4	i->9	n->2	o->94	t->2	v->1	y->1	ä->35	ö->45	
bes	 ->2	e->2	i->4	k->35	l->222	p->5	t->226	v->32	y->1	ä->3	ö->11	
bet	 ->12	"->2	,->3	-->1	.->2	?->1	a->233	e->228	h->1	j->1	o->46	r->96	s->224	t->5	u->1	v->3	y->122	ä->268	
beu	n->3	
bev	a->28	e->1	i->92	
bex	p->1	
bi 	d->1	n->1	
bib	e->11	l->2	
bid	r->111	
bie	f->2	
bif	a->5	
big	a->1	o->1	å->6	
bih	a->1	
bik	m->2	
bil	 ->12	,->2	-->1	.->3	a->95	b->2	d->108	e->7	i->67	j->1	k->4	l->6	m->1	p->7	s->7	t->17	v->6	ä->1	å->1	
bin	,->1	a->1	d->37	e->3	
bio	 ->1	g->1	l->4	p->1	s->3	
bis	e->2	k->12	t->23	
bit	 ->1	e->1	i->26	t->3	
bje	k->2	
bju	d->42	
bjö	d->2	
bl.	a->27	
bla	 ->22	"->1	,->1	.->4	d->1	m->1	n->102	r->2	s->1	
ble	k->1	m->184	r->15	s->1	v->15	
bli	 ->129	,->1	.->1	c->30	g->14	k->20	n->9	o->2	r->115	v->27	x->1	
blo	c->6	m->6	n->1	t->3	
blu	n->4	
bly	 ->1	,->2	.->1	g->4	
blå	 ->1	s->2	
bni	n->1	
bo 	i->1	k->1	v->1	
boa	r->1	
boc	k->2	
bod	a->3	
boe	l->1	n->3	
bog	s->1	
boj	k->1	
bok	 ->16	,->1	.->5	e->36	s->2	
bol	 ->2	a->12	i->7	l->1	
bom	b->9	u->1	
bon	 ->4	,->1	.->1	d->2	m->2	
bor	 ->6	a->3	d->79	g->174	r->1	t->47	
bos	a->3	n->2	t->5	ä->4	
bot	 ->2	a->2	t->9	
bou	r->5	
bov	a->1	e->1	
box	n->1	
bpl	a->1	
bra	 ->64	!->1	,->8	.->6	n->10	
bre	d->17	i->1	p->1	t->7	v->6	
bri	e->4	g->1	k->3	n->13	s->62	t->31	
bro	 ->2	a->1	d->2	k->2	m->10	n->1	r->1	t->55	
bru	a->16	k->80	n->1	t->6	
bry	g->3	o->1	r->2	t->18	
brä	n->15	s->2	
brå	d->20	k->1	s->2	
brö	d->3	s->1	t->7	
bse	r->2	
bsi	d->23	
bso	l->40	r->1	
bst	a->6	r->1	
bsu	r->3	
bt 	f->5	g->2	h->1	k->3	l->1	m->2	o->1	p->1	s->14	t->1	u->1	v->2	
bt,	 ->3	
bt.	J->1	M->1	O->2	T->1	V->1	
bu 	i->1	
bud	 ->22	,->4	.->3	d->1	e->9	g->106	o->1	s->27	
bug	g->1	
buk	t->2	
bul	 ->1	a->2	t->1	
bun	d->28	
bur	e->1	g->11	i->1	n->1	
bus	 ->1	s->2	
but	i->2	
bva	r->1	
bve	n->12	
bvä	r->1	
by,	 ->1	
bya	r->1	
byb	i->1	
bye	n->1	
byg	d->45	g->100	r->2	
byi	s->2	
bym	a->1	
byn	 ->3	
byr	å->35	
byt	a->2	e->17	t->1	
byv	e->1	
byx	f->1	
bäl	t->10	
bän	k->1	
bär	 ->106	,->1	.->2	a->30	l->4	s->2	
bäs	t->42	
bät	t->153	
bäv	n->10	
båd	a->26	e->46	
båt	a->8	e->1	
bé 	a->1	
béb	é->1	
böc	k->3	
böd	e->1	
böj	e->1	t->1	
böl	d->1	
bör	 ->208	,->1	.->1	a->1	d->26	j->115	l->10	s->2	
böt	e->1	
c -	 ->1	
c B	r->1	
c b	l->1	ö->1	
c d	å->1	
c i	 ->2	
c l	'->1	
c o	s->1	
c s	e->1	
c",	 ->1	
c) 	l->1	
c, 	d->1	
c-d	i->1	
c-s	y->1	
c-t	r->1	
c. 	o->1	Ä->2	
c.D	e->1	
c.E	n->1	
c?A	t->1	
cCa	r->1	
cNa	l->5	
ca 	3->1	C->1	M->3	s->1	
ca,	 ->1	
ca.	 ->1	
cal	 ->1	v->1	
can	c->2	n->1	t->1	
cao	 ->1	
cap	 ->1	i->10	
cas	 ->1	e->1	
cay	a->6	
cce	p->89	s->5	
ce 	b->1	d->4	f->1	n->1	o->12	t->2	
ce,	 ->1	
ce.	.->1	A->1	D->1	J->2	O->1	S->1	
ced	o->1	u->1	
cek	o->1	v->1	
cel	o->2	
cem	b->19	e->2	i->1	
cen	 ->1	,->1	a->5	e->1	n->7	s->2	t->226	
cep	t->102	
cer	!->1	,->1	a->75	b->1	i->13	n->2	t->6	
ces	s->114	
ceu	t->1	
ch 	"->3	(->1	-->6	0->1	1->21	2->13	3->7	4->10	5->3	6->2	7->6	8->11	9->4	A->4	B->6	C->4	D->4	E->36	F->15	G->7	H->3	I->14	J->2	K->9	L->8	M->5	N->2	O->2	P->15	R->3	S->26	T->8	U->1	V->2	W->1	X->1	a->292	b->119	c->10	d->609	e->212	f->321	g->92	h->162	i->234	j->162	k->198	l->93	m->279	n->84	o->98	p->115	r->188	s->448	t->153	u->106	v->237	y->7	Ö->7	ä->55	å->37	ö->43	
ch!	 ->1	
ch)	D->1	
ch,	 ->14	
ch.	E->1	J->1	
ch/	e->1	
ch:	 ->1	
ch?	F->1	
chI	 ->1	I->1	
cha	b->1	n->13	p->1	r->4	
che	 ->1	c->1	f->17	m->1	n->16	r->6	z->1	
chh	o->1	
chi	e->1	s->1	
chl	e->4	
chn	e->12	
cho	c->4	k->1	
chr	e->3	o->14	ö->1	
chs	 ->1	
cht	 ->2	.->1	e->2	f->3	i->1	
chu	l->3	
chw	a->1	e->1	i->1	
chy	r->1	
chö	r->1	
chü	s->4	
cia	l->220	
cid	e->1	
cie	l->49	n->4	r->1	t->1	
cif	i->29	
cil	 ->1	l->1	o->1	
cin	e->1	
cio	 ->8	,->3	.->2	:->1	e->3	s->2	
cip	 ->28	,->3	.->4	e->151	i->8	l->14	s->1	
cir	k->10	
cis	 ->39	-->1	a->1	e->11	m->3	t->11	
cit	.->1	a->9	e->14	
civ	i->19	
ck 	-->1	K->1	a->21	b->3	d->6	e->9	f->29	g->4	h->7	i->17	j->5	k->8	l->2	m->10	n->6	o->12	p->3	s->29	t->17	u->2	v->17	ä->2	å->2	
ck"	 ->1	
ck,	 ->28	
ck-	p->1	
ck.	 ->1	A->1	D->2	F->1	H->2	J->2	K->2	Ä->1	
cka	 ->157	"->1	,->5	.->2	?->1	d->19	n->45	r->25	s->28	t->25	
ckb	a->5	i->1	ä->1	
ckd	e->8	
cke	 ->22	-->19	.->3	l->8	n->21	r->115	t->476	
ckf	r->1	ö->7	
ckh	e->15	o->3	
cki	t->1	
ckl	a->78	e->4	i->281	
ckn	a->29	e->1	i->47	
cko	r->39	s->1	
ckp	r->3	
ckr	a->6	
cks	 ->21	.->2	;->1	a->9	b->1	c->1	d->3	f->2	i->3	k->1	o->2	r->2	v->1	å->587	ö->1	
ckt	 ->13	e->22	s->4	
cku	p->5	
ckv	i->3	
ckö	n->5	
cli	n->1	
co,	 ->1	
co-	a->1	
cob	 ->2	
com	b->1	m->1	p->1	
con	d->1	t->2	
cop	y->1	
cor	e->1	p->4	r->1	
cos	t->5	
cou	p->1	r->1	
cov	e->1	
cqu	e->3	i->1	
cri	c->1	
ct.	 ->1	
ctn	e->1	
cto	r->2	
cu 	m->1	
cu,	 ->1	
cy,	 ->1	
cya	v->1	
cyc	l->1	
cyd	e->1	
cyf	ö->1	
cyk	e->3	l->4	
cèt	e->1	
d "	a->2	e->1	
d (	a->2	e->1	k->1	r->1	
d -	 ->11	
d 1	2->2	3->2	4->1	6->1	9->1	
d 2	 ->3	0->2	4->1	7->2	8->1	
d 3	0->1	6->1	
d 5	 ->1	
d 7	 ->1	0->1	
d 8	0->2	
d A	.->1	d->1	m->2	
d B	N->1	S->1	a->3	y->3	
d C	o->1	
d D	a->2	
d E	-->1	D->1	G->3	U->3	r->4	u->17	
d F	P->1	r->4	
d G	A->1	e->1	u->1	
d H	a->5	
d I	n->3	s->2	
d J	ö->1	
d K	o->3	u->2	y->1	
d L	T->1	a->4	e->1	i->2	
d M	a->3	e->1	i->1	
d O	L->1	s->1	
d P	a->2	
d R	y->1	
d S	a->1	v->1	y->5	
d T	h->1	i->1	u->2	
d U	S->4	
d V	a->1	e->1	
d W	i->1	
d a	)->1	c->1	d->2	l->42	n->72	r->15	t->188	u->2	v->159	
d b	a->6	e->59	i->10	l->5	o->2	r->10	u->1	y->2	ä->1	å->2	ö->7	
d c	a->1	i->1	
d d	a->9	e->341	i->8	o->5	r->3	u->2	y->2	ä->9	å->4	
d e	f->11	k->2	l->13	n->118	r->16	t->42	u->5	v->1	x->5	
d f	a->8	e->2	i->7	l->10	o->7	r->64	u->11	y->2	ä->1	å->4	ö->176	
d g	a->2	e->15	i->2	j->2	l->2	o->7	r->10	ä->60	ö->2	
d h	a->40	e->4	i->1	j->26	o->4	u->5	ä->23	å->1	ö->6	
d i	 ->90	b->1	d->3	f->1	m->2	n->65	s->2	v->2	
d j	a->15	o->3	u->3	ä->3	
d k	a->22	i->1	l->3	n->1	o->75	r->11	u->5	v->13	ä->3	ö->1	
d l	a->5	e->4	i->9	u->1	ä->5	ö->4	
d m	a->26	e->100	i->42	o->18	y->9	ä->1	å->19	ö->7	
d n	a->18	e->3	i->5	o->1	u->4	y->7	ä->10	å->11	ö->8	
d o	c->107	e->1	f->2	j->1	l->5	m->81	p->1	r->8	s->14	t->1	
d p	a->18	e->8	l->3	o->8	r->17	s->1	u->6	å->50	
d r	a->1	e->32	i->3	o->3	ä->16	å->7	ö->2	
d s	.->1	a->19	e->11	i->39	j->5	k->25	l->4	m->4	n->2	o->145	p->5	t->54	u->3	v->2	y->12	ä->20	å->16	
d t	.->2	a->60	e->4	i->112	j->1	o->4	r->13	u->2	v->8	y->1	ä->4	
d u	n->13	p->15	r->3	t->38	
d v	a->28	e->15	i->68	o->1	ä->2	å->22	
d y	r->3	t->5	
d Ö	V->1	s->1	
d ä	n->13	r->48	v->2	
d å	r->4	t->13	
d ö	k->2	m->1	p->2	s->1	v->33	
d! 	L->1	N->1	
d) 	i->1	
d),	 ->3	
d, 	"->1	5->1	D->1	E->1	F->1	I->2	N->1	S->2	a->6	b->3	d->13	e->9	f->7	g->1	h->9	i->4	k->3	l->1	m->20	n->3	o->29	p->3	r->2	s->22	t->5	u->4	v->9	ä->3	
d- 	(->1	
d-a	f->1	
d-f	ö->1	
d-k	o->1	
d. 	V->1	Ö->1	ö->1	
d."	J->1	M->1	
d.(	S->1	
d.,	 ->1	
d.-	 ->1	
d..	 ->1	(->1	
d.A	l->1	n->1	t->2	
d.B	e->1	
d.D	e->49	i->2	ä->3	å->1	
d.E	f->1	m->1	n->1	u->3	
d.F	a->1	r->2	ö->5	
d.G	e->1	
d.H	a->2	e->13	u->1	
d.I	 ->6	n->3	r->1	
d.J	a->23	
d.K	a->1	o->6	
d.L	å->2	
d.M	a->1	e->8	i->1	o->1	ä->1	å->1	
d.N	a->1	i->2	u->2	ä->2	
d.O	m->17	r->1	
d.P	a->1	å->1	
d.R	e->3	
d.S	a->1	o->2	u->1	å->1	
d.T	a->1	i->1	r->1	
d.U	n->1	p->1	t->2	
d.V	a->2	e->1	i->13	
d.Ä	n->1	v->1	
d.Å	 ->2	r->1	
d: 	"->2	d->1	e->1	
d; 	d->3	i->2	
d? 	H->1	
d?-	 ->2	
d?.	 ->1	
d?D	ä->1	
d?F	ö->1	
d?H	e->1	
d?J	a->1	
d?V	i->1	
d?Ä	r->1	
da 	-->1	1->1	2->1	6->1	C->5	E->6	F->1	G->1	a->59	b->14	c->3	d->60	e->41	f->60	g->9	h->12	i->39	j->4	k->22	l->14	m->45	n->12	o->31	p->35	r->28	s->73	t->52	u->16	v->18	ä->7	å->8	ö->4	
da!	D->1	
da"	 ->1	
da,	 ->39	
da.	 ->1	B->1	D->6	E->1	F->3	H->5	I->2	J->3	K->1	M->3	N->2	O->2	R->1	V->5	Ä->2	
da?	D->2	F->1	I->1	
dab	o->2	
dac	 ->3	"->1	-->1	
dad	 ->8	.->1	e->31	
daf	o->1	r->2	
dag	 ->165	,->32	.->33	:->2	a->18	e->36	l->8	o->53	s->25	
dah	å->43	
dai	r->1	
dak	i->3	t->3	
dal	!->1	,->1	a->5	e->5	y->2	ö->1	
dam	 ->10	,->3	.->1	a->1	e->46	f->27	m->4	o->74	r->1	å->13	ö->84	
dan	 ->404	,->17	.->18	?->3	a->53	b->2	d->106	f->1	g->1	h->1	i->1	m->1	o->1	r->6	s->33	t->93	
dap	e->1	
dar	 ->38	,->2	.->2	b->2	d->24	e->120	f->1	i->31	n->23	s->4	
das	 ->38	,->5	.->14	?->1	t->86	
dat	 ->24	,->4	.->2	a->4	e->11	i->33	l->12	o->3	p->9	s->8	u->13	
dba	r->9	
dbe	d->1	l->1	s->17	t->1	
dbo	r->170	
dbr	o->1	u->56	ä->1	
dbu	l->1	
dbä	v->10	
dd 	a->22	b->2	e->1	f->18	h->1	i->2	m->5	o->4	s->4	t->3	u->2	v->2	ä->2	ö->1	
dd)	,->1	
dd,	 ->4	
dd.	D->2	J->2	M->1	N->1	R->1	V->1	
dda	 ->58	.->2	d->6	g->13	n->1	r->3	s->2	t->1	
dde	 ->37	,->1	l->63	n->3	r->1	s->11	t->18	
ddh	i->1	
ddi	g->2	n->2	t->1	
ddn	i->4	
dds	 ->1	m->4	n->6	o->2	p->1	s->2	t->1	
de 	"->9	(->30	-->20	1->10	2->6	4->2	8->1	9->1	A->5	B->2	C->2	D->2	E->8	F->1	G->5	H->3	I->2	J->1	K->6	L->2	M->5	N->2	O->2	P->20	R->3	S->6	T->2	V->2	W->1	a->376	b->163	c->4	d->169	e->199	f->423	g->94	h->130	i->274	j->27	k->229	l->70	m->272	n->137	o->326	p->228	r->192	s->447	t->182	u->102	v->163	y->14	Ö->1	ä->76	å->78	ö->46	
de!	 ->6	A->1	J->1	N->1	
de"	,->1	
de(	A->1	
de,	 ->172	
de-	 ->1	F->2	L->1	l->1	
de.	 ->6	-->1	.->1	A->4	D->43	E->9	F->10	G->2	H->15	I->6	J->35	K->4	L->4	M->18	N->4	O->6	P->4	R->1	S->12	T->10	U->2	V->13	Å->1	
de:	 ->39	
de;	 ->5	
de?	D->1	F->1	H->3	J->1	V->1	
deH	e->1	
deP	r->1	
dea	d->1	l->5	u->1	
deb	a->170	e->1	u->9	ä->1	
dec	e->41	
ded	e->2	
dee	l->2	r->2	
def	i->36	o->1	r->1	u->7	ö->13	
deg	e->4	r->1	
deh	ö->1	
dei	r->2	
dek	o->9	r->1	v->5	
del	 ->201	,->23	.->20	?->1	a->187	b->19	e->79	f->1	g->1	h->4	l->17	n->43	p->2	r->1	s->286	t->60	u->2	v->11	ö->1	
dem	 ->143	,->11	.->32	:->2	?->1	a->6	e->5	i->3	o->153	
den	 ->2311	"->1	)->5	,->121	.->169	:->7	;->4	?->6	N->1	a->83	b->2	i->2	n->527	s->73	t->57	
deo	l->5	
dep	a->9	
der	 ->1049	"->1	)->7	,->69	-->1	.->92	:->1	;->1	?->3	a->178	b->14	d->6	e->3	g->5	h->5	i->62	k->5	l->59	m->6	n->294	o->4	r->3	s->124	t->19	u->3	v->2	ä->3	ö->1	
des	 ->208	,->8	.->9	a->2	b->1	d->2	g->1	k->115	p->7	s->487	t->5	v->2	
det	 ->3568	!->2	)->2	,->119	.->154	:->3	;->1	?->9	a->35	s->121	t->829	
deu	r->2	t->1	
dev	a->6	i->2	
dez	,->1	-->2	
dfi	l->1	n->2	
dfr	å->10	
dfu	l->1	
dfä	l->4	
dfö	d->1	r->248	
dga	 ->28	,->1	?->1	d->6	n->10	r->5	s->13	t->3	
dge	 ->4	r->10	s->5	t->108	
dgi	v->28	
dgn	i->71	
dgo	r->1	
dgr	ä->1	ö->1	
dgä	n->2	
dgå	n->2	r->2	t->1	
dgö	r->3	
dhe	t->25	
dhi	s->1	
dhj	ä->1	
dhå	l->4	
dhö	l->1	
di 	-->1	a->3	b->1	h->2	i->1	l->2	o->5	r->1	s->2	t->2	
di,	 ->1	
di.	D->1	S->1	V->1	
di:	 ->1	
di;	 ->1	
dia	 ->5	l->32	r->21	s->1	t->1	
dic	a->1	e->1	i->1	
did	a->14	
die	 ->3	,->1	b->1	k->1	n->7	p->1	r->14	t->4	
dif	f->5	i->5	
dig	 ->46	,->2	.->5	a->157	e->2	h->250	n->1	r->2	s->1	t->235	
dik	a->29	e->1	t->10	
dil	e->3	
dim	e->13	
din	a->1	b->1	f->1	g->11	s->3	ä->1	
dio	l->2	x->7	
dip	l->11	
dir	e->248	i->1	l->2	
dis	 ->8	c->14	e->9	k->213	p->4	t->4	
dit	 ->13	a->1	e->2	h->1	i->22	s->1	
diu	m->4	
div	e->4	i->14	
diz	 ->3	,->1	-->1	
diä	r->1	
dja	 ->69	.->2	n->6	r->6	s->8	
dje	 ->63	,->4	:->1	d->6	k->2	l->6	r->1	
djo	r->1	
dju	n->2	p->39	r->17	
djä	r->7	v->2	
dka	r->1	
dko	m->24	r->1	
dku	r->1	s->2	
dkv	i->1	
dkä	n->94	
dla	 ->23	.->2	d->11	g->2	n->1	r->122	s->14	t->7	
dle	m->343	n->12	t->1	
dli	d->2	g->199	n->193	s->1	
dlä	g->79	
dlö	s->1	
dma	k->1	
dme	d->4	
dmi	n->25	u->3	
dmo	n->3	t->1	
dmä	n->1	
dmå	l->2	n->1	
dna	 ->13	c->2	d->10	n->2	p->1	r->5	s->2	t->3	
dni	n->407	v->1	
do 	R->1	a->4	
do,	 ->1	
do.	D->1	F->1	H->1	O->1	
doc	k->61	
doe	f->1	
dof	i->1	
dog	 ->1	.->2	j->1	m->2	ö->9	
dok	u->45	
dol	f->2	l->9	
dom	 ->18	,->5	.->1	/->1	a->28	e->10	i->8	l->3	r->14	s->98	
don	 ->33	,->10	.->10	?->1	N->1	e->7	s->7	t->1	
dor	 ->16	,->4	.->4	d->1	e->2	n->11	s->1	
dos	a->1	e->1	k->3	t->2	
dou	 ->1	
dov	i->4	
dox	,->1	a->5	
doä	m->1	
dpe	l->1	
dpo	l->1	
dpr	i->1	
dpu	n->119	
dra	 ->434	,->23	.->7	:->4	;->2	b->55	d->25	g->417	h->1	k->1	m->8	n->14	r->70	s->33	t->27	
dre	 ->59	,->2	.->2	?->1	k->1	n->3	s->2	t->1	v->1	
dri	a->2	c->3	d->3	f->8	g->32	k->3	n->315	v->54	
dro	g->10	l->2	m->1	n->1	p->1	t->4	
dru	c->2	n->3	s->1	
dry	f->1	g->3	
drä	g->37	n->3	
drå	p->1	
drö	j->8	m->1	
ds 	a->9	b->7	d->3	e->3	f->5	g->2	i->9	j->1	l->2	m->6	n->1	o->3	p->26	r->4	s->7	t->3	u->2	v->2	ä->1	å->4	ö->2	
ds,	 ->4	
ds-	 ->2	i->2	n->1	s->1	
ds.	 ->1	B->1	D->1	J->1	U->1	
ds/	i->1	
ds;	 ->1	
dsN	ä->1	
dsa	k->17	m->7	n->5	r->5	t->1	v->6	
dsb	e->12	u->1	y->43	
dsc	e->1	
dsd	e->13	i->3	o->1	u->1	ö->1	
dse	f->4	k->15	n->2	t->2	
dsf	a->1	r->15	ö->8	
dsg	r->1	
dsh	a->6	
dsi	n->8	t->1	
dsj	u->1	
dsk	 ->5	-->1	a->65	o->6	r->8	t->1	ä->3	
dsl	a->12	i->3	ä->2	å->1	ö->2	
dsm	a->11	e->11	i->1	y->2	ä->5	å->1	ö->2	
dsn	i->8	
dso	m->8	r->23	
dsp	a->5	e->10	l->11	o->3	r->34	u->1	
dsr	a->5	e->7	y->2	ä->1	ö->1	
dss	a->4	k->2	t->30	y->2	ä->1	
dst	a->4	e->1	i->1	j->2	o->4	r->1	u->2	ä->5	
dsu	p->2	t->3	
dsv	e->1	i->3	ä->1	
dsy	f->1	s->4	
dsä	n->1	
dså	l->2	t->1	
dsö	d->1	
dt 	f->1	h->1	o->3	s->1	t->1	u->1	
dt,	 ->4	
dta	 ->44	.->1	b->6	g->24	l->1	r->11	s->21	
dte	r->14	s->1	
dti	d->1	
dto	g->4	
dty	c->6	s->1	
du 	b->2	c->1	m->1	ä->2	
dua	l->1	
dub	b->17	
duc	e->35	
due	l->7	r->1	
dug	a->1	l->6	
duk	a->1	t->54	
dum	h->3	p->4	t->1	
dun	a->1	k->1	
dup	p->4	
dur	r->1	
dus	s->1	t->114	
dut	s->1	y->1	
dva	g->1	l->24	t->1	
dve	r->19	t->42	
dvi	k->39	n->2	s->3	
dvo	k->5	
dvr	i->12	ä->1	
dvs	.->45	
dvu	n->1	
dvä	n->126	r->1	s->2	
dwi	l->1	
dyk	a->2	e->5	
dyl	i->3	
dyn	a->5	
dyr	 ->1	a->4	k->1	t->2	
dys	t->1	
dzi	o->4	
dzj	i->5	
däc	k->1	
däm	p->2	
där	 ->214	!->1	,->10	.->14	?->1	a->2	e->20	f->184	h->1	i->24	m->40	p->2	r->1	t->1	v->8	
då 	2->1	A->1	D->1	E->3	a->19	b->16	d->17	e->6	f->14	g->4	h->7	i->16	j->3	k->15	l->1	m->9	o->11	p->4	r->4	s->16	t->12	u->5	v->14	ä->4	ö->1	
då,	 ->3	
då.	.->1	D->1	
då?	I->1	
dål	i->19	
dåt	g->6	
dåv	a->1	
dé 	-->1	a->2	j->1	k->1	o->1	s->3	ä->1	
dé,	 ->1	
dée	,->1	r->8	
dén	 ->14	,->1	
dö 	i->1	
död	 ->5	.->3	a->10	f->1	s->2	
döe	n->1	
döl	j->10	
döm	a->37	b->1	d->3	e->11	l->2	n->28	s->3	t->5	
döp	a->1	e->2	t->1	
dör	 ->5	r->9	
dös	t->1	
döt	t->3	
döv	t->1	
e "	a->2	d->1	f->1	k->2	l->2	s->1	
e (	A->29	B->1	C->2	K->2	a->1	f->1	m->1	
e -	 ->42	,->1	
e 1	0->1	1->2	2->1	4->4	5->3	8->1	9->5	
e 2	0->2	1->1	5->4	6->1	
e 3	5->1	
e 4	,->1	0->1	1->1	
e 8	 ->1	
e 9	 ->1	
e A	h->1	l->2	m->3	
e B	 ->1	N->1	a->2	e->2	u->1	
e C	e->2	u->1	
e D	a->1	e->1	i->1	u->1	
e E	M->1	U->4	k->1	u->23	
e F	N->1	o->2	r->2	u->1	
e G	a->3	r->4	
e H	a->1	e->1	i->1	o->1	
e I	m->1	r->1	s->1	t->1	
e J	a->1	o->1	
e K	a->2	i->3	o->3	
e L	a->1	o->1	
e M	a->4	e->1	
e N	a->2	
e O	L->1	i->1	u->1	
e P	a->7	l->1	r->15	
e Q	u->1	
e R	a->1	e->1	o->4	
e S	a->1	c->2	e->1	v->1	w->1	
e T	r->1	u->1	
e V	a->1	e->1	
e W	e->1	
e a	b->2	c->11	d->7	f->1	g->4	i->1	k->10	l->81	m->5	n->124	p->2	r->29	s->5	t->241	u->4	v->232	
e b	a->110	e->188	i->30	l->49	o->7	r->19	u->4	y->11	ä->9	å->11	é->1	ö->18	
e c	e->4	h->4	i->1	o->2	
e d	a->26	e->297	i->26	j->1	o->15	r->17	u->1	y->2	ä->36	å->12	ö->3	
e e	f->15	g->6	j->1	k->27	l->24	m->5	n->141	p->2	r->23	t->52	u->65	v->3	x->28	
e f	a->70	e->13	i->57	j->4	l->35	o->35	r->173	u->14	y->11	ä->2	å->58	ö->406	
e g	a->20	e->69	i->3	j->8	l->11	o->22	r->55	ä->16	å->32	ö->42	
e h	a->247	e->67	i->13	j->6	o->15	u->11	y->2	ä->30	å->12	ö->17	
e i	 ->237	a->2	c->8	d->4	f->4	g->2	l->1	m->1	n->242	s->4	t->6	
e j	a->73	e->1	o->7	u->9	ä->4	
e k	a->132	e->1	i->5	l->10	n->3	o->231	r->36	u->116	v->11	ä->11	ö->1	
e l	a->54	e->29	i->20	o->11	u->1	y->10	ä->64	å->13	ö->10	
e m	a->130	e->215	i->67	o->20	u->4	y->30	ä->38	å->89	ö->14	
e n	a->56	e->5	i->18	o->19	u->21	y->32	ä->46	å->42	ö->15	
e o	a->1	b->4	c->282	e->1	f->16	l->58	m->173	n->2	p->4	r->44	s->14	t->1	v->5	
e p	a->42	e->51	i->1	l->10	o->44	r->90	u->16	å->193	
e q	u->2	
e r	a->23	e->160	i->29	o->11	u->5	y->1	ä->63	å->23	ö->6	
e s	a->51	e->88	i->51	j->13	k->139	l->11	m->22	n->12	o->229	p->11	t->148	u->5	v->17	y->37	ä->72	å->32	ö->5	
e t	.->2	a->89	e->12	i->259	j->13	o->10	r->32	u->8	v->32	y->12	ä->9	
e u	l->1	n->38	p->80	r->9	t->145	
e v	a->168	e->53	i->263	o->8	r->1	ä->37	å->8	
e y	r->3	t->11	
e Ö	s->1	
e ä	g->4	l->1	m->1	n->86	r->163	v->9	
e å	 ->1	k->1	l->1	r->52	s->5	t->76	
e ö	a->1	k->7	m->1	n->11	p->11	s->3	v->65	
e! 	J->5	N->2	
e!A	l->1	
e!D	e->1	
e!J	a->1	
e!M	e->1	
e!N	i->1	
e!S	k->1	
e!Ä	v->1	
e" 	s->2	
e",	 ->3	
e(A	5->1	
e) 	f->1	i->1	o->1	
e, 	,->1	A->1	B->1	D->3	E->2	F->2	G->1	H->1	L->2	R->1	S->1	a->20	b->13	d->24	e->13	f->15	g->3	h->21	i->24	j->4	k->14	l->3	m->30	n->15	o->48	p->10	r->1	s->33	t->9	u->8	v->30	ä->11	å->4	ö->1	
e- 	o->6	p->1	
e-A	l->1	r->1	t->1	
e-F	r->2	
e-L	e->1	o->1	
e-M	a->1	
e-N	o->1	
e-a	l->1	v->3	
e-d	a->1	e->2	i->2	
e-f	a->1	o->1	ö->1	
e-l	o->1	ä->1	
e-m	a->1	e->1	
e-p	r->2	
e-s	p->3	t->11	
e. 	D->6	M->1	O->2	V->2	Ä->1	
e.-	 ->2	
e..	 ->3	(->1	.->1	
e.A	k->1	l->2	n->1	t->2	v->3	
e.B	e->2	å->1	
e.D	e->83	ä->8	å->2	
e.E	f->5	m->1	n->8	t->1	u->4	
e.F	P->1	r->5	ö->15	
e.G	e->2	r->1	
e.H	a->2	e->13	o->1	u->5	
e.I	 ->9	d->1	m->1	n->2	
e.J	a->60	
e.K	a->2	o->7	
e.L	i->2	y->1	ä->1	å->4	
e.M	a->8	e->19	i->7	å->1	
e.N	i->4	u->2	ä->3	
e.O	c->3	f->1	m->7	
e.P	a->1	l->1	o->1	r->2	å->2	
e.R	e->2	o->1	å->2	
e.S	a->2	c->1	e->1	k->1	l->2	o->8	t->2	å->3	
e.T	V->1	a->4	i->3	o->1	r->3	v->1	
e.U	n->2	p->1	r->1	
e.V	a->6	i->27	å->3	
e.d	.->1	
e.Ä	n->2	r->1	v->2	
e.Å	 ->1	r->1	t->2	
e.Ö	s->1	
e: 	"->2	A->3	D->2	F->3	G->3	H->1	I->1	J->2	K->3	M->1	N->3	P->1	S->2	T->1	U->1	V->4	b->2	d->1	f->1	h->1	i->2	k->1	t->1	u->1	v->1	Å->2	
e; 	d->2	h->1	j->1	m->1	p->1	
e?D	e->2	
e?E	n->1	
e?F	ö->2	
e?H	e->4	u->1	ä->1	
e?I	 ->1	
e?J	a->1	
e?K	a->1	
e?O	c->1	
e?S	o->1	
e?V	i->2	
eEn	 ->1	
eFr	u->1	
eHe	r->1	
eNä	s->2	
ePr	o->1	
ea 	b->1	o->3	
ead	-->1	e->5	i->1	l->1	
eag	e->16	
eak	e->1	t->53	
eal	 ->1	,->2	a->1	e->2	i->17	
eam	i->8	
ean	-->1	u->1	
ear	b->3	v->1	
eat	e->1	i->2	o->22	t->4	ö->1	
eau	 ->2	"->1	,->2	x->1	
eb,	 ->1	
eba	l->1	n->1	r->1	s->2	t->170	
ebb	e->1	p->1	
ebe	f->3	h->1	n->1	s->4	t->12	
ebi	l->1	
ebo	a->1	e->2	l->4	r->1	
ebr	e->1	o->1	u->16	å->2	ö->1	
ebu	d->9	
eby	g->25	
ebä	l->10	n->1	r->108	
ebå	d->1	
ebö	r->8	
ec 	l->1	
ece	d->1	m->19	n->22	
eci	a->14	e->42	f->29	r->1	s->49	
eck	 ->3	a->24	e->15	l->248	n->32	o->17	
eco	v->1	
ect	n->1	
ecu	 ->1	,->1	
ecy	c->1	
ed 	"->3	(->1	-->1	1->6	2->8	3->2	5->1	8->1	A->3	B->2	D->2	E->19	F->4	G->1	H->4	I->3	J->1	K->2	L->3	M->4	O->2	P->1	R->1	S->5	T->3	U->4	V->2	a->200	b->24	d->264	e->142	f->91	g->20	h->58	i->54	j->3	k->58	l->16	m->73	n->39	o->59	p->52	r->38	s->125	t->84	u->30	v->54	y->5	Ö->2	ä->9	å->6	ö->15	
ed,	 ->15	
ed.	D->5	E->1	F->1	H->2	I->1	J->1	K->1	V->2	
eda	 ->74	,->3	g->1	k->1	m->158	n->327	r->25	s->8	t->1	
edb	e->16	o->170	r->1	
edd	 ->24	a->19	e->83	
ede	 ->3	.->1	l->236	n->3	p->2	r->97	s->44	t->3	
edf	i->2	ö->20	
edg	a->1	e->20	i->2	å->2	ö->2	
edh	j->1	
edi	 ->1	.->1	a->8	c->1	e->9	g->3	n->9	t->3	
edj	a->3	e->73	o->1	
edk	v->1	ä->5	
edl	a->4	e->356	i->14	ä->4	
edm	o->3	
edn	i->83	
edo	 ->4	f->1	g->10	m->12	v->4	
edr	a->172	e->1	i->15	o->1	u->1	ä->37	
eds	 ->8	,->1	.->1	a->4	b->2	e->2	f->3	k->6	p->23	s->28	t->5	u->1	
edt	 ->2	,->2	e->14	
edu	c->4	r->1	
edv	e->61	r->12	ä->1	
edö	m->55	
ee-	f->1	l->1	
ee.	D->1	
eel	a->2	l->6	
een	d->63	h->5	
eer	 ->3	,->4	J->1	b->3	i->1	s->5	
ees	 ->1	
eex	e->1	
ef 	h->1	
efa	d->1	l->20	n->1	r->5	t->12	
efe	l->1	n->1	r->22	
eff	e->148	i->1	
efi	n->78	t->5	
efl	e->7	ä->1	
efo	g->32	l->43	n->2	r->149	
efr	a->10	i->12	ä->1	å->2	
eft	e->373	
efu	l->18	s->2	
efä	l->1	n->1	r->10	s->10	
efö	l->1	r->22	
eg 	a->1	b->1	f->11	g->1	h->2	i->13	j->1	l->2	m->4	n->2	o->2	p->3	s->7	t->4	u->1	v->1	
eg,	 ->3	
eg.	D->2	
ega	 ->36	!->4	,->3	.->1	d->2	g->4	l->22	n->16	p->1	s->2	t->45	
egd	r->1	
ege	.->1	?->1	l->50	m->3	n->111	r->423	t->27	
egi	 ->17	,->4	.->3	c->1	e->19	m->3	n->8	o->252	p->1	s->37	t->18	u->3	
egl	a->24	e->126	i->1	
egn	a->45	i->1	
ego	i->2	r->12	
egr	a->21	e->36	i->25	u->2	ä->68	
egu	r->1	
egä	r->60	
egå	 ->2	e->15	n->4	r->3	s->3	t->3	
eha	b->1	g->2	n->88	r->2	v->2	
ehi	n->1	
eho	v->67	
ehr	e->7	
ehä	f->1	
ehå	l->120	
ehö	j->1	l->5	r->18	v->147	
eid	o->2	
eij	s->2	
eik	.->1	h->4	
eil	l->1	
ein	.->1	c->1	d->3	e->6	s->3	z->2	
eir	a->5	
eis	e->2	k->711	m->2	
eiv	r->1	
eix	a->5	
eiz	,->1	
ej 	a->3	b->3	i->1	k->1	l->2	n->1	t->1	ä->1	
ej,	 ->10	
ej.	(->1	E->1	I->1	R->1	
ejd	a->3	o->1	
ejo	r->3	
eju	d->4	
ejä	l->3	
ek 	h->1	o->1	s->1	
eka	 ->27	,->2	.->2	d->12	n->39	r->17	s->7	t->16	
eke	l->4	n->4	r->2	
ekh	e->4	
eki	n->1	s->8	
ekl	a->59	e->2	ö->1	
ekn	i->49	o->3	
eko	d->8	k->1	l->15	m->72	n->291	r->3	s->5	
ekr	e->16	i->1	y->1	ä->30	
eks	a->6	
ekt	 ->113	"->1	,->8	.->12	:->1	;->1	?->2	a->21	e->131	i->373	o->107	r->12	u->3	y->1	ö->7	
eku	l->4	n->3	
ekv	a->7	e->62	o->1	ä->16	
eky	m->16	
ekä	m->41	n->1	
el 	(->2	-->5	1->16	2->14	3->8	4->9	5->6	6->12	7->8	8->16	9->3	B->1	H->1	K->1	N->1	P->1	R->1	a->104	b->8	d->9	e->2	f->39	g->5	h->10	i->25	k->9	l->4	m->11	n->7	o->48	p->30	r->5	s->31	t->9	u->7	v->6	ä->18	å->1	ö->1	
el!	 ->2	M->1	T->1	
el,	 ->54	
el-	 ->3	I->2	S->6	
el.	B->1	D->12	E->3	F->1	G->1	I->1	J->4	M->4	N->2	S->3	T->1	V->10	Ä->2	
el:	 ->5	
el;	 ->1	
el?	E->1	J->1	
ela	 ->146	,->1	?->1	d->12	g->6	k->24	n->57	r->97	s->21	t->55	y->2	
elb	a->20	e->1	r->1	u->15	y->1	
ele	d->2	f->2	g->21	k->14	m->9	n->40	r->10	s->23	t->1	v->11	
elf	e->1	r->3	t->1	u->1	
elg	a->1	e->1	i->18	
elh	a->3	e->21	j->8	o->1	
eli	g->42	k->1	l->1	m->6	n->1	s->15	
elk	r->1	u->1	v->1	
ell	 ->101	"->2	,->4	-->3	.->10	a->564	b->2	e->449	f->3	i->10	m->1	r->10	s->1	t->116	å->4	ö->2	
elm	a->2	e->1	s->1	ä->2	
eln	 ->16	,->2	.->1	i->42	s->2	
elo	d->1	g->2	n->2	p->16	r->3	
elp	l->1	r->1	u->2	
elr	a->1	e->4	i->1	o->1	u->1	y->1	ä->3	
els	 ->24	-->1	a->1	d->1	e->408	f->4	h->2	i->23	k->18	l->6	m->12	n->1	o->10	p->6	s->46	t->92	u->3	v->1	y->3	ä->102	
elt	 ->184	,->1	.->12	;->1	?->1	a->56	i->3	o->2	r->1	ä->4	
elu	t->2	x->1	
elv	a->3	e->21	i->40	ä->4	
ely	s->4	
elz	e->1	
elä	g->31	m->3	n->1	t->1	
elö	n->2	s->4	
em 	-->2	2->1	a->14	b->3	d->14	e->11	f->34	g->4	h->6	i->29	j->1	k->8	l->2	m->28	n->5	o->26	p->13	r->1	s->109	t->6	u->5	v->8	ä->8	å->15	ö->2	
em,	 ->35	
em.	 ->3	(->1	.->1	A->2	B->2	D->15	E->2	F->3	G->1	H->5	I->1	J->7	K->1	M->5	N->3	O->1	P->1	R->1	S->2	T->1	U->1	V->9	
em:	 ->5	
em;	 ->2	
em?	D->1	M->1	
ema	 ->3	,->1	g->4	l->1	n->24	r->1	s->1	t->17	
emb	a->1	e->45	l->1	r->1	u->6	y->1	
eme	d->2	l->67	n->457	s->4	t->117	
emf	ö->1	
emh	ö->14	
emi	,->1	g->2	k->6	n->6	s->15	t->3	ä->10	
eml	a->3	i->6	ä->3	ö->5	
emm	a->26	e->1	
emo	g->3	k->137	m->3	n->14	t->101	
emp	e->114	l->8	o->2	u->1	
ems	 ->3	-->1	a->2	k->7	l->36	r->1	s->284	
emt	 ->4	e->16	i->3	o->5	
emv	i->1	
emy	n->1	
emä	n->37	r->5	s->1	
emå	l->16	n->1	r->3	
emö	d->3	j->4	n->1	t->7	
en 	"->14	(->14	,->1	-->53	1->50	2->25	3->11	4->4	5->1	6->1	7->3	9->3	A->6	B->7	C->3	D->5	E->19	F->3	G->4	H->1	I->5	J->4	K->12	L->3	M->1	N->2	P->6	R->5	S->5	T->5	U->2	V->1	W->1	X->1	a->1039	b->352	c->22	d->407	e->467	f->904	g->358	h->458	i->774	j->111	k->448	l->129	m->587	n->229	o->856	p->364	r->268	s->1060	t->377	u->213	v->390	w->1	y->5	z->2	Ö->1	ä->274	å->59	ö->116	
en!	 ->4	N->2	R->1	
en"	 ->5	,->3	.->4	
en)	 ->4	(->2	,->1	.->2	J->1	N->1	
en,	 ->715	
en-	S->1	
en.	 ->20	"->1	(->2	)->11	.->13	1->1	A->22	B->4	C->1	D->221	E->35	F->45	G->3	H->63	I->32	J->102	K->27	L->9	M->52	N->20	O->28	P->18	R->9	S->40	T->19	U->10	V->87	Ä->8	Å->2	Ö->2	
en:	 ->24	F->1	
en;	 ->17	
en?	.->1	D->7	E->1	F->4	H->2	I->1	J->2	K->2	N->1	V->8	Ä->3	
enF	r->3	
enH	e->2	
enI	 ->1	
enJ	a->2	
enN	ä->5	
ena	 ->119	,->16	.->13	;->1	?->1	d->33	n->9	r->89	s->89	t->3	u->1	v->3	
enb	a->66	e->8	u->2	
enc	e->1	
end	 ->6	!->2	,->2	-->1	a->158	b->1	e->400	i->1	o->5	r->1	s->2	t->7	é->1	ö->1	
ene	f->5	l->1	m->1	n->3	r->177	t->3	z->1	
enf	r->1	ä->1	ö->7	
eng	a->74	e->20	u->2	ä->1	ö->3	
enh	a->2	e->193	ä->32	å->1	
eni	 ->2	.->1	e->2	g->14	n->89	s->2	
enj	ö->2	
enk	e->36	l->19	o->2	ä->1	
enl	i->134	ö->1	
enn	a->578	d->1	e->34	i->24	
eno	m->450	r->32	v->3	
enp	r->1	
enr	e->3	y->1	ö->1	
ens	 ->906	!->1	,->22	-->2	.->13	/->1	:->1	?->2	a->215	b->12	d->5	e->237	f->8	h->4	i->53	k->408	m->11	n->9	o->3	p->81	r->20	s->27	t->8	u->2	v->12	ä->2	
ent	 ->287	,->28	.->35	a->144	e->644	f->6	i->101	k->1	l->207	o->1	p->2	r->128	s->47	t->1	u->25	v->2	y->13	ä->2	
enu	m->5	s->1	t->1	
env	e->1	i->5	ä->8	
enz	 ->12	)->2	,->3	F->1	b->1	
enÄ	r->1	
enä	g->1	m->1	t->1	
enå	d->1	
enè	v->3	
enö	r->3	
eog	r->8	
eol	o->5	
eom	r->3	
eon	a->1	i->1	l->1	
eor	d->1	e->2	
eos	t->2	
eot	e->1	
ep 	a->1	m->1	
epa	 ->15	,->1	d->8	r->31	s->7	t->5	
epe	s->1	
eph	e->3	
epn	i->1	
epo	k->4	l->2	s->1	t->5	
epp	 ->12	,->1	a->1	e->11	s->8	
epr	e->24	i->2	o->2	
eps	i->1	k->1	
ept	 ->2	.->2	a->44	e->64	i->14	
epu	b->19	
er 	(->4	-->48	1->31	2->7	3->2	4->3	5->2	6->1	7->2	8->3	9->3	A->6	B->5	C->2	D->2	E->36	F->7	G->7	H->2	I->10	J->5	K->3	L->9	M->3	N->4	O->3	P->2	R->2	S->9	T->6	U->4	V->1	[->1	a->996	b->131	c->12	d->573	e->320	f->515	g->96	h->183	i->470	j->121	k->187	l->70	m->354	n->107	o->611	p->219	r->92	s->746	t->238	u->145	v->272	y->1	Ö->4	ä->140	å->36	ö->34	
er!	 ->71	"->2	D->5	E->1	J->3	M->1	V->2	
er"	 ->4	)->1	,->1	.->1	
er)	 ->4	F->2	J->1	K->1	T->1	
er,	 ->476	
er-	b->1	k->1	n->1	p->11	r->1	
er.	 ->17	(->2	)->1	-->3	.->5	9->1	A->11	B->8	C->1	D->124	E->23	F->26	G->3	H->18	I->23	J->59	K->23	L->5	M->22	N->12	O->15	P->8	R->3	S->14	T->16	U->6	V->48	Ä->9	Å->2	
er:	 ->19	
er;	 ->7	
er?	-->1	.->1	B->1	D->1	E->1	H->3	J->1	K->1	M->1	P->1	T->1	V->2	Ä->1	
erH	e->1	
erJ	a->1	
erM	e->1	
erN	ä->2	
era	 ->629	!->1	"->1	,->12	.->27	d->235	h->1	l->78	n->97	r->278	s->250	t->170	y->1	
erb	,->1	a->5	e->18	i->7	j->20	l->3	r->4	ö->12	
erc	e->1	
erd	a->41	e->4	o->3	r->14	s->3	ö->1	
ere	 ->2	.->1	d->59	g->3	l->16	n->265	r->20	s->1	t->8	x->6	
erf	a->30	e->7	i->6	l->3	o->27	r->8	u->2	ö->27	
erg	 ->4	a->2	e->33	i->121	n->1	r->19	ä->1	å->16	
erh	a->6	e->284	u->2	ä->3	å->12	ö->17	
eri	 ->17	,->7	-->1	.->3	a->23	b->4	e->54	f->7	g->26	k->28	l->2	m->9	n->745	o->86	p->1	s->5	t->1	u->1	ö->8	
erk	 ->27	,->3	.->4	?->1	a->207	e->46	l->211	n->15	o->7	r->2	s->71	t->8	u->1	ä->42	
erl	a->8	e->10	i->121	y->2	ä->61	å->11	
erm	a->12	e->4	i->11	o->3	å->1	ö->2	
ern	 ->50	,->9	.->12	/->2	a->1570	d->3	e->14	f->1	i->27	s->13	t->6	ö->1	
ero	d->5	e->69	g->1	i->1	m->1	n->1	p->1	r->24	t->1	
erp	a->2	o->4	r->2	
err	 ->494	a->48	e->9	i->147	o->12	ä->1	å->14	ó->3	ö->1	
ers	 ->65	,->1	-->1	a->10	e->8	h->1	i->42	k->51	l->1	m->1	o->298	p->22	t->147	u->3	v->7	y->1	ä->35	å->1	ö->48	
ert	 ->66	!->1	,->4	.->1	a->26	e->37	g->3	h->2	i->81	k->17	o->2	r->11	u->1	y->38	ä->2	
eru	p->34	s->2	t->3	
erv	a->36	e->13	i->82	j->3	r->1	t->1	u->3	ä->48	
ery	,->1	k->1	
erä	g->1	k->4	n->17	t->35	
erå	r->12	t->1	
erö	m->2	r->42	s->5	v->3	
es 	-->2	1->3	2->1	3->1	A->1	D->3	G->1	S->1	V->1	W->1	a->47	b->11	d->20	e->20	f->42	g->3	h->11	i->54	j->2	k->15	l->5	m->15	n->12	o->21	p->10	r->16	s->24	t->20	u->15	v->12	y->1	ä->4	å->1	ö->7	
es"	.->1	
es,	 ->17	
es-	 ->6	C->1	
es.	)->1	A->1	D->2	F->1	H->1	I->1	J->1	K->1	M->2	O->1	R->2	U->1	V->2	
es;	 ->1	
esa	 ->14	,->2	.->1	m->7	n->1	r->2	t->7	u->1	
esb	e->2	
esd	i->2	
ese	 ->1	g->2	k->3	n->49	r->11	t->1	
esf	o->1	r->4	ö->1	
esg	e->1	i->1	å->3	
esh	a->4	
esi	d->15	k->2	s->12	t->2	
esk	a->120	e->3	i->3	r->51	v->1	y->6	å->1	
esl	a->26	i->2	o->11	u->241	ä->1	å->69	ö->3	
esm	a->2	i->10	ä->3	
esn	å->4	
eso	l->100	n->4	r->1	
esp	.->2	a->5	e->88	o->7	r->9	
esq	u->1	
esr	a->2	ö->1	
ess	 ->134	"->1	,->2	.->13	?->1	a->402	b->5	e->176	h->1	i->19	k->3	m->1	n->1	o->6	r->3	t->1	u->62	v->4	
est	 ->47	,->1	?->1	a->42	e->44	i->23	n->1	o->6	r->11	s->1	u->7	y->1	ä->181	å->61	ö->1	
esu	l->116	r->50	t->7	
esv	a->18	i->10	ä->7	
esy	n->1	s->1	
esä	t->6	
esö	k->9	r->2	
et 	"->11	(->19	,->1	-->33	1->14	2->2	A->5	B->3	C->1	D->2	E->15	F->1	G->2	I->2	K->4	L->2	M->4	P->4	R->2	S->5	T->2	V->3	a->772	b->224	c->9	d->116	e->204	f->947	g->353	h->336	i->496	j->35	k->283	l->100	m->402	n->136	o->517	p->203	r->117	s->773	t->207	u->112	v->374	y->7	Ö->1	ä->832	å->30	ö->38	
et!	(->1	.->2	H->1	K->1	P->1	
et"	 ->5	,->2	.->2	
et)	 ->6	,->3	.->4	N->1	
et,	 ->512	
et-	 ->1	f->1	
et.	 ->17	(->3	)->4	-->1	.->3	1->1	A->12	B->4	D->126	E->28	F->28	H->34	I->27	J->80	K->7	L->6	M->42	N->17	O->14	P->12	R->4	S->18	T->12	U->3	V->56	Ä->2	Å->3	Ö->1	
et:	 ->13	
et;	 ->6	
et?	 ->1	.->2	A->1	D->3	H->3	I->1	J->2	K->2	N->3	O->1	R->1	S->1	V->3	Ä->1	
etJ	a->1	
eta	 ->128	,->4	.->3	?->1	b->13	d->2	g->207	k->1	l->136	n->36	p->5	r->42	s->2	t->14	
etb	e->1	
etc	.->5	?->1	
etd	e->1	
ete	 ->116	,->11	.->29	?->3	c->12	e->3	n->501	r->448	s->12	t->63	
etf	r->2	ö->9	
eth	 ->1	
eti	k->2	n->2	s->9	t->1	
etj	ä->1	
etk	o->16	r->1	
etl	i->36	
etm	a->1	ä->1	
etn	a->17	i->14	
eto	d->29	n->46	r->3	
etp	l->3	o->11	
etr	a->25	o->13	u->1	y->4	ä->153	
ets	 ->339	,->2	-->5	.->1	a->22	b->12	c->4	d->4	e->6	f->31	g->19	h->2	i->3	k->15	l->51	m->25	n->9	o->16	p->97	r->30	s->12	t->92	u->5	v->7	y->1	å->2	
ett	 ->1488	,->7	.->10	:->2	a->1041	e->21	i->7	o->4	s->15	v->1	
etu	n->1	t->10	
etv	i->30	
ety	 ->1	-->1	d->129	
etä	n->293	r->6	
etå	r->10	
etê	t->2	
etö	v->1	
eug	e->2	
eum	 ->1	
eun	d->3	
eur	o->416	
eus	s->1	
eut	b->1	i->1	r->3	s->3	v->4	
ev 	a->3	d->4	f->3	i->3	k->1	n->1	o->4	s->1	t->3	u->2	
ev.	F->1	
eva	 ->17	,->1	?->1	k->6	l->6	n->12	r->22	t->2	
evd	e->2	
eve	b->1	k->1	l->2	n->21	r->20	
evi	d->18	g->3	l->48	s->70	t->1	
evl	i->3	å->1	
evn	a->12	
evo	l->1	
evs	 ->6	
evt	 ->4	
evä	c->3	r->14	
evå	n->2	
ew 	Y->1	
ewi	e->1	
ewo	o->2	
ex 	a->6	e->1	f->1	m->11	p->2	t->2	ö->1	
ex,	 ->1	
ex.	 ->20	J->1	
exa	,->1	k->18	m->16	n->2	s->2	
exc	e->5	
exe	m->117	
exi	b->27	k->1	l->2	s->20	
exk	l->3	
exm	å->1	
exp	a->6	e->45	l->3	o->6	
ext	 ->13	,->5	.->1	e->34	o->1	r->36	
exu	e->3	
exv	ä->1	
ey 	C->3	
eye	r->3	
eyh	u->1	
ez 	G->1	a->1	o->1	t->1	
ez,	 ->2	
ez-	k->2	
ezu	e->1	
eäg	a->2	
eåt	e->1	
f -	 ->1	
f H	i->2	
f a	v->1	
f e	l->1	x->1	
f f	ö->5	
f h	a->3	
f i	 ->1	n->2	
f k	u->1	
f l	i->1	
f n	o->1	
f o	c->4	m->1	
f s	o->4	
f t	h->1	
f u	t->1	
f ä	g->1	
f, 	h->1	m->1	o->1	p->1	s->1	
f- 	o->2	
f-M	a->2	
f.D	e->1	ä->1	
f.E	n->1	
f.J	a->1	
f.d	.->2	
fa 	a->3	b->1	d->2	e->5	f->3	i->1	k->3	m->1	o->1	r->1	s->2	u->2	
fa,	 ->2	
fa.	M->1	
fab	e->1	r->1	
fac	k->4	
fad	d->1	e->10	
fae	l->3	
fai	l->1	
fak	t->136	
fal	a->1	d->15	l->231	s->4	
fam	i->15	
fan	d->42	n->16	t->14	
far	 ->36	,->4	.->9	:->1	?->1	a->182	e->26	h->2	i->2	l->59	m->1	n->1	o->4	s->1	t->81	v->9	
fas	 ->4	,->2	.->1	c->11	e->4	n->3	o->1	t->112	
fat	 ->5	.->4	s->2	t->257	
fau	n->1	
fav	o->1	
fax	a->1	
fbe	s->1	
fdr	a->1	
feb	r->16	
fed	e->12	
fek	t->162	
fel	 ->11	!->1	,->4	.->4	a->13	b->2	e->1	k->1	r->1	s->1	
fem	 ->27	,->1	:->1	p->1	t->24	å->3	
fen	 ->17	,->5	-->1	.->4	o->3	s->4	t->80	
fer	 ->30	"->1	,->10	.->6	a->4	e->182	i->2	n->12	t->2	
fes	s->8	t->1	
fet	y->1	
ff 	n->1	o->2	
ff,	 ->1	
ff-	 ->2	
ffa	 ->25	,->2	.->1	d->9	n->42	r->51	s->5	t->10	
ffb	e->1	
ffe	k->153	n->86	r->18	
ffi	c->7	
ffl	a->1	i->2	
ffp	r->2	
ffr	a->9	e->14	o->15	ä->28	
ffä	r->12	
fhj	ä->1	
fi 	o->1	p->1	s->1	
fi,	 ->1	
fi.	D->1	V->1	
fic	e->39	i->8	k->27	
fid	e->2	
fie	n->34	r->27	
fik	 ->5	-->1	.->2	a->22	e->3	l->1	t->7	
fil	 ->1	.->2	m->2	o->5	s->1	t->1	
fin	 ->2	-->3	.->1	a->83	g->2	i->38	l->5	n->416	s->6	t->10	
fiq	u->1	
fir	a->3	
fis	k->61	
fit	-->5	
fjo	l->4	r->9	
fjä	r->11	
fkr	i->1	
fla	g->30	m->4	
fle	k->7	r->99	s->25	x->27	
fli	c->1	g->2	k->16	r->1	t->2	
flo	d->4	r->1	t->4	
flu	t->14	
fly	g->14	k->16	r->1	t->30	
flä	c->1	k->1	
flö	d->4	
fma	n->1	
fob	i->1	
fod	e->10	
fog	 ->1	a->30	e->27	
fok	u->5	
fol	k->122	
fon	,->1	d->126	e->1	
for	 ->2	a->1	c->1	d->89	m->351	s->81	t->194	u->5	ê->1	
fos	s->3	t->1	
fot	b->1	f->1	s->2	
fpr	o->2	
fra	 ->4	,->3	d->1	k->11	m->658	n->38	r->1	s->16	
fre	d->93	e->3	k->1	n->14	s->5	
fri	 ->15	,->1	-->8	a->31	e->6	g->6	h->115	k->7	s->16	t->5	v->12	
fro	d->4	n->4	r->15	
fru	 ->67	,->1	k->16	s->2	t->1	
fry	s->3	t->2	
frä	c->1	m->144	t->28	
frå	g->816	n->617	
fsi	t->1	
fst	r->4	ö->2	
ft 	2->1	a->9	b->2	d->5	e->5	f->14	g->1	h->1	i->6	k->2	l->1	m->6	n->4	o->6	p->5	r->1	s->18	t->5	u->2	v->4	ä->4	
ft!	H->1	
ft,	 ->13	
ft.	 ->1	A->1	D->3	E->1	H->1	J->1	M->1	O->1	V->4	
ft:	 ->1	
ft?	 ->1	N->1	
fta	 ->70	,->1	.->1	d->6	n->7	r->44	s->9	t->8	
ftb	u->1	
fte	 ->20	,->1	.->2	l->1	n->42	r->496	t->26	
ftf	u->12	
fti	g->49	
ftl	i->8	
ftn	i->113	
fto	m->1	n->1	r->3	
fts	-->1	a->4	f->2	l->2	m->1	o->1	p->4	r->1	s->2	t->1	v->1	ä->1	
ftt	a->1	r->4	
ftv	e->8	
ful	l->149	t->1	
fun	d->18	g->54	k->32	n->12	
fus	e->1	i->8	k->1	
fut	t->1	
fyl	l->62	
fyr	a->25	t->3	
fys	i->9	
fäd	e->1	
fäk	t->1	
fäl	h->1	l->114	t->6	
fän	g->2	
fär	 ->9	a->1	d->36	e->12	g->3	l->2	r->2	s->2	
fäs	t->25	
få 	1->1	E->1	G->1	a->5	b->8	d->16	e->41	f->13	g->2	h->2	i->7	k->6	l->7	m->9	n->3	o->6	p->9	r->5	s->25	t->22	u->3	v->11	ä->1	å->1	ö->1	
få,	 ->3	
få.	E->1	G->1	V->1	
fåg	e->3	l->6	
fån	g->14	
får	 ->182	,->2	?->1	k->1	
fås	 ->1	
fåt	a->1	t->57	
fér	e->1	
föd	d->2	e->4	n->1	o->1	s->1	
fög	a->2	
föl	j->158	l->7	
fön	s->1	
för	 ->3683	"->1	,->27	.->17	:->3	;->1	?->5	a->512	b->224	d->276	e->789	f->135	g->6	h->191	i->16	k->93	l->123	m->69	n->74	o->79	p->26	r->60	s->1251	t->159	u->78	v->156	ä->73	å->3	ö->8	
föt	t->3	
g (	1->1	E->1	a->2	r->1	å->1	
g -	 ->23	,->2	
g 1	 ->2	,->2	0->5	1->1	2->1	3->1	5->1	7->2	8->2	9->5	
g 2	,->2	0->2	2->3	3->1	6->1	
g 3	 ->1	4->1	7->1	8->3	
g 4	 ->1	.->2	3->1	4->1	5->3	
g 5	,->2	
g 6	 ->2	0->1	8->1	
g 8	0->2	
g D	e->1	
g E	c->1	u->2	
g F	ä->1	
g G	a->1	
g H	a->14	
g I	N->1	V->2	r->1	
g O	L->1	
g T	a->1	
g V	I->1	
g [	K->1	
g a	b->1	c->3	j->1	k->1	l->12	n->113	r->7	s->2	t->203	v->371	
g b	a->22	e->83	i->3	l->13	o->5	r->4	y->3	ä->2	ö->10	
g c	i->2	
g d	a->1	e->73	i->6	j->1	o->5	r->3	y->1	ä->17	å->1	ö->3	
g e	.->1	f->8	k->1	l->22	m->10	n->34	r->15	t->20	u->1	v->1	x->4	
g f	a->4	e->1	i->12	o->7	r->118	u->7	ä->1	å->16	ö->297	
g g	a->5	e->22	i->3	j->5	l->12	o->1	r->27	ä->12	å->2	ö->4	
g h	a->155	e->14	i->4	j->3	o->58	u->4	ä->25	å->15	ö->8	
g i	 ->210	,->1	.->1	a->1	h->1	n->163	r->1	v->1	
g j	a->2	o->1	u->5	ä->3	
g k	a->80	l->5	n->2	o->85	r->5	u->8	v->2	ä->11	ö->1	
g l	a->12	e->7	i->9	y->7	ä->14	å->3	ö->6	
g m	a->18	e->117	i->28	o->27	y->14	ä->3	å->41	ö->2	
g n	a->7	e->4	i->14	o->8	r->2	u->8	y->3	ä->26	å->2	ö->3	
g o	b->3	c->264	e->1	f->5	l->1	m->113	n->2	r->4	s->1	
g p	a->2	e->11	l->2	o->13	r->12	u->7	å->116	
g r	a->5	e->41	i->7	o->8	u->1	y->1	ä->11	å->5	ö->15	
g s	a->24	e->25	i->23	j->25	k->186	l->2	o->233	p->2	t->41	u->1	v->3	y->10	ä->50	å->11	
g t	.->1	a->61	e->3	i->222	o->3	r->120	v->6	y->49	ä->17	
g u	n->27	p->57	r->1	t->62	
g v	a->39	e->35	i->295	o->1	ä->33	å->2	
g y	r->1	t->1	
g Ö	s->2	
g ä	g->2	l->1	n->14	r->164	v->6	
g å	 ->3	k->1	s->4	t->31	
g ö	k->3	n->6	p->1	v->18	
g!"	.->1	
g!H	a->1	
g!J	a->1	
g" 	a->1	o->1	s->1	
g",	 ->2	
g".	E->1	J->1	N->1	
g) 	i->2	o->2	
g),	 ->1	
g).	V->1	
g)N	ä->1	
g, 	B->1	I->1	O->1	a->14	b->8	d->24	e->33	f->40	g->7	h->14	i->22	j->7	k->7	l->8	m->34	n->15	o->40	p->9	r->2	s->59	t->11	u->17	v->28	ä->10	å->3	ö->1	
g-P	M->1	
g. 	D->3	E->1	F->1	H->1	M->1	P->1	S->2	
g.(	A->2	
g.)	F->2	H->1	
g..	 ->3	(->1	
g.A	l->4	n->2	r->1	v->6	
g.B	e->2	i->1	r->1	
g.D	a->2	e->100	i->1	o->2	ä->10	
g.E	f->4	m->1	n->7	r->2	t->1	u->3	
g.F	l->1	r->9	ö->19	
g.G	e->4	r->1	
g.H	a->2	e->20	u->2	y->1	ä->1	ö->1	
g.I	 ->20	n->3	
g.J	a->62	u->1	
g.K	a->2	o->13	
g.L	e->1	i->2	å->3	
g.M	a->9	e->9	i->1	y->1	å->4	ö->1	
g.N	a->2	i->3	u->3	ä->3	å->1	
g.O	a->1	c->11	f->1	m->10	
g.P	P->1	a->2	r->2	å->2	
g.R	a->1	e->2	
g.S	a->3	e->1	k->2	l->4	y->1	å->1	
g.T	a->2	i->4	r->1	
g.U	n->2	
g.V	a->6	i->29	å->2	
g.a	.->1	
g.Ä	r->4	
g: 	D->1	d->3	e->1	f->1	h->1	i->1	j->1	
g:D	e->2	
g; 	d->2	e->1	f->3	m->1	s->1	
g?D	e->4	ä->1	
g?F	i->1	r->1	ö->1	
g?H	u->1	ä->1	
g?J	a->1	o->1	
g?O	l->1	
g?T	y->1	
g?V	a->1	
g?Ä	r->1	
gNä	s->1	
ga 	"->2	-->8	2->1	3->1	B->3	E->8	F->7	H->3	I->1	J->3	K->1	L->1	M->1	N->2	R->2	S->3	a->189	b->75	c->2	d->64	e->39	f->228	g->41	h->33	i->68	j->3	k->69	l->31	m->84	n->59	o->201	p->48	r->116	s->199	t->60	u->44	v->49	y->2	ä->42	å->26	ö->14	
ga!	 ->1	D->1	F->2	J->1	Ä->1	
ga,	 ->91	
ga.	 ->2	(->1	-->1	A->4	D->13	E->3	F->6	H->5	I->6	J->14	M->6	N->3	O->3	P->2	S->2	T->1	U->1	V->12	Ä->1	
ga/	h->1	
ga:	 ->11	
ga;	 ->1	
ga?	.->1	D->1	F->1	
gad	 ->21	,->1	.->4	e->40	o->1	
gag	e->18	n->11	å->6	
gak	t->1	
gal	 ->19	,->4	a->7	e->1	i->2	l->1	n->1	s->7	t->9	u->3	
gam	 ->1	,->1	l->28	m->4	
gan	 ->217	"->1	,->20	.->18	:->5	;->1	?->1	d->388	e->9	i->66	s->30	t->6	
gap	r->1	
gar	 ->418	!->1	"->1	)->1	,->64	-->1	.->96	:->7	;->1	?->1	a->96	d->2	e->337	i->17	l->3	m->14	n->286	s->12	v->1	ä->1	
gas	 ->41	,->8	.->10	a->1	e->5	k->2	t->56	ä->19	
gat	 ->24	,->3	.->2	a->1	e->2	i->43	o->15	s->7	
gau	 ->7	,->5	.->1	M->1	b->1	s->3	
gav	 ->14	,->1	a->1	s->5	
gba	r->15	
gbe	r->1	
gbl	a->1	
gbo	x->1	
gbr	o->1	
gby	g->1	
gd 	a->2	b->2	f->5	g->1	i->4	l->1	n->1	o->6	p->2	s->2	y->1	ä->1	å->1	
gd,	 ->1	
gd.	D->2	
gda	 ->8	.->1	
gde	 ->4	n->36	r->5	s->1	
gdo	m->27	
gdp	u->4	
gdr	a->2	
gds	b->1	k->1	o->4	r->2	t->1	u->1	
gdy	r->1	
ge 	E->1	F->2	a->15	b->7	d->19	e->32	f->4	g->3	h->6	i->6	j->1	k->7	m->7	n->4	o->19	p->12	r->10	s->25	t->4	u->13	v->10	ä->2	å->1	
ge,	 ->4	
ge.	 ->1	H->1	J->2	O->1	V->1	
ge?	H->1	
ged	i->6	
gef	ä->10	
gek	o->1	
gel	 ->4	,->1	b->16	i->1	l->2	m->3	n->8	r->2	s->32	v->20	ä->23	
gem	a->13	e->386	
gen	 ->1426	!->1	"->3	,->130	.->134	:->9	;->3	?->7	I->1	a->20	b->1	d->13	e->39	f->5	g->1	h->39	j->2	k->2	o->419	r->1	s->119	t->99	u->1	ä->1	
geo	g->8	s->2	
ger	 ->392	!->65	,->30	.->16	:->6	;->1	M->1	a->130	b->1	e->6	i->327	k->1	l->3	m->1	n->29	p->2	s->1	v->1	
ges	 ->29	,->3	-->1	.->1	b->1	f->1	r->2	t->12	
get	 ->252	)->4	,->28	.->46	:->1	;->1	?->1	a->3	b->1	d->1	e->18	f->11	k->17	m->1	p->14	s->29	t->25	u->10	å->10	ö->1	
gfa	l->15	
gfl	ö->1	
gfo	n->1	r->20	
gfr	i->1	u->1	
gfu	n->1	
gfä	r->2	
gfö	r->5	
gg 	d->2	f->2	g->1	h->2	i->5	k->1	l->1	m->2	o->1	p->3	s->2	t->4	u->4	v->1	
gg"	 ->1	
gg,	 ->8	
gg.	D->1	F->2	K->1	M->1	N->1	
gg;	 ->1	
gga	 ->144	,->1	d->3	n->111	s->14	
ggb	o->1	
ggd	 ->2	e->2	
gge	 ->1	l->1	n->8	r->133	t->6	
ggh	e->6	
ggi	g->3	
ggj	o->13	
ggl	i->1	
ggn	a->19	i->28	
ggo	r->2	
ggr	a->13	e->1	
ggs	 ->19	,->1	b->1	f->1	k->1	t->1	
ggt	 ->4	s->1	
ggå	 ->1	s->1	
ggö	r->21	
gh 	l->1	m->1	
gh.	V->1	
ghe	t->851	
ght	 ->2	s->1	
ghå	l->2	
gi 	-->2	b->1	f->5	g->2	h->2	i->1	k->1	l->1	m->2	o->8	s->7	t->2	
gi,	 ->6	
gi-	,->1	
gi.	.->1	A->1	D->1	E->2	F->2	J->1	M->1	V->1	
gia	g->1	n->6	
gib	e->3	
gic	e->1	k->22	
gie	f->4	n->11	r->18	t->2	
gif	o->1	t->101	ö->4	
gig	a->5	g->1	t->4	
gii	m->1	
gik	 ->1	,->2	.->3	a->1	e->2	o->1	ä->37	
gil	l->2	t->26	
gim	e->3	i->1	y->1	
gin	 ->8	,->2	.->2	a->7	e->1	s->1	ä->1	
gio	n->252	r->2	
gip	l->1	o->2	r->5	
gis	e->4	i->70	k->66	n->1	s->1	t->20	ä->7	
git	 ->96	,->2	.->5	a->1	i->18	s->27	
giu	m->3	
giv	a->63	e->32	i->15	l->1	n->11	
giz	i->5	
giä	k->1	
giå	t->1	
giö	s->4	
gjo	r->136	
gkr	a->3	
gku	l->1	
gkö	r->1	
gla	 ->7	d->30	n->1	r->19	s->5	
gle	d->5	r->126	s->1	w->2	
gli	g->87	n->2	
glj	u->1	
glo	b->12	
glu	p->1	
glä	d->40	n->1	
glö	m->21	
gm 	e->1	
gma	r->1	t->3	
gme	t->6	
gmä	r->1	s->2	
gmå	l->1	
gn 	f->3	o->1	
gna	 ->97	,->3	.->2	d->24	l->14	n->1	r->31	s->3	t->7	
gne	 ->8	-->1	l->1	n->2	r->3	s->1	
gni	,->1	n->223	s->1	t->1	v->3	
gno	r->4	
gnu	t->2	
gnä	l->1	
go 	g->1	s->1	å->1	
god	 ->23	.->1	a->37	k->89	o->4	s->38	t->46	
gof	e->1	
gog	e->1	i->4	
goi	s->2	
gol	f->4	v->1	y->1	
gom	 ->4	.->1	å->3	
gon	 ->142	,->5	.->7	b->15	d->3	s->15	t->39	
gor	 ->182	)->1	,->38	.->28	:->4	;->1	?->2	d->52	i->9	l->1	n->31	s->2	ö->4	
gos	k->1	l->1	
got	 ->185	,->2	.->6	?->1	t->20	
gou	 ->1	
gpl	a->4	
gpo	l->2	
gra	 ->158	d->37	f->17	m->238	n->85	r->6	s->1	t->69	v->6	
gre	 ->82	,->1	.->9	d->2	k->7	m->1	n->4	p->26	r->24	s->4	
gri	f->1	k->1	n->1	p->66	t->3	
gro	d->1	g->1	t->1	u->1	v->1	
gru	n->297	p->184	v->1	
gry	m->1	
grä	l->3	m->1	n->134	v->4	
grå	 ->1	z->1	
grö	d->1	j->1	n->18	v->1	
gs 	-->1	a->14	b->2	d->5	e->3	f->15	g->1	h->2	i->11	k->3	m->5	n->2	o->5	p->9	r->2	s->7	t->1	u->7	v->4	
gs,	 ->5	
gs-	 ->12	
gs.	F->1	J->1	L->1	
gsa	k->3	l->1	m->13	n->8	r->9	v->8	
gsb	a->2	e->13	i->11	o->4	r->6	u->1	
gsc	e->5	h->8	
gsd	e->1	i->2	o->1	r->1	
gse	k->6	n->3	r->2	t->5	
gsf	a->9	e->2	i->31	l->1	o->22	r->16	u->12	ä->1	ö->235	
gsg	i->8	r->8	
gsh	a->1	e->1	o->1	
gsi	d->4	k->7	n->12	
gsj	u->2	
gsk	a->1	l->3	o->173	r->16	u->1	v->1	ä->2	
gsl	a->2	i->60	o->1	ä->8	ö->5	
gsm	a->4	e->7	i->1	o->5	ä->4	å->4	ö->4	
gsn	a->6	e->1	i->5	o->1	y->1	ä->2	
gso	m->12	r->2	
gsp	a->4	e->3	l->23	o->22	r->46	u->11	å->1	
gsr	e->23	i->15	u->1	ä->2	å->3	
gss	a->2	e->8	i->3	k->22	p->1	t->23	y->24	ä->16	
gst	 ->14	,->1	.->1	a->28	e->6	i->131	j->5	m->2	r->1	ä->2	
gsu	m->1	t->7	
gsv	e->4	i->33	ä->7	å->2	
gsy	s->2	
gsä	g->3	n->3	r->1	t->1	
gså	r->1	t->5	
gsö	v->1	
gt 	-->7	4->2	:->1	D->1	E->2	G->1	I->1	K->1	R->1	S->1	T->1	a->242	b->34	d->38	e->36	f->129	g->47	h->33	i->55	j->3	k->30	l->15	m->97	n->26	o->81	p->39	r->22	s->149	t->32	u->26	v->48	y->2	ä->17	å->3	ö->6	
gt!	L->1	M->1	
gt,	 ->73	
gt.	 ->1	A->1	D->12	E->3	F->8	G->2	H->5	I->1	J->12	L->2	M->10	N->2	O->3	P->1	S->4	U->1	V->14	Ö->1	
gt:	 ->1	
gt;	 ->1	
gt?	A->1	
gta	r->1	
gte	k->2	r->8	x->2	
gtg	å->11	
gti	d->8	
gto	n->5	
gtr	a->2	
gts	 ->37	,->2	
gtv	i->108	ä->4	
gud	s->2	
gue	,->1	i->1	r->2	s->1	
gul	d->1	t->1	
gum	e->17	m->1	
gur	o->1	
gus	t->1	
guv	e->1	
gva	r->6	t->1	
gve	r->1	
gyn	n->19	
gyp	t->2	
gäc	k->1	
gäl	d->1	l->405	
gän	g->24	
gär	 ->11	.->1	a->34	d->248	n->33	s->1	t->10	
gäv	e->1	
gå 	K->1	a->2	b->2	d->2	e->5	f->9	g->2	h->1	i->27	l->6	m->3	o->3	p->1	s->7	t->13	u->5	v->4	å->1	
gå.	A->1	D->1	F->1	N->1	O->1	S->1	V->1	
gåe	n->101	
gån	g->259	
går	 ->142	,->4	.->8	d->6	
gås	 ->4	,->1	:->1	
gåt	t->36	
gåv	o->2	
göm	m->3	t->1	
gör	 ->190	,->2	.->4	a->389	e->5	i->2	l->2	s->28	
h "	U->1	s->1	t->1	
h (	A->1	
h -	 ->3	o->3	
h 0	 ->1	
h 1	-->1	0->2	3->1	4->1	6->1	7->2	9->13	
h 2	 ->1	,->1	.->1	0->3	1->3	2->1	5->1	7->1	9->1	
h 3	.->1	0->2	3->1	4->1	5->1	:->1	
h 4	.->1	1->2	5->4	7->1	8->2	
h 5	 ->1	.->1	3->1	
h 6	0->1	8->1	
h 7	 ->4	,->2	
h 8	 ->1	,->1	2->6	6->2	9->1	
h 9	 ->2	2->1	4->1	
h A	l->2	m->1	n->1	
h B	P->1	a->1	e->1	r->2	u->1	
h C	.->1	E->1	a->1	y->1	
h D	a->2	e->2	
h E	L->2	U->4	d->1	l->2	m->1	r->1	t->1	u->24	
h F	N->1	P->1	i->2	r->11	
h G	a->2	e->1	o->1	r->3	
h H	e->1	i->1	u->1	
h I	I->2	n->4	r->2	s->5	t->1	
h J	a->1	ö->1	
h K	a->1	i->6	o->1	u->1	
h L	a->3	e->5	
h M	A->1	a->3	e->1	
h N	o->1	y->1	
h O	L->1	n->1	
h P	P->1	S->2	a->9	e->1	o->3	r->1	
h R	a->3	
h S	a->10	c->2	i->1	j->1	o->1	p->1	t->2	w->1	y->8	
h T	a->4	s->1	u->1	y->2	
h U	z->1	
h V	i->1	ä->1	
h W	y->1	
h X	 ->1	
h a	b->1	c->1	d->2	g->2	k->4	l->18	m->4	n->58	p->1	r->15	s->4	t->150	v->32	
h b	a->13	e->52	i->10	l->8	o->5	r->15	u->3	y->2	ä->4	å->1	ö->6	
h c	a->2	e->6	h->2	
h d	a->4	e->467	i->11	j->4	o->9	r->4	u->1	y->1	ä->83	å->24	ö->1	
h e	f->34	g->1	j->1	k->22	l->1	n->90	r->17	t->33	u->9	x->4	
h f	a->14	e->3	i->12	l->10	o->7	r->83	u->9	y->2	ä->1	å->12	ö->168	
h g	a->7	e->43	i->4	j->1	l->3	o->2	r->10	ä->1	å->4	ö->17	
h h	a->46	e->54	i->1	j->4	o->11	u->15	y->2	ä->9	å->16	ö->6	
h i	 ->74	b->3	c->2	d->5	f->1	k->1	l->1	m->2	n->142	r->1	s->2	
h j	a->149	o->5	u->7	ä->1	
h k	a->21	i->1	l->4	n->1	o->129	r->18	u->7	v->10	ä->6	ö->1	
h l	a->17	e->17	i->11	j->1	o->9	u->1	y->3	ä->14	å->19	ö->2	
h m	a->21	e->144	i->39	o->24	u->1	y->8	ä->12	å->22	ö->9	
h n	a->11	e->8	i->9	o->5	u->11	y->13	ä->17	å->5	ö->6	
h o	a->4	b->2	c->10	d->1	e->2	f->6	j->1	k->4	l->8	m->41	n->1	p->2	r->8	s->5	t->1	u->3	
h p	a->25	e->9	l->3	o->17	r->32	å->29	
h r	a->7	e->66	i->9	o->4	u->1	ä->61	å->39	ö->1	
h s	a->43	e->29	i->10	j->6	k->30	l->24	m->2	n->4	o->134	p->9	t->61	u->5	v->12	y->16	ä->33	å->28	ö->2	
h t	.->1	a->20	e->6	h->1	i->60	j->4	o->6	r->18	u->17	v->3	y->14	ä->3	
h u	n->25	p->24	t->57	
h v	a->52	e->23	i->123	ä->26	å->12	ö->1	
h y	n->1	r->1	t->5	
h Ö	V->1	s->6	
h ä	g->2	n->12	r->10	v->31	
h å	 ->4	k->1	s->3	t->29	
h ö	k->3	m->1	n->1	p->13	r->1	s->4	v->20	
h! 	U->1	
h)D	e->1	
h, 	a->1	d->1	f->3	h->1	i->1	n->1	o->1	r->1	s->4	t->1	u->1	
h-B	e->7	
h-a	v->1	
h.D	e->1	
h.E	f->1	
h.F	ö->1	
h.J	a->1	
h.V	i->1	
h/e	l->1	
h: 	V->1	
h?F	r->1	
hI 	o->1	
hII	.->1	
ha 	a->5	b->5	d->10	e->55	f->6	g->5	h->7	i->3	k->10	l->4	m->12	n->10	o->2	p->2	r->3	s->14	t->11	u->5	v->14	y->1	ä->2	å->1	ö->3	
ha,	 ->1	
ha.	A->1	
hab	i->1	l->1	
had	e->85	
haf	t->37	
hag	l->2	
hak	a->1	
hal	l->1	t->1	v->25	
ham	b->1	e->1	m->1	n->39	p->1	
han	 ->117	,->2	;->1	d->509	g->47	k->1	s->88	t->43	
hap	e->1	p->1	
har	 ->1674	"->1	,->14	.->2	:->1	?->1	a->2	d->2	m->24	t->1	
has	 ->1	t->4	
hat	 ->1	e->2	i->1	t->1	
hau	s->1	
hav	 ->2	,->1	a->4	e->27	s->20	
he 	B->1	R->1	c->1	i->1	o->1	
he,	 ->1	
hea	d->1	t->21	
heb	r->1	
hec	k->1	
hed	e->3	r->5	
hee	r->14	
hef	 ->1	e->16	
hei	k->5	
hej	d->2	
hek	t->2	
hel	 ->11	a->105	g->1	h->29	i->1	l->55	m->1	s->47	t->143	
hem	 ->6	.->2	a->1	b->1	f->1	l->15	m->10	s->5	v->1	
hen	 ->7	,->1	.->1	;->1	g->10	n->27	s->2	
hep	h->3	
her	 ->3	"->1	a->2	d->3	e->1	n->10	o->1	r->210	
hes	 ->1	
het	 ->589	!->1	"->3	,->116	.->114	:->1	;->1	?->6	J->1	a->1	e->729	l->36	s->188	t->3	
heu	g->2	
hez	 ->1	
hho	f->1	
hie	l->1	r->4	s->2	
hig	h->1	
hil	l->1	
hin	d->86	g->3	n->2	
hip	 ->1	
hiq	u->1	
his	t->36	
hit	 ->4	,->1	t->58	
hja	m->1	
hjä	l->108	r->27	
hle	r->4	
hne	,->1	r->12	
ho 	f->1	p->1	s->1	v->1	
ho.	 ->1	
hob	b->2	
hoc	-->2	k->4	
hoe	k->1	
hof	e->1	
hok	l->1	
hol	,->1	k->4	m->3	
hom	 ->3	o->4	
hon	 ->29	o->28	
hop	 ->8	,->2	.->3	p->112	
hor	d->2	i->3	m->1	
hos	 ->50	p->1	
hot	 ->11	a->19	b->1	e->8	f->1	
hov	 ->31	,->2	.->3	e->39	s->5	
how	 ->1	
hre	n->7	y->3	
hrk	o->1	
hro	e->14	
hrö	d->1	
hs 	i->1	
ht 	k->1	m->1	o->1	t->1	
ht.	D->1	
hta	l->1	
hte	r->2	
htf	ö->3	
hti	d->1	
hts	.->1	
hu 	o->1	
hud	 ->2	
hug	g->3	
hul	d->1	z->3	
hum	a->6	l->1	ö->2	
hun	 ->1	d->20	
hur	 ->196	.->2	u->14	
hus	 ->6	,->5	.->3	e->6	g->4	h->1	l->1	ö->1	
huv	u->47	
hwa	r->1	
hwe	i->1	
hwi	t->1	
hy 	o->1	
hyc	k->5	
hyg	i->2	
hyl	l->2	
hyp	o->2	
hyr	d->1	e->1	
hys	a->3	e->5	s->5	t->1	
häf	t->2	
häl	e->1	f->3	l->81	s->34	
häm	m->4	n->2	t->8	
hän	;->1	d->79	f->1	g->22	s->80	t->8	v->35	
här	 ->261	,->14	.->10	;->1	?->1	d->6	e->1	i->2	j->2	l->1	m->3	r->4	t->1	v->1	
häs	t->1	
häv	a->7	d->28	e->1	s->2	t->1	
håg	 ->15	.->1	o->2	
hål	 ->2	,->1	:->1	e->1	l->472	
hån	 ->1	a->1	
hår	d->18	e->1	k->1	t->9	
håv	a->1	
hôn	e->1	
hög	 ->21	,->1	a->17	e->32	h->2	l->1	n->3	r->20	s->29	t->17	
höj	a->6	d->12	e->1	n->2	s->1	t->1	
höl	l->18	
hön	a->1	
hör	 ->38	.->1	a->32	d->8	i->19	l->1	n->3	t->27	
hös	t->1	
höv	a->16	d->2	e->99	l->1	s->27	t->3	
hüs	s->4	
i "	g->1	
i -	 ->11	
i 1	5->1	9->15	
i 2	0->13	
i 5	5->1	
i 8	 ->2	
i A	B->1	d->2	f->3	k->2	l->1	m->17	s->1	u->1	v->1	
i B	N->1	e->11	i->5	o->1	r->11	u->1	
i C	E->1	a->1	e->6	u->1	
i D	D->1	a->9	u->4	
i E	C->1	G->8	K->3	M->1	U->15	k->1	t->1	u->173	
i F	a->1	e->1	i->2	o->1	r->11	ö->14	
i G	U->1	a->2	e->2	o->2	r->4	u->2	
i H	a->1	e->14	
i I	C->2	n->2	r->10	s->2	t->6	
i J	o->1	
i K	a->3	f->1	i->3	o->35	y->1	ä->1	ö->1	
i L	a->13	e->1	i->9	o->6	u->5	
i M	a->5	c->1	e->16	i->1	o->3	
i N	e->5	o->1	
i O	L->1	m->1	
i P	P->3	a->3	e->1	o->5	r->1	
i R	a->1	o->1	y->2	
i S	a->3	c->4	e->3	h->4	k->2	r->3	t->15	v->2	y->4	
i T	V->1	a->17	e->1	h->5	i->5	u->7	y->5	
i U	E->1	S->3	r->1	
i V	a->2	e->1	ä->1	
i W	a->4	i->1	
i Y	a->1	
i a	)->1	b->4	c->2	g->3	i->1	k->5	l->96	n->80	r->44	t->78	v->24	
i b	a->6	e->133	i->18	l->7	o->12	r->8	u->9	y->1	ä->2	å->3	ö->44	
i c	e->2	i->1	
i d	a->168	e->560	i->41	o->6	r->3	ä->7	å->9	
i e	f->16	g->15	k->6	m->5	n->161	r->20	t->82	u->6	v->1	x->3	
i f	.->1	a->22	e->10	i->7	j->2	l->7	o->46	r->154	u->6	y->2	ä->4	å->33	ö->234	
i g	a->3	e->42	i->1	j->6	l->5	o->14	r->11	ä->3	å->23	ö->26	
i h	a->291	e->33	i->7	j->3	o->10	u->7	y->1	ä->27	å->12	ö->11	
i i	 ->74	a->1	b->2	c->2	g->2	n->171	t->1	
i j	a->2	o->1	u->26	ä->3	
i k	a->125	e->1	l->8	n->2	o->126	r->39	u->13	v->5	ä->13	
i l	a->21	e->5	i->25	j->5	o->2	y->6	ä->14	å->3	ö->2	
i m	a->12	e->81	i->51	j->1	o->46	y->8	ä->1	å->168	ö->4	
i n	a->7	i->4	o->7	u->24	y->4	ä->25	å->14	ö->3	
i o	b->2	c->100	f->6	k->2	l->6	m->24	n->1	r->9	s->10	t->1	u->1	ö->1	
i p	a->40	e->5	l->12	o->10	r->43	u->2	å->16	
i r	a->13	e->54	i->9	o->1	u->3	ä->16	å->35	ö->16	
i s	a->76	e->42	i->105	j->30	k->107	l->24	m->2	n->11	o->46	p->3	t->133	u->1	v->6	y->61	ä->20	å->19	ö->1	
i t	.->2	a->45	e->2	i->43	j->1	o->7	r->21	v->12	y->11	ä->8	
i u	n->45	p->31	r->3	t->57	
i v	a->49	e->59	i->131	ä->37	å->65	
i y	r->2	t->3	
i z	o->2	
i Ö	V->1	s->37	
i ä	g->5	k->1	m->3	n->20	r->72	v->6	
i å	l->1	r->13	s->1	t->10	
i ö	k->1	n->7	p->1	r->1	s->3	v->22	
i! 	J->2	U->1	
i!H	e->1	
i!J	a->1	
i" 	s->1	
i, 	M->1	b->2	d->6	e->4	f->4	g->1	h->4	i->2	j->3	k->3	l->5	m->11	n->2	o->11	p->1	s->11	t->4	u->2	v->3	ä->4	
i- 	o->10	
i-,	 ->1	
i-g	e->1	
i-i	r->1	
i-r	a->1	
i.(	P->1	
i..	 ->1	.->1	
i.A	l->2	n->1	
i.B	å->1	
i.D	e->11	ä->1	
i.E	f->1	n->1	t->1	u->1	
i.F	o->2	r->1	ö->1	
i.H	a->1	e->1	u->1	ä->1	
i.I	 ->1	
i.J	a->3	
i.K	a->1	u->1	
i.L	i->1	
i.M	a->2	i->1	
i.N	ä->1	
i.S	e->1	o->1	å->1	
i.U	t->1	
i.V	i->5	å->1	
i: 	f->1	
i; 	m->1	
i? 	O->1	
i?.	H->1	
ia 	-->2	B->1	E->1	P->1	R->1	a->4	b->1	d->3	e->1	f->2	h->1	i->2	k->1	m->1	o->4	r->10	s->6	t->3	u->1	v->4	å->1	
ia,	 ->4	
ia-	R->1	
ia.	D->1	Ä->1	
iag	e->1	
iak	t->8	
ial	 ->44	,->3	-->1	.->6	a->78	b->2	d->16	e->4	f->28	i->42	o->31	p->5	t->18	u->1	
ian	 ->1	e->3	o->1	s->8	v->6	
iar	i->21	
ias	 ->4	m->3	
iat	 ->2	.->1	i->84	ä->1	
iba	k->1	n->6	
ibb	i->1	
ibe	d->1	h->11	k->4	l->11	r->32	s->5	t->31	
ibi	 ->1	l->11	
ibl	a->31	i->2	
ibu	t->1	
iby	e->1	
ic 	-->1	B->1	i->1	
ica	l->1	n->1	p->1	
ice	 ->19	.->4	k->2	n->3	r->57	
ich	a->1	e->1	i->1	t->8	y->1	
ici	e->10	n->1	o->1	t->3	
ick	 ->52	,->3	.->5	a->15	b->5	e->48	f->1	l->1	n->1	o->2	p->3	s->5	
icy	,->1	a->1	d->1	f->1	
id 	1->1	7->1	B->3	E->8	G->1	H->1	K->1	L->1	M->1	P->1	a->43	b->19	c->1	d->49	e->26	f->39	g->6	h->22	i->17	j->3	k->17	l->5	m->22	n->10	o->18	p->13	r->7	s->36	t->20	u->16	v->14	y->1	ä->11	å->5	ö->2	
id,	 ->19	
id.	.->1	D->5	E->1	F->1	H->1	J->1	K->1	M->1	N->1	O->1	S->1	T->2	V->1	
id:	 ->1	
ida	 ->64	,->9	.->8	?->1	g->1	k->2	n->61	r->75	s->1	t->14	
idd	 ->5	.->1	a->13	e->2	
ide	 ->1	a->5	e->2	m->1	n->150	o->5	r->98	s->2	
idg	a->38	n->71	
idh	å->4	ö->1	
idi	a->21	g->170	s->31	t->4	ä->1	
idk	a->1	
idl	a->2	i->5	
idm	a->1	
idn	a->1	i->22	
ido	e->1	r->8	s->2	
idp	u->10	
idr	a->108	o->7	
ids	 ->6	,->1	-->1	a->4	b->2	d->4	f->11	g->1	i->2	m->2	o->1	p->17	r->7	s->2	t->1	å->3	ö->1	
idt	a->68	o->2	
idu	a->1	e->8	t->1	
idé	 ->10	,->1	e->8	n->14	
ie 	C->1	R->1	a->1	o->1	
ie,	 ->1	
ie-	 ->1	s->1	
ieb	e->2	ö->1	
iec	k->1	
ied	 ->1	.->1	e->2	
ief	f->6	i->1	u->1	
iek	t->1	
iel	 ->1	a->4	f->1	l->119	s->12	
iem	i->3	
ien	 ->66	,->23	.->13	?->2	d->1	f->1	n->1	s->29	t->46	
iep	r->1	
ier	 ->86	,->16	.->11	a->62	b->2	d->1	i->43	n->44	s->2	
ies	 ->3	k->2	m->1	t->1	
iet	 ->42	"->1	)->4	,->9	.->9	n->3	s->22	y->1	
ieu	r->1	
ieä	g->2	
ifa	l->5	r->2	s->3	
ife	r->6	s->1	
iff	e->5	r->22	
ifi	c->40	e->27	k->32	n->2	q->1	
ifo	l->1	n->2	r->1	
ifr	å->61	
ift	 ->26	!->1	,->2	.->7	:->1	a->16	e->78	i->3	l->8	n->113	s->11	
ifu	l->1	
ifö	r->4	
ig 	-->2	E->1	O->1	a->100	b->36	d->48	e->35	f->124	g->20	h->26	i->79	j->5	k->35	l->16	m->65	n->21	o->102	p->60	r->35	s->76	t->60	u->39	v->29	y->2	ä->14	å->25	ö->10	
ig!	"->1	H->1	
ig"	.->1	
ig,	 ->50	
ig.	 ->2	A->1	B->1	D->10	E->4	G->2	H->2	I->1	J->13	K->1	M->4	N->1	O->3	P->1	S->1	T->1	U->1	V->5	Ä->1	
ig:	 ->3	
ig;	 ->1	
ig?	D->1	H->1	J->1	V->1	
iga	 ->904	,->34	.->31	/->1	;->1	?->1	d->11	n->16	r->170	s->58	t->27	
igd	o->12	
ige	 ->6	.->2	n->571	r->5	s->1	t->12	
igg	a->23	e->87	j->13	ö->21	
igh	 ->1	e->830	t->3	å->2	
igi	e->1	n->2	t->2	ö->4	
igj	o->1	
igl	a->1	i->4	
igm	a->1	
ign	a->15	e->2	o->4	
igo	r->4	t->1	u->1	
igr	a->12	e->1	
igs	e->1	h->1	s->1	t->1	
igt	 ->1085	!->2	,->62	.->77	:->1	;->1	?->1	v->108	
igv	a->1	
igå	 ->1	e->4	n->7	s->1	
igö	r->6	
iha	n->3	
ihe	t->116	
ihj	ä->1	
iho	p->12	
ihä	r->1	
ihå	g->16	
iik	a->3	
iim	p->1	
iin	n->1	t->1	
iis	-->2	
ij-	v->1	
ijs	 ->1	.->1	
ik 	-->2	D->1	J->1	a->5	e->5	f->19	h->5	i->11	k->3	m->13	n->3	o->31	p->5	r->2	s->35	t->1	u->3	v->3	ä->5	å->1	ö->1	
ik!	O->1	
ik"	 ->1	
ik,	 ->35	
ik-	 ->2	
ik.	.->1	B->1	D->11	E->2	F->4	G->1	H->4	I->1	J->1	M->1	R->2	T->1	V->3	Ä->1	
ik:	 ->1	
ik?	H->1	V->1	
ika	 ->251	,->9	-->1	.->8	b->2	d->2	f->1	l->25	n->31	p->8	r->15	s->20	t->30	
ike	 ->56	,->15	.->21	:->1	E->1	F->1	N->1	d->10	l->100	n->168	r->43	s->50	t->18	
ikg	i->2	
ikh	 ->1	-->1	.->2	e->35	
iki	s->54	t->3	
ikl	a->15	e->1	i->6	
ikm	e->2	
ikn	a->22	i->44	
iko	,->1	l->1	m->7	n->3	
ikr	a->7	i->4	o->4	y->2	
iks	 ->1	o->55	t->2	
ikt	 ->123	,->13	.->12	;->1	a->69	e->91	f->1	i->464	l->78	n->55	p->2	s->5	
ikv	ä->9	
ikä	l->37	
il 	-->2	1->1	P->1	e->4	f->2	g->2	i->1	k->1	m->2	n->1	o->1	s->7	u->2	v->1	
il,	 ->2	
il-	 ->2	D->1	R->1	p->1	
il.	 ->1	D->2	J->1	L->1	T->1	
ila	 ->6	g->7	n->1	r->85	t->9	
ilb	e->3	r->1	
ild	 ->21	,->1	.->3	a->67	e->11	n->66	r->6	
ile	d->1	g->6	m->3	n->7	r->1	
ilf	ö->2	
ilh	e->1	
ili	a->1	e->1	g->1	k->1	n->30	s->15	t->35	
ilj	 ->1	a->253	e->26	o->65	t->1	ö->190	
ilk	a->106	e->235	o->1	y->1	ö->2	
ill	 ->2304	!->1	,->25	.->16	:->1	?->3	a->13	b->56	d->13	e->31	f->144	g->49	h->53	i->29	k->79	m->5	n->51	o->6	r->77	s->129	t->11	v->118	ä->197	å->55	
ilm	e->2	ä->1	
ilo	 ->3	,->1	b->1	m->1	s->5	t->4	v->1	
ilp	a->6	r->1	
ilr	e->1	ä->1	
ils	 ->2	e->4	k->8	p->1	t->1	
ilt	 ->133	,->1	i->44	o->1	r->1	
ilu	r->1	
ilv	e->3	r->6	
ilä	g->1	n->1	
ilå	t->1	
ilö	n->1	
ima	 ->5	,->1	.->1	g->2	l->11	n->3	t->15	
imb	u->1	
ime	n->17	r->9	t->1	
imi	b->2	f->1	i->1	k->4	l->2	n->36	r->5	s->7	t->12	x->1	å->1	
iml	i->23	
imm	a->9	e->5	i->6	u->1	
imo	r->1	
imp	l->1	o->10	s->1	u->6	
ims	a->2	b->2	o->1	p->1	r->2	å->1	
imt	 ->3	,->1	
imu	l->13	m->4	s->1	
imy	n->1	
imå	l->1	
imö	g->1	
in 	-->1	1->1	2->1	E->1	F->1	a->19	b->21	d->19	e->22	f->45	g->34	h->23	i->40	k->37	l->5	m->30	n->10	o->42	p->40	r->27	s->53	t->13	u->30	v->14	w->1	y->1	ä->3	å->12	ö->4	
in!	H->1	
in"	,->1	
in,	 ->31	
in-	r->3	
in.	 ->2	A->1	B->1	C->1	D->6	F->2	H->2	I->1	J->3	L->2	M->1	N->1	O->2	S->3	V->5	
in:	 ->1	
in?	P->1	
ina	 ->246	,->1	-->1	.->2	f->2	l->11	n->84	r->2	s->2	t->8	v->1	
inb	a->1	e->12	j->7	l->14	u->1	y->1	
inc	i->203	
ind	 ->1	a->17	e->62	f->4	i->28	r->111	u->113	
ine	 ->6	,->1	f->3	l->4	n->14	r->57	s->9	t->3	z->1	
inf	e->2	i->3	l->12	o->92	r->17	ö->164	
ing	 ->1313	!->1	"->5	)->6	,->196	-->1	.->241	:->4	;->4	?->7	a->645	d->1	e->938	f->22	g->2	i->6	o->4	p->2	r->20	s->990	t->9	å->34	
inh	e->2	o->6	ä->6	
ini	e->17	f->1	m->27	n->1	o->4	p->1	r->1	s->99	t->103	v->1	
inj	e->93	
ink	e->11	l->22	o->16	r->2	t->3	ö->3	
inl	a->6	e->73	i->1	ä->28	å->2	ö->1	
inm	ä->1	
inn	a->155	e->301	i->50	l->2	o->91	s->330	
ino	 ->3	,->2	.->2	m->284	r->25	s->5	t->1	
inp	r->1	
inr	a->13	e->86	i->57	y->1	ä->55	å->1	
ins	 ->21	a->49	b->1	e->43	i->10	k->92	l->6	p->15	t->350	y->13	
int	 ->1	-->1	a->13	e->1777	i->1	l->10	o->7	r->170	y->4	ä->5	
inu	c->1	e->2	s->5	t->16	
inv	a->19	e->25	i->1	o->9	ä->13	å->9	
inz	 ->2	
inä	r->12	
inö	v->1	
io 	S->1	V->4	b->2	f->4	g->3	h->1	l->1	m->9	p->1	s->4	t->1	u->1	ä->1	å->7	
io,	 ->3	
io-	P->4	
io.	J->1	N->1	
io:	 ->1	
io;	 ->1	
iod	 ->23	,->5	.->2	?->1	e->41	i->14	
ioe	k->3	l->1	
iof	e->1	ö->1	
iog	r->1	
iol	a->1	o->6	
ion	 ->323	"->1	)->2	,->48	.->80	:->3	;->1	?->6	a->135	d->2	e->2253	i->5	j->1	s->148	ä->248	
iop	i->3	l->1	
ior	.->1	g->2	i->39	
ios	 ->2	f->1	j->1	ä->2	
iot	 ->2	a->6	e->2	i->1	u->1	
iox	i->7	
ip 	a->3	e->3	f->1	i->7	m->1	o->4	r->1	s->5	ä->4	
ip,	 ->3	
ip.	J->1	S->1	V->2	
ipa	 ->17	,->1	.->2	n->20	r->1	s->1	
ipe	n->105	r->63	s->1	t->3	
ipi	e->8	t->2	
ipl	a->1	i->20	o->11	
ipn	a->1	i->9	
ipo	l->4	t->1	
ipp	a->3	e->2	
ipr	o->7	
ips	 ->1	k->1	
iqu	e->3	i->1	
ir 	E->2	a->10	b->3	d->14	e->10	f->6	g->1	h->3	i->5	j->2	k->1	l->5	m->11	n->5	o->4	r->3	s->13	t->5	u->2	v->4	ä->1	å->1	ö->1	
ir,	 ->2	
ir:	 ->1	
ira	 ->3	,->2	.->1	k->2	r->3	t->1	
ire	 ->1	,->1	-->1	.->1	f->4	g->3	k->257	r->4	
irg	i->5	
iri	g->1	
irk	a->4	e->4	l->2	u->3	
irl	ä->11	
irm	a->1	o->1	
iro	n->2	
irr	a->7	e->1	g->1	i->12	v->1	
irt	a->1	
is 	(->1	-->3	A->1	B->1	G->1	M->1	P->1	W->1	a->27	b->9	d->14	e->9	f->21	g->9	h->16	i->28	j->2	k->8	l->10	m->12	n->3	o->26	p->15	r->4	s->53	t->4	u->8	v->14	ä->21	å->4	ö->3	
is!	 ->1	
is)	 ->1	
is,	 ->22	
is-	J->2	f->1	n->1	p->1	
is.	 ->1	D->4	E->1	F->2	H->1	J->2	M->1	S->2	V->1	Ä->1	
is:	 ->1	
is;	 ->1	
is?	Ä->1	
isa	 ->67	,->8	.->14	?->1	b->1	d->19	k->1	n->8	r->71	s->10	t->82	v->1	
isb	a->1	e->10	ö->7	
isc	a->6	e->1	h->5	i->14	
isd	a->2	i->5	o->1	
ise	 ->1	e->1	k->8	m->3	n->19	r->205	s->2	t->15	
isf	i->3	ö->1	
ish	 ->1	e->3	
isi	o->27	s->70	t->1	ä->1	
isk	 ->344	,->7	-->2	.->11	a->1373	b->8	e->102	f->4	h->6	k->3	n->1	o->91	r->21	t->262	u->143	v->5	
isl	ä->2	
ism	 ->35	,->11	.->20	?->1	e->33	i->2	y->2	
isn	i->15	å->1	
iso	l->7	m->1	n->3	r->5	
isp	e->1	l->1	o->3	
isr	a->20	
iss	 ->43	,->5	.->2	a->155	b->10	e->18	f->7	g->7	h->5	i->1152	k->6	l->20	n->3	o->6	r->2	t->37	u->2	y->1	ä->1	
ist	 ->54	!->1	,->5	.->1	a->146	d->11	e->184	f->9	g->3	h->1	i->92	k->1	l->1	n->2	o->36	p->5	r->53	s->3	y->4	ä->2	å->25	
isu	a->1	e->1	m->1	t->1	
isv	ä->1	
isy	s->1	
isä	k->7	r->4	
it 	-->2	F->1	a->16	b->8	d->13	e->39	f->29	g->2	h->18	i->16	k->5	l->8	m->21	n->8	o->9	p->12	r->3	s->35	t->22	u->25	v->8	ä->1	å->1	ö->7	
it,	 ->8	
it-	a->5	
it.	F->5	I->1	M->2	N->1	P->1	
ita	 ->13	,->1	.->3	d->1	l->35	m->8	n->17	r->13	s->1	t->14	u->1	
itb	o->53	
ite	 ->5	l->7	n->22	r->70	t->311	
ith	ö->1	
iti	a->80	c->1	e->8	k->325	m->21	n->2	o->80	s->260	v->85	ö->12	
itl	a->2	e->7	i->5	ä->1	
itn	i->1	
ito	r->25	
itr	a->5	e->1	o->1	u->2	
its	 ->54	,->4	.->5	
itt	 ->179	,->3	.->1	a->40	e->30	i->61	l->1	n->7	r->6	s->2	é->59	
itu	 ->20	a->129	d->1	e->1	l->2	m->1	t->158	
ity	d->5	
itz	 ->1	.->1	
itä	r->7	
ium	 ->13	!->1	,->4	.->9	
iut	s->1	
iv 	(->1	-->3	9->8	E->1	a->7	b->3	d->4	e->7	f->18	g->1	h->8	i->14	k->12	l->8	m->6	o->32	p->8	r->4	s->49	t->17	u->3	v->6	ä->6	å->2	ö->1	
iv,	 ->27	
iv.	 ->1	.->2	A->2	B->1	D->6	E->1	F->4	I->3	L->1	M->2	O->1	R->1	S->1	V->2	Y->1	
iv:	 ->2	
iv;	 ->1	
iv?	F->1	N->1	
iva	 ->146	,->4	.->3	d->1	n->24	r->63	s->10	t->26	v->7	
ivb	e->1	o->1	
ive	 ->32	l->38	n->26	r->51	s->1	t->159	
ivf	ö->4	
ivi	d->14	e->2	l->38	s->4	t->88	
ivk	r->3	
ivl	a->10	i->5	
ivn	a->9	i->11	
ivr	a->1	i->1	ä->4	
ivs	 ->13	,->1	.->1	c->3	d->2	k->6	m->91	u->1	v->1	
ivt	 ->111	,->7	.->7	
ivä	g->3	
ivå	 ->46	,->13	.->21	;->1	?->1	e->14	g->3	n->12	
iwa	n->1	
ix.	D->1	
ixa	s->5	
ixe	n->1	
ixt	r->1	
iz 	e->1	f->2	s->1	
iz,	 ->2	
iz-	k->1	
izi	s->5	
iäk	e->1	
iär	,->1	a->1	e->4	m->10	p->1	
iål	d->1	
iåt	e->1	
ièr	e->1	
ié 	u->1	
iös	 ->4	,->1	a->13	t->6	
j 1	9->3	
j 2	0->1	
j L	i->1	
j a	n->1	t->1	v->1	
j b	e->2	o->1	
j f	ö->3	
j i	 ->1	
j k	o->1	
j l	å->1	ö->1	
j m	o->1	
j n	ä->1	
j o	m->1	
j t	i->1	
j ä	r->1	
j ö	v->1	
j, 	b->2	d->1	h->1	j->1	m->2	n->1	o->2	s->2	ä->1	
j-v	a->1	
j.(	A->1	
j.D	e->1	
j.E	x->1	
j.I	 ->1	
j.J	a->1	
j.R	å->1	
j.T	o->1	
j.V	i->1	
ja 	-->3	D->1	F->1	H->2	J->1	M->1	a->32	b->18	c->2	d->48	e->27	f->39	g->19	h->14	i->6	k->15	l->7	m->41	n->4	o->17	p->13	r->7	s->47	t->35	u->23	v->11	y->2	Ö->1	å->6	ö->1	
ja,	 ->11	
ja.	.->1	H->1	J->2	K->1	M->1	T->1	V->1	
jad	e->18	
jag	 ->1069	,->15	.->2	a->2	
jak	t->24	
jal	a->2	i->5	
jam	o->1	
jan	 ->32	,->3	a->1	d->77	u->16	
jap	a->1	
jar	 ->39	.->2	b->1	d->15	e->8	n->6	
jas	 ->25	,->4	.->6	
jat	 ->16	.->2	a->1	s->4	
jd 	-->1	a->19	g->1	m->1	p->1	s->1	u->1	
jd.	J->1	
jda	 ->7	,->3	s->1	t->1	
jde	 ->6	n->1	r->19	s->2	
jdo	s->1	
jdp	u->2	
jdr	i->1	
jds	k->2	
jdå	t->1	
je 	(->1	-->1	1->1	B->1	E->2	a->5	b->5	d->11	e->7	f->19	g->8	h->2	i->3	k->3	l->33	m->20	n->1	o->5	p->6	r->5	s->11	v->4	ä->1	å->11	ö->3	
je,	 ->4	
je-	 ->1	
je.	G->1	J->1	
je:	 ->1	
jeb	e->1	o->4	ä->10	
jed	e->6	o->1	
jef	a->1	ö->2	
jei	n->3	
jej	o->3	
jek	o->2	t->68	
jel	a->6	i->1	s->4	
jem	ä->1	
jen	 ->3	.->1	
jer	 ->82	"->1	,->10	.->4	:->1	a->16	n->35	
jes	k->1	t->1	
jet	 ->2	a->9	r->2	t->2	
jeu	t->2	
jev	ä->3	
jeå	t->1	
jfl	ö->1	
jik	i->5	
jka	n->1	
jko	n->2	t->1	
jli	g->309	
jni	n->19	
job	b->4	
joc	k->2	
jol	 ->2	,->1	.->1	
jon	 ->1	e->63	i->1	t->1	
jor	 ->1	.->1	d->113	i->42	n->1	t->104	
jos	 ->1	
jou	r->3	
jov	i->17	
js 	a->1	k->1	o->1	t->1	u->2	
js,	 ->1	
js.	(->1	
jsm	å->2	
jt 	i->1	o->1	s->1	u->1	v->1	
jts	 ->3	,->1	
ju 	E->1	M->1	a->11	b->2	d->5	e->2	f->2	g->1	h->1	i->12	l->1	m->7	o->8	p->4	r->3	s->7	t->1	u->1	v->1	ä->7	
ju,	 ->3	
jua	d->1	
jub	l->1	
jud	a->23	d->1	e->18	i->6	l->1	n->3	
jug	e->1	o->4	
juk	.->1	a->2	d->1	f->1	h->7	n->2	v->3	
jul	 ->1	f->1	i->10	k->1	
jun	d->4	g->3	i->12	k->10	
jup	 ->1	a->13	e->5	g->7	n->5	s->1	t->7	
jur	 ->2	,->2	-->2	.->2	a->1	e->2	f->4	i->47	l->2	
jus	 ->1	.->1	e->8	t->111	
jut	a->13	e->8	i->5	n->1	s->5	t->2	v->1	
juv	e->2	
jäl	 ->1	,->1	.->2	e->2	p->107	t->3	v->170	
jäm	f->16	k->2	l->13	n->11	s->24	t->3	v->2	
jän	a->21	s->123	t->29	
jär	a->1	d->11	e->1	n->19	t->27	v->7	
jät	t->21	
jäv	u->2	
jö 	f->2	i->1	k->1	m->1	s->2	v->1	
jö!	D->1	
jö,	 ->11	
jö-	 ->2	
jö.	D->3	M->1	U->1	V->1	
jöa	n->3	v->1	
jöb	e->3	r->1	
jöd	 ->1	e->1	i->1	s->1	
jöe	r->4	
jöf	a->10	r->4	ö->4	
jöi	n->1	
jök	a->11	o->6	r->8	v->1	
jöl	a->1	
jöm	i->1	ä->13	å->3	
jön	 ->15	!->1	,->9	.->11	k->4	o->2	s->2	
jöo	m->4	v->1	
jöp	e->1	o->8	r->4	å->1	
jör	 ->2	å->1	ö->2	
jös	e->1	i->1	k->15	s->4	t->5	y->6	
jöt	r->1	
jöu	t->1	
jöv	ä->10	
k -	 ->6	
k D	e->1	
k J	ö->1	
k K	i->1	
k T	V->1	
k a	 ->1	g->1	l->9	n->7	r->3	s->1	t->24	v->13	
k b	a->7	e->12	i->4	l->2	o->2	r->1	y->3	ö->1	
k c	i->2	
k d	a->2	e->14	i->7	
k e	f->3	g->1	j->1	k->1	l->4	m->1	n->7	r->1	t->2	
k f	e->1	i->4	l->2	o->3	r->12	y->1	å->3	ö->50	
k g	a->1	e->5	j->1	l->1	r->4	ä->3	å->2	
k h	a->17	e->1	j->2	o->3	u->2	ä->2	ö->3	
k i	 ->31	d->1	m->1	n->29	
k j	a->4	o->1	u->4	ä->2	
k k	a->15	l->2	o->30	u->5	v->1	ä->2	
k l	a->5	e->5	i->5	o->1	y->1	ä->3	ö->1	
k m	a->6	e->17	i->5	o->7	y->5	å->6	ö->2	
k n	a->3	e->1	i->14	j->1	u->1	y->1	ä->5	å->3	
k o	c->74	f->4	j->1	m->11	p->1	r->1	s->3	
k p	a->3	e->2	l->2	o->20	r->5	u->1	å->13	
k r	a->3	e->11	i->1	o->5	ä->1	å->1	ö->2	
k s	a->3	e->3	i->5	j->1	k->8	m->1	n->1	o->60	t->16	v->1	y->6	ä->3	å->17	
k t	e->1	i->30	r->3	v->2	y->1	ä->1	
k u	n->8	p->6	r->1	t->17	
k v	a->11	e->1	i->19	ä->4	
k ä	n->2	r->12	
k å	k->13	t->3	
k ö	v->5	
k!A	n->1	
k!O	m->1	
k" 	-->1	f->1	o->1	
k, 	1->1	R->1	a->1	b->1	d->13	e->5	f->10	g->2	h->8	i->6	k->6	m->9	n->4	o->3	s->11	t->13	u->1	v->5	ä->1	
k- 	e->1	o->2	
k-b	r->1	
k-d	a->1	
k-f	r->1	
k-i	s->1	
k-p	o->1	
k-s	k->1	
k. 	D->1	J->1	M->1	a->1	i->1	s->2	
k..	(->1	
k.A	t->2	v->1	
k.B	e->1	y->1	
k.D	e->20	ä->1	å->2	
k.E	n->1	t->1	u->1	
k.F	a->1	r->4	ö->1	
k.G	e->1	
k.H	a->2	e->7	i->1	u->1	ä->1	
k.I	 ->3	n->1	
k.J	a->7	
k.K	i->1	o->1	
k.M	e->3	
k.N	i->1	
k.O	c->1	m->1	
k.R	e->1	i->1	
k.S	y->1	
k.T	a->1	r->1	v->1	y->1	
k.V	a->1	i->9	
k.Ä	v->2	
k: 	g->1	v->1	
k?H	e->1	
k?N	e->1	
k?R	e->1	
k?V	a->1	
ka 	"->1	-->4	1->1	2->1	A->1	B->1	E->6	F->2	G->2	K->3	L->1	P->5	S->1	T->1	a->105	b->88	c->3	d->95	e->56	f->198	g->66	h->48	i->121	j->6	k->202	l->56	m->143	n->31	o->183	p->129	r->138	s->204	t->67	u->298	v->85	ä->22	å->32	ö->12	
ka"	,->1	
ka,	 ->44	
ka-	o->1	
ka.	(->1	B->1	D->4	E->4	F->1	H->2	I->3	J->5	L->1	M->2	O->1	P->2	R->1	T->1	V->5	Å->1	
ka:	 ->2	
ka?	"->1	I->1	
kab	a->1	e->3	i->3	
kad	 ->38	.->1	a->27	e->60	i->1	l->10	m->3	o->26	r->3	
kaf	f->26	r->1	
kag	å->4	
kak	a->2	
kal	 ->10	:->1	a->43	d->1	e->1	i->12	l->716	p->1	t->7	v->1	y->1	
kam	 ->2	!->1	,->1	l->2	m->61	p->31	r->1	
kan	 ->862	,->6	.->7	a->11	d->384	e->17	i->11	o->1	s->71	t->7	
kao	s->2	
kap	 ->75	"->3	,->16	.->17	:->1	a->186	e->244	i->25	l->37	p->6	r->1	s->92	t->2	
kar	 ->177	,->8	.->8	:->1	a->18	e->58	g->1	k->2	l->6	n->52	p->2	r->2	s->1	t->18	
kas	 ->84	!->1	,->10	.->10	k->1	m->1	s->3	t->44	u->3	å->4	
kat	 ->56	,->8	.->7	a->92	e->10	i->18	o->12	s->32	t->66	
kav	i->4	
kay	 ->3	,->3	.->1	D->1	b->1	s->2	
kba	r->12	
kbe	d->4	s->4	
kbi	l->1	
kbo	r->1	
kbä	r->1	
kda	m->1	
kde	l->8	
kdo	m->1	
kdö	r->1	
ke 	(->1	-->4	I->1	a->6	b->7	d->6	e->9	f->9	g->5	h->4	i->21	k->12	l->8	m->8	n->4	o->20	p->48	r->3	s->14	t->14	u->7	v->8	ä->11	ö->1	
ke!	Ä->1	
ke)	 ->2	
ke,	 ->24	
ke-	a->2	d->3	f->1	m->1	s->12	
ke.	 ->1	-->1	.->2	D->6	F->4	H->1	I->1	J->2	M->2	N->1	O->1	V->4	Ö->1	
ke:	 ->1	
keE	n->1	
keF	r->1	
keN	ä->1	
keb	a->1	
ked	 ->3	.->1	a->4	e->7	j->4	o->10	
kef	r->1	ö->1	
keg	å->1	
kek	v->1	
kel	 ->109	,->4	.->4	:->2	f->3	m->1	n->8	p->1	r->2	s->11	t->29	v->2	
kem	e->1	i->7	å->3	ö->4	
ken	 ->279	,->30	.->38	:->3	?->3	H->1	s->39	
keo	m->2	
kep	o->2	p->8	s->1	t->8	
ker	 ->297	,->13	.->14	:->2	a->28	e->1	h->235	i->10	l->15	n->33	s->26	t->30	ä->2	
kes	 ->26	-->4	a->1	e->2	f->5	h->4	i->1	k->2	l->4	m->10	p->3	t->1	u->7	v->1	
ket	 ->699	!->1	,->35	.->12	:->1	;->3	?->1	e->3	i->2	m->1	r->3	s->14	t->15	
kev	a->2	
kfa	k->1	r->7	
kfo	r->1	
kfr	i->2	o->1	
kfy	l->1	
kfö	r->11	
kgi	l->2	
kgr	u->33	
kh 	h->1	
kh-	a->1	
kh.	D->1	F->1	
kha	n->6	
khe	e->14	t->41	
kho	l->3	
khu	s->7	
khä	l->9	
ki 	L->2	
ki.	D->1	
kic	k->17	
kid	n->1	
kie	n->3	t->35	
kif	t->6	
kig	 ->1	t->4	
kil	d->62	j->21	l->47	o->5	t->130	
kin	 ->4	.->1	e->12	g->4	l->1	
kip	a->3	n->9	
kir	e->1	
kis	 ->3	!->1	b->1	k->67	s->4	t->12	
kit	 ->4	i->2	s->1	
kiv	 ->1	e->1	
kju	t->31	
kka	p->1	
kki	 ->2	
kko	m->2	
kku	n->2	y->2	
kkö	y->1	
kl.	 ->20	1->1	
kla	 ->41	.->1	d->12	g->94	m->3	n->44	p->2	r->284	s->47	t->7	u->6	v->1	
kle	d->1	r->5	t->1	
kli	b->1	e->1	g->385	m->14	n->177	
klo	a->1	c->2	k->7	
klu	d->4	k->1	s->20	
kly	f->5	v->1	
klä	g->1	
klö	s->1	
km 	l->1	m->1	
km,	 ->1	
km.	T->1	
kme	n->2	t->2	
kmo	d->1	
kna	 ->13	,->1	.->1	d->204	n->20	p->16	r->38	s->30	t->19	
kne	e->1	l->1	s->1	
kni	k->13	n->349	p->4	s->36	v->1	
kno	l->3	w->1	
knu	s->1	t->7	
kny	t->9	
knä	c->2	
ko 	C->5	
ko,	 ->1	
ko.	T->1	
koa	l->14	
kod	 ->7	e->6	i->2	
koe	f->1	
kof	f->1	i->2	ö->2	
kog	 ->3	a->10	e->5	r->1	s->20	å->1	
koh	a->3	e->1	o->1	
kok	a->1	o->1	
kol	-->1	a->6	d->5	e->1	i->4	l->234	o->21	
kom	 ->48	,->1	.->1	a->1	b->1	l->9	m->2160	n->45	p->90	r->16	s->18	
kon	 ->1	a->2	c->42	f->193	g->1	j->1	k->329	o->286	s->238	t->224	v->27	
koo	p->1	
kop	 ->1	,->3	i->2	o->5	p->6	
kor	 ->96	,->12	.->10	a->1	d->2	e->22	l->2	n->34	r->39	s->15	t->98	
kos	a->1	l->1	t->116	y->4	
kot	i->7	t->172	
kou	r->1	
kov	 ->2	e->1	
kpa	r->10	
kpr	o->4	
kra	 ->37	d->3	f->149	n->1	r->10	s->10	t->171	v->91	
kre	a->3	d->2	g->1	n->2	p->3	r->1	t->85	v->8	
kri	d->21	f->22	g->23	k->44	m->27	n->55	s->35	t->70	v->61	
kro	a->1	e->5	f->2	k->2	m->3	n->1	p->1	s->2	t->27	v->15	
kry	.->1	g->1	p->5	s->1	t->1	
krä	c->9	d->1	f->30	k->1	m->5	n->29	p->1	t->1	v->139	
krå	n->2	
krö	n->1	
ks 	a->4	b->2	d->3	e->1	f->1	g->1	i->1	m->3	n->1	o->6	p->2	r->1	s->4	t->3	u->2	v->3	ö->1	
ks,	 ->1	
ks.	D->1	O->1	P->1	U->1	V->1	
ks;	 ->1	
ksa	k->1	m->129	n->1	
ksb	o->1	å->1	
ksc	e->1	h->1	
ksd	r->3	
kse	k->2	
ksf	a->2	o->1	r->1	
ksi	l->3	
ksk	ö->1	
ksl	o->1	u->1	
kso	d->1	m->57	n->2	
ksp	o->6	r->3	
ksr	e->2	i->2	
kss	e->5	y->1	
kst	a->2	y->1	ä->22	
ksv	a->1	
ksw	a->1	
ksä	g->1	
kså	 ->572	,->10	.->5	
ksö	d->1	
kt 	(->2	-->5	1->3	2->3	4->2	5->1	6->1	7->1	D->1	E->6	F->2	K->1	M->1	a->64	b->39	c->2	d->20	e->21	f->81	g->13	h->27	i->42	j->1	k->29	l->11	m->43	n->8	o->59	p->52	r->8	s->114	t->20	u->20	v->38	ä->25	å->1	ö->6	
kt!	N->1	
kt"	,->1	
kt,	 ->47	
kt.	 ->1	(->1	A->2	B->4	D->20	F->2	G->1	H->1	I->3	J->6	K->1	M->7	N->2	O->4	P->1	R->1	S->2	T->2	U->1	V->6	Å->1	
kt:	 ->4	
kt;	 ->2	
kt?	E->1	T->1	U->1	
kta	 ->90	,->2	.->4	b->3	d->24	g->1	i->2	k->3	l->1	n->18	r->44	s->19	t->25	
ktb	a->5	e->2	
ktd	e->1	i->1	
kte	 ->31	,->3	.->2	l->13	n->195	r->230	s->5	t->16	
ktf	a->1	ö->2	
kth	a->1	e->1	å->1	
kti	e->3	g->491	k->12	n->16	o->124	s->74	v->415	
ktk	o->1	
ktl	i->92	ö->3	
ktm	e->2	i->1	
ktn	i->55	
kto	b->8	r->137	
ktp	u->2	
ktr	a->1	i->1	o->9	u->2	
kts	 ->11	!->1	a->3	b->1	f->4	m->1	p->2	
ktt	a->8	
ktu	a->1	e->34	m->68	r->154	
kty	g->8	r->1	
ktä	r->9	
ktö	r->23	
kub	i->2	
kug	g->3	
kul	a->7	d->3	e->2	i->1	l->505	o->1	t->121	ä->1	
kum	e->46	u->2	
kun	d->33	g->15	n->261	s->17	
kup	a->2	e->3	p->1	
kur	 ->1	a->1	r->285	s->17	
kus	 ->2	.->1	e->3	s->61	t->31	
kut	a->7	e->78	
kuu	m->2	
kuy	u->2	
kva	,->1	l->53	n->7	r->35	t->6	
kve	n->62	s->3	
kvi	c->3	d->3	n->59	s->1	
kvo	t->16	
kvä	l->14	m->16	r->18	v->2	
kvå	r->3	
ky 	f->1	
kyd	d->109	
kyf	a->1	
kyh	ö->1	
kyl	a->2	d->29	i->1	l->5	
kym	m->6	r->10	t->1	
kyn	d->15	
kyr	k->1	
kyv	ä->1	
käl	 ->35	,->1	.->4	e->12	i->1	l->47	
käm	d->1	m->2	n->1	p->46	t->1	
kän	d->40	k->2	n->151	s->43	t->29	
kär	 ->2	a->53	e->1	l->3	n->56	p->11	s->1	
kåd	a->3	l->6	n->1	
kål	e->1	
kår	,->1	
kåt	 ->2	s->1	
kök	s->1	
köl	 ->1	,->1	a->1	d->2	
kön	e->3	h->1	s->6	
köp	 ->2	a->4	e->1	k->1	s->2	t->1	
kör	 ->1	.->1	a->4	d->3	n->2	s->3	t->3	
köt	 ->2	a->7	e->1	s->8	t->11	
köv	l->1	
köy	 ->1	
l "	M->1	
l (	B->1	k->2	
l -	 ->13	,->1	
l 1	 ->4	,->2	-->11	.->1	0->2	1->1	2->2	3->5	4->1	5->4	6->1	9->4	
l 2	 ->6	,->3	-->3	.->3	2->1	5->5	8->5	9->2	
l 3	 ->1	.->2	0->2	3->2	7->2	9->1	
l 4	 ->6	.->1	2->1	8->2	
l 5	 ->1	.->1	0->3	2->1	6->1	b->2	
l 6	 ->9	,->1	.->1	2->1	7->1	
l 7	 ->7	,->2	0->1	5->1	7->1	
l 8	1->10	2->2	3->1	5->1	7->2	8->2	
l 9	 ->1	.->1	1->1	4->3	5->1	
l A	l->1	
l B	a->2	o->2	r->2	
l C	h->1	o->2	
l D	e->1	i->1	
l E	G->3	U->6	f->1	u->25	
l F	r->3	ö->4	
l G	e->1	r->1	
l H	e->1	i->1	
l I	n->2	r->1	
l K	a->3	i->3	o->10	u->1	
l L	o->2	
l M	c->1	i->1	o->2	
l N	i->2	y->1	
l O	L->1	
l P	P->1	a->3	e->1	o->1	u->1	
l R	a->1	i->1	
l S	c->1	h->1	o->3	t->2	y->1	
l T	h->1	i->1	r->1	y->2	
l U	l->1	
l V	e->1	
l W	a->2	i->1	u->1	
l a	b->1	c->1	g->1	l->37	n->38	p->1	r->14	t->300	v->152	
l b	a->17	e->94	i->13	l->26	o->6	r->6	u->1	y->2	ä->6	å->2	ö->14	
l c	a->1	e->1	i->2	o->1	
l d	a->1	e->299	i->28	o->4	r->4	u->3	ä->17	å->4	
l e	f->6	g->3	k->3	l->7	m->3	n->117	r->15	t->32	u->3	x->46	
l f	a->14	e->3	i->8	l->3	o->13	r->56	u->14	y->2	ä->2	å->13	ö->222	
l g	a->8	e->38	i->1	l->1	o->10	r->21	ä->15	å->13	ö->25	
l h	a->94	e->12	i->5	j->6	o->2	u->6	y->1	ä->9	å->2	ö->7	
l i	 ->78	c->1	d->1	n->110	s->1	
l j	a->109	o->1	u->6	ä->2	
l k	a->19	l->4	n->1	o->88	r->6	u->58	v->6	ä->3	ö->1	
l l	a->3	e->6	i->14	u->1	y->7	ä->16	å->3	ö->3	
l m	a->23	e->63	i->26	o->7	u->1	y->8	ä->2	å->16	ö->6	
l n	a->14	i->16	o->2	u->4	y->13	ä->18	å->12	ö->2	
l o	a->1	c->154	e->1	f->3	i->1	j->1	l->6	m->49	p->1	r->9	s->4	ä->2	
l p	a->11	e->11	i->1	l->5	o->8	r->24	u->2	å->46	
l r	a->4	e->40	i->7	o->4	y->1	ä->23	å->20	ö->4	
l s	a->25	e->19	i->40	j->7	k->47	l->17	m->2	n->1	o->112	p->4	t->81	u->6	v->4	y->7	ä->57	å->6	ö->1	
l t	a->53	e->3	i->45	o->3	r->18	u->1	v->8	y->3	ä->2	
l u	-->1	n->19	p->24	r->6	t->57	
l v	a->60	e->24	i->71	o->6	ä->7	å->16	
l y	r->2	t->3	
l Ö	s->1	
l ä	g->1	n->23	r->41	v->6	
l å	k->2	r->2	s->3	t->22	
l ö	k->6	n->1	p->3	s->1	v->20	
l! 	I->1	J->1	
l!H	e->1	ä->1	
l!J	a->1	
l!M	e->1	
l!T	i->1	
l" 	m->1	o->1	
l",	 ->2	
l".	I->1	
l'e	a->1	
l, 	A->1	R->1	T->1	a->8	b->1	d->9	e->9	f->8	g->2	h->6	i->8	j->3	k->5	l->3	m->20	n->9	o->32	p->3	r->3	s->23	t->4	u->5	v->11	ä->4	å->3	ö->1	
l- 	o->18	
l-2	-->1	
l-D	e->1	
l-F	i->3	
l-H	e->1	
l-I	)->1	I->1	
l-R	o->1	
l-S	h->6	y->1	
l-f	ö->1	
l-p	r->1	
l-s	o->2	
l. 	1->17	2->3	D->1	E->1	J->1	o->1	
l.1	2->1	
l.A	l->1	n->1	v->1	
l.B	e->1	i->1	ä->1	
l.D	e->44	ä->3	
l.E	U->1	f->1	n->3	t->3	u->2	
l.F	i->2	r->5	ö->8	
l.G	e->1	
l.H	a->1	e->8	u->1	ä->1	
l.I	 ->8	n->2	
l.J	a->22	
l.K	a->1	o->4	u->1	ä->1	
l.L	y->1	
l.M	a->1	e->9	i->1	å->1	
l.N	ä->4	
l.O	m->1	r->1	
l.P	e->1	r->1	å->1	
l.R	e->1	
l.S	a->4	c->1	j->1	m->1	o->1	t->1	å->4	
l.T	a->1	r->1	v->1	ä->1	
l.U	t->1	
l.V	i->23	o->1	å->1	
l.a	.->27	
l.Ä	n->2	r->1	v->1	
l: 	"->1	E->1	F->1	O->1	U->1	V->2	a->1	d->1	e->1	j->1	p->1	
l; 	a->1	f->1	i->1	
l?.	 ->1	
l?D	a->1	
l?E	l->1	
l?H	u->1	
l?J	a->2	
l?K	o->1	
lFi	n->1	
la 	-->2	9->1	A->1	B->1	E->24	F->1	H->1	K->2	L->1	M->1	P->1	S->1	U->1	a->87	b->61	d->158	e->87	f->128	g->26	h->39	i->58	j->7	k->74	l->30	m->116	n->24	o->159	p->75	r->63	s->178	t->53	u->54	v->50	ä->9	å->16	ö->8	
la!	H->1	
la"	 ->2	.->2	;->1	
la,	 ->24	
la.	B->1	D->12	H->2	I->1	J->3	K->1	M->2	N->1	S->1	V->4	Ö->1	
la:	F->1	
la?	A->1	D->3	
laa	m->1	
lab	o->3	
lac	e->17	i->15	
lad	 ->30	,->1	a->4	d->3	e->100	
laf	r->1	
lag	 ->347	,->40	.->44	;->1	?->3	a->97	d->12	e->159	f->5	g->28	i->16	l->18	n->33	o->10	r->3	s->146	t->75	
lai	 ->7	
lak	 ->1	t->25	
lam	 ->3	,->1	e->602	o->2	p->1	s->4	t->1	
lan	 ->226	"->2	,->6	.->10	:->1	?->1	N->1	a->4	c->1	d->642	e->101	g->8	h->4	k->4	l->1	n->1	s->51	t->13	ö->19	
lap	p->8	
lar	 ->377	,->30	.->32	:->1	;->1	?->2	a->83	b->1	e->57	f->2	g->17	h->12	i->27	l->5	m->4	n->62	s->3	t->99	v->1	y->1	
las	 ->96	,->8	.->8	:->1	h->1	i->6	p->1	s->22	t->29	
lat	 ->58	,->5	.->3	e->14	h->4	i->34	l->1	o->3	s->65	t->1	
lau	d->1	s->6	t->2	
lav	a->4	e->1	i->1	t->1	
law	,->1	.->1	
lay	a->1	e->2	
lba	c->1	k->52	n->19	r->47	
lbe	f->2	l->1	r->2	s->8	
lbi	l->1	
lbl	o->1	
lbo	r->3	
lbr	a->1	i->5	o->1	
lbu	n->15	
lby	r->1	
ld 	W->1	a->3	b->4	f->6	i->4	k->4	m->3	o->2	p->5	r->3	s->1	t->3	u->2	ä->1	å->1	
ld,	 ->10	
ld.	D->1	F->1	J->2	N->1	
lda	 ->68	,->5	.->6	?->1	d->3	g->1	n->6	r->6	s->10	t->5	
ldb	e->2	
lde	 ->25	,->1	.->1	l->42	m->16	n->46	r->15	s->12	t->2	z->3	
ldg	r->1	
ldh	e->23	
ldi	g->54	o->5	r->17	s->1	
ldj	u->1	
ldn	i->66	
ldo	m->1	
ldr	a->10	e->7	i->32	
lds	a->3	d->1	e->1	f->1	h->6	k->6	l->1	m->1	n->1	o->1	u->1	
ldt	a->2	
le 	-->1	E->3	K->1	a->25	b->21	d->41	e->8	f->31	g->17	h->23	i->26	j->44	k->66	l->5	m->5	n->4	o->14	p->7	r->5	s->30	t->14	u->16	v->123	ä->4	å->2	ö->2	
le,	 ->3	
le-	d->2	
le.	J->1	V->1	
led	 ->2	a->246	d->23	e->84	i->1	n->74	s->9	
lef	a->1	o->1	
leg	a->105	e->133	i->26	o->4	
leh	a->3	
lei	d->2	
lej	d->2	
lek	a->1	e->3	o->7	s->1	t->33	
lel	e->3	l->5	s->9	
lem	 ->79	,->14	.->23	:->1	;->2	?->1	a->5	e->85	i->1	l->1	m->17	o->3	s->323	
len	 ->174	"->3	,->32	.->38	?->1	F->2	a->10	n->7	s->12	t->1	u->5	Ä->1	ä->1	
leo	t->1	
ler	 ->1029	,->20	-->1	.->22	;->1	?->1	a->197	e->7	i->30	k->3	m->1	n->52	s->6	t->73	å->12	
les	 ->38	.->2	;->1	a->7	e->1	k->1	m->2	n->4	t->47	ä->2	
let	 ->227	!->1	,->31	.->38	:->1	a->1	s->6	t->37	
leu	m->1	r->3	
lev	 ->15	a->31	d->2	e->23	i->1	n->12	s->3	t->4	
lew	o->2	
lex	 ->1	.->1	a->3	i->27	t->1	
lez	 ->1	
lf 	H->2	
lf-	M->2	
lfa	b->1	
lfe	d->1	n->4	r->1	
lfi	n->1	
lfk	r->1	
lfo	g->6	n->15	r->3	
lfr	a->3	e->27	i->2	å->9	
lfs	t->3	
lft	e->4	
lfu	n->3	
lfä	l->97	r->9	
lfå	n->4	
lfö	l->3	r->39	
lga	d->1	r->1	
lge	m->1	n->1	r->1	
lgi	e->9	s->8	v->1	
lgj	o->1	
lgo	d->1	
lgr	i->2	u->2	
lgä	n->21	
lgå	n->25	v->1	
lgö	r->2	
lha	n->43	v->4	
lhe	l->1	t->24	
lhj	ä->8	
lho	e->1	
lhö	r->8	
li 	-->1	1->4	2->3	a->11	b->5	d->5	e->31	f->13	g->1	h->2	j->1	k->4	l->4	m->21	n->5	o->3	p->3	r->1	s->9	t->3	u->1	v->4	ä->1	ö->2	
li!	J->1	
li,	 ->3	
li.	U->1	
lia	-->1	n->7	
lib	a->2	b->1	e->29	i->1	
lic	 ->1	a->1	e->17	i->4	k->25	y->4	
lid	a->33	e->10	i->3	
lie	n->38	r->6	s->1	
lif	i->15	
lig	 ->267	!->1	,->13	.->15	:->2	?->2	a->771	e->481	g->142	h->335	i->5	s->1	t->831	
lih	o->1	
lik	 ->4	.->1	:->1	a->186	e->15	g->2	h->35	n->65	r->3	s->49	t->57	v->8	
lil	l->6	
lim	a->17	e->1	i->6	s->1	
lin	 ->12	,->3	.->2	a->1	b->1	d->63	e->4	f->1	g->440	i->2	j->93	k->2	o->1	r->6	s->1	t->3	ä->4	
lio	t->2	
lip	p->2	
lir	 ->112	,->2	:->1	a->1	t->1	
lis	 ->1	,->1	.->1	;->1	a->3	e->85	i->4	k->26	m->16	s->3	t->137	v->1	
lit	 ->22	,->1	a->27	e->137	i->547	l->5	s->6	t->12	ä->6	
liv	 ->9	,->4	.->5	a->22	e->25	i->27	s->101	
lix	t->1	
lj 	L->1	o->1	ö->1	
lj,	 ->2	
lj.	V->1	
lja	 ->228	,->5	.->4	d->3	k->18	n->60	r->35	s->16	t->8	
ljd	 ->18	.->1	e->21	r->1	s->2	å->1	
lje	-->1	b->15	d->1	f->3	i->3	j->3	k->2	l->4	m->1	r->63	s->2	t->11	u->2	å->1	
ljf	l->1	
ljk	o->2	
ljn	i->13	
ljo	n->65	
ljs	 ->4	,->1	
ljt	 ->3	s->2	
lju	d->3	g->1	s->10	
ljö	 ->8	!->1	,->11	-->2	.->6	a->4	b->4	d->2	e->4	f->10	i->1	k->26	l->1	m->15	n->39	o->5	p->14	r->3	s->24	u->1	v->9	
lk 	a->1	b->2	h->1	i->2	o->2	r->1	s->3	t->1	u->1	
lk,	 ->1	
lk.	A->1	D->1	M->1	O->1	V->4	
lka	 ->108	d->1	n->7	r->5	s->10	t->1	
lke	m->1	n->61	s->1	t->194	
lkf	r->1	
lkg	r->2	
lkh	ä->9	
lkl	a->3	i->2	
lkn	i->57	
lko	h->1	m->67	n->2	r->65	
lkp	a->10	
lkr	e->8	i->1	ä->1	
lks	 ->3	t->1	w->1	ä->1	
lku	r->1	
lkv	a->2	o->1	
lky	r->1	
lkä	n->12	
lkö	p->2	
ll 	"->1	-->3	1->5	2->4	3->2	4->1	5->1	7->4	8->2	9->4	A->1	B->5	C->2	D->1	E->35	F->7	G->2	I->1	K->15	L->2	M->4	N->2	O->1	P->5	R->1	S->7	T->5	V->1	W->4	a->397	b->161	c->4	d->337	e->220	f->255	g->119	h->122	i->119	j->117	k->165	l->44	m->104	n->65	o->121	p->60	r->84	s->309	t->106	u->73	v->165	y->5	Ö->1	ä->37	å->24	ö->26	
ll!	H->1	J->1	
ll"	,->2	.->1	
ll,	 ->71	
ll-	 ->4	
ll.	 ->2	A->2	B->1	D->22	E->3	F->5	H->5	I->5	J->11	K->3	M->3	O->2	P->2	R->1	S->5	T->2	U->1	V->10	Ä->1	
ll:	 ->3	
ll?	.->1	D->1	H->1	J->1	K->1	
lla	 ->946	!->1	,->13	.->10	:->1	d->10	m->1	n->375	r->30	s->48	t->5	v->1	
llb	a->78	e->1	i->1	o->3	r->4	
lld	 ->5	a->23	e->66	h->23	r->1	
lle	 ->532	,->3	.->1	g->206	h->3	k->13	l->17	n->111	r->1072	s->11	t->187	u->2	
llf	i->1	o->6	r->27	u->1	ä->98	ö->20	
llg	j->1	o->1	r->2	ä->21	å->26	ö->1	
llh	a->43	e->3	ö->8	
lli	 ->1	!->1	a->7	b->1	e->1	g->88	h->1	n->2	s->5	t->29	v->1	
llk	a->1	l->2	o->75	ä->9	
llm	a->1	o->1	y->2	ä->128	ö->6	
lln	a->45	i->141	ä->6	
llo	 ->5	b->2	j->2	k->1	l->1	m->1	r->41	
llp	o->1	
llr	a->10	e->6	i->2	ä->81	
lls	 ->85	,->4	.->9	?->1	a->35	b->1	e->16	f->1	h->1	i->1	k->14	l->3	m->4	o->1	r->2	s->4	t->78	v->5	y->5	ä->5	
llt	 ->353	,->17	.->10	:->1	;->1	a->3	f->40	i->83	j->3	m->1	r->8	s->77	
llu	t->15	
llv	a->75	e->87	i->2	ä->31	
lly	 ->1	!->1	.->1	b->1	s->1	w->1	
llä	g->20	m->177	n->2	
llå	n->4	t->55	
llö	s->2	
lm 	d->1	
lm,	 ->1	
lm.	H->1	
lma	j->1	k->1	n->427	r->2	s->1	
lme	d->3	n->3	r->1	
lmo	s->1	
lms	h->1	
lmy	n->2	
lmä	n->125	r->2	s->2	t->2	
lmå	e->2	
lmö	j->2	s->1	t->3	
ln 	"->1	a->1	f->3	i->2	k->1	m->1	o->3	t->5	ä->2	
ln,	 ->2	
ln.	D->1	
lna	 ->1	,->1	d->44	
lni	n->212	s->1	
lns	 ->2	
lnä	r->6	
lo 	g->2	i->1	m->1	o->3	r->1	å->1	
lo,	 ->3	
loa	k->1	
lob	a->12	b->10	
loc	k->10	
lod	 ->2	e->2	l->1	
log	 ->31	,->2	.->7	e->10	i->45	s->4	
loj	a->7	
lok	 ->1	a->46	e->1	t->5	
lol	a->1	j->1	
lom	a->11	e->1	m->3	r->1	s->3	ä->1	
lon	a->2	i->1	m->1	
loo	i->1	
lop	p->21	
lor	 ->25	,->6	.->13	a->21	e->19	g->1	n->5	s->3	
los	 ->5	i->2	o->5	s->3	
lot	 ->1	e->1	p->2	t->12	
lov	 ->2	a->15	e->1	o->3	v->2	y->1	
loy	d->1	
lp 	a->27	d->1	f->6	n->1	o->2	p->1	s->2	t->5	v->2	ö->1	
lp,	 ->2	
lp.	D->1	H->1	I->1	J->1	V->1	
lpa	 ->37	n->3	r->8	t->1	
lpe	 ->1	n->4	r->2	s->1	
lpl	a->1	i->1	
lpo	l->45	
lpr	o->4	
lps	.->1	
lpt	 ->1	a->1	e->1	
lpu	n->2	
lpv	i->1	
lra	 ->9	n->1	p->1	
lre	 ->6	g->5	s->4	
lri	k->5	n->1	s->1	
lro	l->1	
lru	m->1	
lry	c->1	
lrä	c->75	k->2	t->11	
ls 	C->1	a->17	b->4	d->5	e->2	f->8	g->1	h->14	i->20	k->3	l->2	m->9	n->1	o->7	p->9	s->11	t->8	u->4	v->9	ä->3	å->6	ö->1	
ls,	 ->4	
ls-	 ->1	
ls.	D->4	F->1	H->1	N->1	T->1	U->1	Y->1	
ls?	V->1	
lsa	 ->15	,->3	.->1	c->3	m->32	n->4	r->1	t->4	v->1	
lsb	e->1	u->1	
lsd	o->1	r->1	
lse	 ->139	,->12	-->1	.->20	a->1	b->1	f->11	h->1	k->13	l->5	m->1	n->55	o->1	r->176	u->1	v->2	x->1	
lsf	a->2	l->2	r->2	ö->2	
lsh	a->2	i->1	
lsi	d->1	g->1	k->1	n->22	t->1	
lsk	-->1	a->31	e->1	i->1	n->1	o->4	r->8	t->3	u->1	v->1	y->5	ö->1	
lsl	a->5	i->1	o->1	u->1	ö->2	
lsm	e->1	y->9	ä->6	
lsn	i->2	y->1	
lso	-->1	c->1	e->1	m->3	n->5	r->5	s->1	v->3	
lsp	a->1	l->2	o->2	r->4	u->6	
lsr	i->2	u->3	
lss	e->2	i->1	j->1	t->5	y->1	ä->43	
lst	 ->35	,->7	.->5	a->7	e->1	h->3	i->9	o->45	r->5	u->1	v->1	ä->41	å->28	ö->2	
lsu	m->1	t->4	
lsv	a->4	i->1	ä->2	
lsy	n->3	s->6	
lsä	m->1	t->123	
lsö	k->6	
lt 	-->2	1->1	2->1	7->1	9->1	E->4	S->2	a->47	b->23	d->54	e->37	f->66	g->16	h->12	i->59	j->2	k->47	l->4	m->33	n->20	o->54	p->29	r->18	s->87	t->26	u->31	v->37	y->1	ä->14	å->4	ö->12	
lt,	 ->24	
lt.	 ->1	D->10	E->1	H->3	I->1	J->2	M->2	O->1	U->1	V->6	
lt:	 ->1	
lt;	 ->2	
lt?	J->1	
lta	 ->25	,->3	g->31	k->1	l->3	r->11	s->1	t->111	
ltb	a->1	
lte	 ->2	,->2	n->40	r->22	s->3	t->9	
ltf	l->1	ö->39	
lth	e->8	
lti	b->1	d->80	e->3	g->26	h->1	l->18	m->1	n->10	s->1	
ltj	ä->3	
ltm	e->1	
ltn	i->48	
lto	g->2	n->1	
ltr	a->3	e->1	o->1	ä->7	
lts	 ->13	.->1	:->1	a->1	e->3	i->1	å->63	
ltu	r->146	
ltä	c->4	
luc	k->5	
lud	d->2	e->4	
luf	t->2	ö->1	
lug	n->6	
luk	a->3	t->2	
lum	p->4	r->1	
lun	c->1	d->15	t->5	
lup	s->1	
lur	a->3	e->1	
lus	 ->2	i->20	s->2	t->10	
lut	 ->140	,->14	.->12	;->1	a->158	b->5	e->78	f->9	g->8	h->2	i->105	k->1	l->72	n->55	p->1	r->3	s->89	v->3	ä->5	
lux	,->1	
lv 	a->5	b->2	d->1	f->5	g->1	h->3	i->3	k->1	m->2	o->3	s->7	t->3	u->2	v->2	ä->3	å->1	
lv,	 ->5	
lv.	D->1	J->1	K->1	V->1	
lva	 ->68	,->3	.->5	l->1	n->1	r->74	
lvb	e->3	i->1	ä->1	
lve	r->126	t->1	
lvf	a->2	ö->1	
lvh	j->2	
lvi	d->1	l->1	n->1	s->40	
lvk	l->20	o->1	
lvm	i->1	
lvn	i->3	
lvo	f->1	l->1	
lvp	l->1	
lvr	a->6	
lvs	t->15	ä->1	
lvt	 ->7	i->3	
lvv	ä->2	
lvä	g->11	n->3	r->2	x->20	
lvå	r->5	
lvö	,->1	.->1	n->1	
ly 	f->1	å->1	
ly!	 ->1	
ly,	 ->2	
ly.	A->1	V->1	
lyb	e->1	
lyc	k->125	
lyd	a->3	e->5	
lyf	t->13	
lyg	,->1	a->2	b->1	e->2	k->1	n->1	p->4	s->4	t->2	
lyk	t->17	
lym	 ->2	e->2	p->2	
lyr	 ->1	
lys	 ->27	,->4	.->5	?->2	a->11	e->23	n->4	s->29	t->2	
lyt	a->12	e->1	t->17	
lyv	e->1	
lyw	o->1	
lz 	e->1	s->2	
lze	n->1	
lzm	a->2	
läc	k->8	
läd	e->22	j->15	s->6	
läg	a->1	e->50	g->293	l->1	n->8	r->11	s->12	
läk	a->5	e->1	t->5	
läm	n->86	p->228	
län	d->215	g->108	k->2	n->1	t->1	
läp	a->1	p->20	
lär	 ->1	a->9	d->8	l->1	o->2	t->3	
läs	 ->3	a->3	b->2	e->6	f->1	k->1	n->2	t->6	
lät	 ->5	t->56	
läx	a->2	o->1	
lå 	E->1	a->6	b->1	e->4	f->6	i->1	k->4	m->2	n->1	p->1	r->1	s->2	v->4	
låd	a->1	e->12	
låe	n->1	
låg	 ->7	a->5	e->1	t->2	
lån	a->1	b->1	g->121	i->1	
lår	 ->43	"->1	.->2	?->1	
lås	 ->25	.->1	e->3	s->1	t->3	
låt	 ->24	a->50	e->30	i->3	l->5	n->6	s->6	
léc	h->1	
löd	e->3	i->1	
löf	t->11	
löj	a->6	e->3	
lök	m->1	
löm	m->16	s->1	t->4	
lön	 ->1	a->2	e->3	s->5	t->4	
löp	a->8	e->10	t->7	
lör	d->1	
lös	 ->5	.->1	a->51	e->5	g->1	h->44	n->52	r->1	t->19	
löt	 ->3	s->4	
löv	s->1	
løn	,->2	
m "	E->2	K->2	n->1	o->1	v->1	ö->1	
m -	 ->19	
m 1	 ->1	5->1	6->1	9->3	
m 2	0->3	8->1	
m 3	-->2	1->1	5->3	
m 4	0->3	5->1	
m 5	0->1	b->1	
m 6	,->1	
m 8	0->1	
m A	g->1	h->1	l->2	m->3	p->1	t->1	
m B	S->1	a->1	e->6	l->1	o->1	r->2	
m C	E->1	e->1	o->2	
m D	a->4	e->2	i->1	u->1	
m E	G->3	M->1	U->20	h->1	l->1	r->1	t->1	u->73	
m F	B->1	P->1	l->1	r->2	ö->4	
m G	U->1	a->1	e->2	o->2	r->2	
m H	a->5	e->1	i->1	
m I	N->1	n->1	r->1	s->1	t->2	
m J	o->2	ö->2	
m K	a->1	o->5	
m L	a->6	i->1	l->1	
m M	a->2	c->2	
m N	e->1	
m O	f->1	
m P	P->1	a->3	o->4	r->1	
m R	a->1	i->1	o->1	
m S	E->1	c->3	e->2	j->1	k->1	p->1	y->1	
m T	a->1	h->3	i->2	o->2	u->4	
m V	ä->1	
m W	a->2	i->1	
m a	 ->1	b->2	c->1	d->2	g->4	l->59	m->2	n->67	p->1	r->22	s->5	t->398	v->80	
m b	)->1	a->7	e->138	i->12	l->11	o->15	r->13	u->4	y->2	ä->7	å->5	ö->16	
m c	)->1	a->1	e->1	h->2	o->2	
m d	a->9	e->666	i->20	j->1	o->6	r->16	u->2	y->1	ä->12	å->8	ö->4	
m e	f->13	g->6	j->1	k->5	l->10	m->18	n->205	r->16	t->126	u->10	x->15	
m f	a->32	e->2	i->44	j->1	l->12	o->23	r->65	u->6	y->2	ä->2	å->9	ö->295	
m g	a->7	e->50	i->4	j->10	l->1	o->8	r->19	ä->22	å->12	ö->37	
m h	a->205	e->57	i->14	j->6	o->14	u->34	y->1	ä->42	å->9	ö->7	
m i	 ->149	c->4	d->1	f->2	g->1	h->1	n->208	s->1	
m j	a->136	o->6	u->14	ä->3	
m k	a->68	e->1	l->2	o->200	r->27	u->9	v->2	ä->12	ö->2	
m l	a->21	e->38	i->41	j->1	o->1	y->6	ä->27	å->4	ö->5	
m m	a->108	e->84	i->33	o->16	u->1	y->17	ä->14	å->40	ö->52	
m n	a->13	e->4	i->71	o->2	u->26	y->7	ä->17	å->30	ö->2	
m o	a->1	b->2	c->92	f->7	g->1	l->6	m->61	n->1	r->17	s->4	t->1	
m p	a->25	e->7	l->4	o->8	r->23	u->4	å->66	
m r	a->57	e->98	i->15	o->1	u->3	y->2	ä->16	å->36	ö->17	
m s	.->1	a->52	c->1	e->17	i->14	j->4	k->140	l->8	m->3	n->3	o->135	p->13	t->89	u->4	v->3	y->21	ä->23	å->29	ö->3	
m t	.->3	a->22	i->126	j->3	o->10	r->30	u->1	v->6	y->11	ä->4	
m u	n->42	p->36	r->9	t->83	
m v	a->65	e->29	i->369	o->5	r->1	u->1	ä->15	å->19	
m y	r->1	t->4	
m Ö	s->4	
m ä	g->4	n->30	r->192	t->1	v->15	
m å	k->2	l->2	r->18	s->7	t->25	
m ö	a->1	k->4	m->1	n->1	p->7	r->1	s->2	v->24	
m!D	e->2	
m!M	e->1	
m!T	r->1	
m".	D->1	
m) 	o->1	
m);	 ->1	
m, 	K->1	a->9	b->4	d->13	e->10	f->7	g->2	h->6	i->7	j->3	k->4	l->1	m->12	n->5	o->23	p->5	r->1	s->17	t->2	u->9	v->13	ä->9	å->1	
m- 	o->1	
m-e	l->1	
m. 	D->3	H->2	M->1	a->2	d->1	i->1	ä->2	
m.(	A->1	
m.,	 ->1	
m..	 ->1	(->1	
m.A	l->1	t->1	v->3	
m.B	e->1	u->1	
m.D	e->38	ä->5	
m.E	G->1	K->1	n->1	u->1	x->1	
m.F	r->5	ö->3	
m.G	e->2	ö->1	
m.H	e->10	u->2	
m.I	 ->4	n->2	
m.J	a->17	
m.K	o->2	u->1	
m.L	å->1	
m.M	a->1	e->12	å->1	
m.N	a->1	e->1	i->1	u->1	ä->3	å->1	
m.O	M->1	c->4	m->2	
m.P	r->2	
m.R	e->2	å->1	
m.S	a->1	l->2	o->2	t->2	y->1	å->1	
m.T	i->1	r->1	y->1	
m.U	r->1	
m.V	a->1	e->1	i->19	
m.m	.->1	
m.Ä	n->1	r->1	
m/r	i->1	
m: 	A->1	N->1	d->3	e->1	p->1	
m; 	d->2	
m?D	e->1	
m?J	a->1	
m?M	e->1	
m?V	i->2	
mI.	 ->1	
ma 	-->2	1->1	B->1	E->1	H->2	M->1	a->25	b->13	d->25	e->12	f->30	g->4	h->12	i->47	j->5	k->18	l->7	m->31	n->9	o->17	p->24	r->17	s->111	t->15	u->15	v->14	ä->3	å->5	ö->9	
ma,	 ->10	
ma.	D->1	H->2	J->4	O->2	V->1	
ma:	 ->2	
mac	e->1	
mad	 ->1	e->10	
maf	f->1	
mag	e->2	h->1	i->1	n->2	o->4	
mai	l->1	n->7	
maj	 ->5	,->1	.->2	o->41	
mak	o->1	r->6	t->46	ä->1	
mal	 ->7	a->7	i->5	t->11	
man	 ->654	!->242	,->171	.->5	:->1	a->54	b->6	d->105	e->9	f->15	g->20	h->101	i->34	j->1	k->12	l->3	n->32	o->2	s->69	t->38	ö->1	
map	l->1	
mar	 ->45	!->1	,->14	.->4	b->88	e->84	g->6	i->3	k->232	l->1	n->26	s->11	
mas	 ->13	,->1	k->9	o->1	s->11	t->15	
mat	 ->14	.->1	c->2	e->36	f->4	i->118	n->1	p->2	s->2	t->4	u->1	
mav	t->3	
max	b->1	i->7	
mb 	h->1	
mb.	A->1	
mba	d->1	l->1	n->47	r->4	s->1	t->2	
mbe	d->1	n->4	r->47	s->2	t->10	x->1	
mbi	n->1	t->26	
mbl	e->1	i->5	
mbn	i->1	
mbo	l->9	r->1	
mbr	o->2	y->1	
mbu	d->12	l->1	r->8	s->1	
mby	g->1	
mbä	r->4	
md 	a->1	h->1	i->1	o->1	t->2	v->1	
md,	 ->2	
mda	 ->8	,->1	
mde	 ->5	.->1	f->1	n->1	s->1	
mdh	e->1	
mdi	r->1	
mdr	i->6	
mdö	m->2	
me 	e->1	f->6	k->1	o->3	s->4	å->2	
me,	 ->1	
me-	f->1	
me.	K->1	
med	 ->1525	,->14	.->6	a->25	b->184	d->59	e->217	f->22	g->22	h->1	i->15	k->5	l->354	v->61	
meg	a->1	
mek	a->11	
mel	l->291	s->146	
men	 ->531	,->26	.->17	;->2	?->1	a->33	d->45	e->5	i->55	s->415	t->862	
mer	 ->1051	!->2	,->15	.->27	a->57	f->22	g->1	i->36	n->22	p->1	s->9	v->5	
mes	,->1	g->1	t->48	
met	 ->152	)->3	,->15	.->28	:->1	?->1	a->11	e->5	o->29	r->1	s->3	
meu	r->4	
mex	i->2	
mfa	r->1	t->83	
mfi	n->1	
mfl	y->1	
mfo	r->4	
mfu	n->5	
mfä	l->1	
mfå	n->2	
mfö	r->362	
mge	r->1	
mgi	c->2	v->2	
mgr	i->4	
mgä	n->1	
mgå	 ->2	.->1	e->1	n->43	r->16	t->3	
mhe	t->100	
mhu	l->1	
mhä	l->49	r->1	v->4	
mhå	l->17	
mhö	g->14	l->2	
mi 	-->1	a->1	m->5	o->12	ä->1	
mi,	 ->3	
mi.	D->2	F->1	
mi?	 ->1	
mib	e->2	
mid	d->13	i->4	
mie	r->8	
mif	i->1	
mig	 ->210	!->1	,->15	.->5	:->1	?->1	a->1	h->2	r->11	t->1	
mii	n->1	
mik	 ->2	a->6	o->1	r->6	
mil	d->4	i->10	j->282	l->7	s->1	ä->1	ö->1	
min	 ->171	,->3	.->5	a->80	d->53	e->47	g->8	i->124	n->50	o->24	s->124	u->21	ä->3	
mip	a->1	
mir	a->1	e->5	
mis	-->2	.->1	k->223	m->5	s->1250	t->20	ä->2	
mit	 ->37	,->3	.->2	a->1	e->7	i->4	n->1	r->5	s->2	t->130	
miu	m->3	
mix	.->1	e->1	
miä	r->10	
miå	l->1	
mja	 ->36	.->1	n->17	r->6	s->1	t->1	
mju	k->3	
mka	 ->1	r->2	s->1	t->2	
mko	m->10	
mkr	i->15	
mla	 ->38	d->2	g->12	n->3	r->3	s->2	t->5	
mle	n->1	v->1	
mli	g->113	k->13	n->59	
mlo	k->2	
mlä	g->8	n->1	s->3	x->1	
mlö	s->5	
mm 	a->1	
mma	 ->406	,->7	.->5	:->2	d->5	l->4	n->320	p->1	r->96	s->7	t->6	
mme	 ->17	,->1	l->143	n->124	r->804	t->79	
mmi	g->11	p->1	s->1150	t->103	
mmo	n->1	r->10	
mmu	n->34	
mmö	b->1	
mn 	K->1	b->1	i->1	k->1	m->3	o->1	p->1	s->3	
mn,	 ->3	
mn.	D->2	M->1	V->1	
mna	 ->70	,->2	.->1	d->10	n->4	r->74	s->14	t->18	v->2	
mnb	e->1	
mnd	a->8	e->18	
mne	 ->3	.->2	:->1	n->21	r->5	t->6	
mni	n->85	
mnk	o->2	
mns	 ->8	.->1	
mnt	 ->9	,->2	.->2	s->6	
mnu	p->4	
mnv	i->1	ä->1	
mo,	 ->2	
mob	i->7	
moc	o->1	
mod	 ->7	e->58	i->7	l->12	
mof	o->1	
mog	e->4	r->3	
mok	o->5	r->137	
mol	n->1	
mom	e->5	r->3	s->1	
mon	 ->1	b->1	e->7	i->19	n->1	o->20	s->7	t->12	
mor	 ->8	,->1	.->1	a->7	d->53	g->39	s->6	u->1	
mos	 ->1	e->1	o->1	
mot	 ->325	!->7	,->17	.->4	a->1	e->26	g->1	i->22	o->9	p->4	s->73	t->17	v->6	å->3	
mou	t->1	
mp 	J->1	a->2	f->2	i->3	m->5	s->1	
mp.	D->1	
mpa	 ->69	d->2	g->1	k->1	n->10	r->13	s->45	t->16	
mpe	l->111	n->26	r->9	t->11	
mpi	c->1	s->1	
mpl	a->11	e->35	i->77	
mpn	i->85	
mpo	n->7	p->1	r->9	
mpr	o->48	ö->8	
mps	o->1	
mpt	o->1	
mpu	l->6	n->1	
mpå	l->1	
mra	 ->3	d->11	n->1	p->2	r->3	s->2	t->2	
mre	 ->6	s->1	
mri	n->1	
mru	m->2	n->1	
mrä	t->1	
mrå	d->325	
mrö	s->57	
ms 	B->1	a->2	e->2	f->1	i->1	s->1	t->1	u->1	v->1	
ms-	 ->3	,->1	
msa	 ->3	n->2	r->1	v->2	
msb	e->2	r->1	
mse	s->5	
msf	r->3	u->1	
msg	r->1	
msh	a->1	e->1	
msi	d->1	g->2	
msk	 ->1	a->7	i->1	j->1	r->1	y->4	
msl	a->12	u->3	ä->27	
msn	i->11	
mso	l->1	r->9	
msp	a->1	l->1	ä->1	
msr	e->1	ä->1	å->2	
mss	t->284	
mst	 ->46	.->1	a->14	e->79	f->1	h->1	k->1	o->86	r->15	ä->74	å->7	ö->1	
msv	e->1	ä->1	
msy	n->3	r->3	
msä	t->8	
mså	t->1	
mt 	A->1	G->1	H->1	W->1	a->22	b->7	d->3	e->11	f->14	h->4	i->5	j->1	k->5	l->3	m->6	n->1	o->15	p->4	r->7	s->13	t->10	u->9	v->4	y->1	ä->3	å->1	ö->3	
mt,	 ->6	
mt.	D->1	P->1	U->1	Å->1	
mta	 ->3	g->5	l->17	n->2	r->1	s->1	t->1	
mte	 ->14	d->2	
mti	d->174	e->1	o->4	
mtl	i->25	
mtn	i->1	
mto	n->5	
mtr	ä->2	
mts	 ->3	a->1	
mtv	i->2	
mty	c->6	
mtä	n->1	
mtå	l->1	
mug	g->1	
mul	a->8	e->26	l->1	t->9	
mum	 ->4	
mun	.->1	a->3	e->10	i->20	t->29	
mur	a->1	
mus	 ->1	-->1	i->4	s->3	
mut	f->1	o->1	s->3	
mva	n->5	
mve	r->4	t->2	
mvi	k->2	l->3	s->1	
mvä	g->2	l->4	n->5	r->1	x->1	
myc	k->452	
myg	g->1	
myl	l->1	
myn	d->162	n->2	
myt	i->1	
mán	,->1	
mäd	e->1	
mäk	t->3	
mäl	a->3	d->1	e->1	n->12	s->2	t->2	
män	 ->63	,->1	.->3	d->3	g->23	h->47	i->1	n->163	s->46	t->17	
mär	k->129	r->1	t->2	
mäs	s->31	t->2	
mät	a->4	e->1	i->1	t->3	
må 	E->1	a->1	b->2	e->1	f->4	h->2	l->2	m->4	o->33	p->1	r->1	s->5	v->1	å->1	
må,	 ->2	
må.	D->1	
måe	n->2	
måf	ö->6	
måg	a->31	r->1	
måh	ä->5	
mål	 ->99	,->16	-->1	.->17	:->1	a->1	e->43	i->5	m->1	s->21	
mån	 ->22	,->1	a->74	d->4	e->2	g->161	i->4	s->1	
mår	.->2	i->1	s->2	
mås	k->1	t->696	
måt	 ->12	,->3	.->7	g->1	t->5	
mé 	o->2	p->1	
méa	v->1	
mék	o->1	
mén	 ->1	.->1	
més	 ->1	
möb	l->2	
möd	a->3	o->1	r->1	
mög	e->1	n->1	
möj	l->307	
mön	s->2	
mör	 ->2	d->5	k->2	
mös	s->1	
möt	a->10	e->130	s->2	t->1	
möv	e->2	
n "	E->1	L->1	T->2	d->2	e->3	h->1	n->1	r->2	s->1	u->1	å->1	
n (	1->3	A->5	B->2	C->2	E->1	F->1	H->21	I->1	K->1	e->1	f->3	i->1	m->1	o->1	s->1	
n ,	 ->1	
n -	 ->72	
n 1	 ->13	,->1	0->7	1->2	2->6	3->4	4->7	5->3	6->2	7->4	8->5	9->42	
n 2	 ->2	,->1	0->17	1->2	3->1	4->1	6->3	8->1	9->1	
n 3	 ->4	,->2	0->3	1->3	4->1	8->1	9->1	
n 4	 ->3	,->2	
n 5	 ->3	0->1	2->1	7->1	
n 6	 ->1	
n 7	 ->2	9->1	
n 8	 ->2	9->1	
n 9	 ->2	0->1	5->1	
n A	B->2	D->1	c->1	f->1	l->3	m->6	n->1	r->1	t->2	u->1	
n B	S->1	a->3	e->4	o->2	r->5	
n C	E->4	a->2	e->1	h->1	r->2	
n D	a->4	e->6	u->1	
n E	G->3	K->1	M->1	U->6	i->1	n->3	r->6	u->50	
n F	E->1	M->1	N->1	l->4	o->2	r->2	ö->2	
n G	U->1	a->3	o->2	r->3	ö->1	
n H	a->4	e->2	u->23	
n I	 ->2	M->1	R->1	X->1	m->2	n->3	s->14	
n J	a->3	o->1	u->2	
n K	a->5	i->4	o->7	y->2	ö->2	
n L	a->3	e->1	i->1	o->2	
n M	a->1	i->1	
n N	a->5	i->1	o->1	
n O	S->1	
n P	P->2	R->1	S->1	a->3	l->1	o->5	r->7	
n R	a->2	e->2	o->3	
n S	P->1	S->1	a->3	c->2	e->1	h->2	o->1	y->5	ã->1	
n T	a->4	e->1	h->1	o->1	y->4	
n U	N->1	S->1	n->2	
n V	I->2	a->3	e->2	i->1	
n W	a->1	i->4	o->18	u->1	
n X	X->1	
n a	 ->1	b->4	c->15	d->8	g->4	k->12	l->71	m->5	n->249	p->2	r->30	s->8	t->429	u->3	v->558	x->1	
n b	a->40	e->223	i->42	l->39	o->30	r->45	u->13	y->11	ä->28	å->3	ö->56	
n c	e->11	h->9	o->6	
n d	a->30	e->557	i->36	j->8	o->15	r->18	u->3	y->2	ä->57	å->18	ö->12	
n e	f->55	g->26	j->2	k->55	l->41	m->7	n->238	p->1	r->23	t->55	u->145	v->4	x->28	
n f	a->43	e->12	i->43	j->7	l->14	o->40	r->239	u->26	y->6	ä->6	å->48	ö->798	
n g	a->36	e->179	i->9	j->14	l->14	n->2	o->35	r->82	u->1	y->1	ä->27	å->75	ö->51	
n h	a->395	e->51	i->13	j->10	o->28	u->17	y->2	ä->111	å->21	ö->35	
n i	 ->592	,->1	b->1	c->4	d->10	f->3	g->1	h->2	l->3	m->1	n->503	r->3	s->12	t->5	
n j	a->133	u->30	ä->8	
n k	a->177	e->2	i->1	l->32	n->3	o->398	r->44	u->30	v->14	y->1	ä->21	ö->4	
n l	a->25	e->24	i->45	o->13	u->1	y->13	ä->50	å->26	ö->24	
n m	.->1	a->86	e->319	i->75	o->67	u->4	y->81	ä->20	å->159	ö->27	
n n	a->36	e->13	i->17	o->14	u->46	y->85	ä->59	å->41	ö->17	
n o	a->6	b->27	c->682	e->4	f->34	h->1	k->5	l->17	m->435	n->4	p->6	r->59	s->6	t->4	u->3	v->5	ä->1	ö->3	
n p	.->1	a->40	e->34	l->26	o->82	r->58	u->29	y->1	å->270	
n r	a->42	e->187	i->41	o->12	u->3	y->1	ä->61	å->27	é->1	ö->24	
n s	a->108	c->2	e->61	i->67	j->34	k->309	l->28	m->5	n->23	o->407	p->30	r->1	t->266	u->9	v->11	y->25	ä->58	å->102	ö->3	
n t	.->1	a->80	e->18	i->371	j->8	o->22	r->60	u->15	v->53	y->47	ä->10	
n u	n->95	p->106	r->13	t->160	
n v	a->120	e->69	i->371	o->4	r->1	u->1	ä->64	å->18	
n w	a->1	e->1	
n y	t->8	
n z	i->2	
n Ö	s->3	
n ä	g->9	l->1	n->53	r->313	v->32	
n å	 ->8	b->1	k->8	l->4	r->10	s->28	t->50	
n ö	d->1	k->32	m->1	n->9	p->8	r->1	s->18	v->80	
n! 	A->5	B->2	D->33	E->6	F->12	G->2	H->1	I->10	J->75	K->5	L->6	M->6	N->6	O->2	P->4	R->4	S->9	T->8	U->4	V->17	Ä->7	Å->3	Ö->1	
n!A	m->1	
n!D	e->3	
n!E	f->1	n->1	
n!H	e->1	
n!J	a->6	
n!M	i->1	
n!N	ä->2	
n!R	ö->1	
n!S	a->1	
n!T	a->1	i->1	
n!U	n->1	
n!V	i->2	
n" 	a->2	e->1	g->1	i->1	o->1	p->1	s->1	
n",	 ->5	
n".	D->3	O->1	R->1	
n) 	(->3	f->1	h->1	z->1	
n)(	P->2	
n),	 ->1	
n).	D->2	H->1	
n)J	a->1	
n)N	ä->1	
n, 	"->1	1->4	5->1	8->1	A->2	B->5	C->1	D->1	E->2	I->2	J->1	K->4	L->2	N->1	O->1	P->4	R->2	S->3	T->2	U->1	V->2	W->1	a->35	b->22	d->69	e->53	f->100	g->9	h->74	i->51	j->12	k->56	l->8	m->85	n->30	o->135	p->18	r->6	s->141	t->32	u->35	v->59	y->1	Î->1	ä->44	å->1	ö->1	
n- 	o->4	
n-C	l->1	
n-H	a->1	
n-K	e->1	
n-S	S->1	
n-g	r->1	
n-r	å->3	
n. 	D->8	F->1	H->2	I->2	J->3	L->1	M->3	N->1	O->3	R->1	V->2	
n."	 ->1	
n.(	E->1	I->1	L->1	P->2	
n.)	 ->2	.->1	A->1	B->4	F->3	G->1	H->1	
n..	 ->10	(->3	H->1	
n.1	4->1	5->1	
n.A	l->11	n->2	r->2	t->4	v->8	
n.B	e->3	i->1	r->2	
n.C	e->1	u->1	
n.D	E->1	e->255	ä->28	å->3	
n.E	U->2	f->4	m->1	n->17	r->2	t->10	u->5	v->1	
n.F	E->1	a->2	i->1	l->1	o->1	r->9	y->1	ö->45	
n.G	e->1	o->1	ä->1	å->1	
n.H	a->8	e->57	i->2	o->2	u->5	ä->7	
n.I	 ->37	l->1	n->7	
n.J	a->135	o->1	u->2	
n.K	a->5	o->25	r->1	u->1	v->1	
n.L	e->1	i->2	å->11	
n.M	a->8	e->40	i->7	o->4	y->1	ä->2	å->1	ö->1	
n.N	a->2	i->9	u->4	y->1	ä->9	
n.O	c->11	m->18	r->5	z->1	
n.P	a->4	e->1	l->1	r->3	å->9	
n.R	e->2	i->1	o->1	ä->1	å->4	
n.S	a->7	c->1	e->4	i->3	k->2	l->11	n->1	o->11	t->4	u->1	y->2	ä->3	å->8	
n.T	a->5	h->2	i->6	o->2	r->3	v->1	y->5	
n.U	n->10	p->1	t->4	
n.V	a->17	e->1	i->98	å->5	
n.W	o->1	
n.Ä	n->3	r->2	v->4	
n.Å	 ->3	
n.Ö	g->2	v->1	
n/N	o->2	
n/å	r->2	
n: 	"->1	A->1	D->2	E->1	H->1	J->2	K->3	R->1	T->1	V->2	a->1	d->3	e->1	f->3	i->2	j->1	m->2	n->2	v->5	
n:F	ö->1	
n; 	J->1	a->1	d->10	e->1	f->2	i->1	m->1	o->1	p->1	s->2	v->1	ä->1	
n? 	2->1	D->1	I->1	
n?.	 ->1	
n?A	n->1	
n?D	e->8	
n?E	f->1	
n?F	o->1	r->2	ö->2	
n?H	e->3	u->1	
n?I	 ->1	
n?J	a->4	
n?K	a->3	o->2	
n?N	ä->1	
n?O	m->1	
n?P	a->1	
n?S	e->1	
n?V	a->1	e->2	i->8	
n?Ä	r->4	v->1	
nFr	å->3	
nHe	r->2	
nI 	d->1	
nJa	g->2	
nNä	s->7	
na 	(->1	-->23	1->5	3->1	6->1	8->8	A->2	B->1	E->2	I->1	L->1	M->1	P->1	T->4	a->172	b->98	c->3	d->154	e->93	f->380	g->102	h->99	i->280	j->5	k->155	l->44	m->149	n->32	o->278	p->113	r->119	s->309	t->128	u->96	v->100	y->4	ä->71	å->28	ö->22	
na!	D->1	H->1	O->1	
na"	.->2	i->1	
na,	 ->258	
na-	I->1	
na.	 ->10	(->1	)->1	-->2	.->1	A->9	B->2	D->68	E->13	F->16	G->2	H->11	I->16	J->31	K->10	L->4	M->19	N->7	O->7	P->5	R->1	S->12	T->5	U->8	V->40	Ä->5	Å->1	
na/	E->1	s->1	
na:	 ->3	
na;	 ->5	
na?	E->1	H->2	I->1	J->2	M->1	P->1	S->1	V->4	Ä->1	
naH	e->1	
nab	b->72	i->1	
nac	k->10	
nad	 ->60	,->11	.->8	:->1	;->1	?->2	a->2	e->406	s->61	
naf	l->1	r->1	
nag	a->3	e->4	i->3	
nai	v->2	
nak	i->2	n->1	r->1	
nal	 ->26	,->3	-->2	.->6	a->47	e->17	f->4	i->38	l->1	p->42	r->4	s->7	t->1	u->1	v->1	y->58	
nam	b->1	i->5	m->4	n->17	
nan	 ->82	,->4	.->1	d->67	e->1	s->89	t->1	
nap	p->18	r->2	
nar	 ->241	,->7	.->13	:->1	a->37	b->1	d->1	e->52	i->6	k->7	l->1	n->17	s->23	t->27	å->1	
nas	 ->336	!->1	,->10	.->10	t->79	
nat	 ->157	,->4	.->6	e->1	i->283	s->15	t->3	u->121	
nau	e->1	
nav	g->2	i->1	t->3	
naz	i->16	
nba	n->1	r->68	
nbe	g->12	h->1	r->5	s->1	t->5	
nbi	l->8	n->1	
nbj	u->6	ö->1	
nbl	a->16	i->16	
nbo	e->1	k->2	
nbr	o->1	y->1	
nbu	d->4	l->1	n->1	r->3	
nby	g->1	
nc 	d->1	
nc,	 ->1	
nca	,->1	s->1	
nce	,->1	.->1	n->31	p->7	r->6	
nch	e->2	t->1	
nci	d->1	l->1	p->195	s->3	t->8	
nck	h->14	
nd 	(->3	-->4	8->1	E->1	L->4	S->1	T->1	a->118	b->10	c->1	d->22	e->15	f->35	g->5	h->13	i->26	j->1	k->9	l->3	m->62	n->7	o->47	p->6	r->2	s->50	t->14	u->8	v->12	ä->18	å->1	ö->1	
nd!	 ->2	
nd)	,->1	
nd,	 ->49	
nd-	 ->1	
nd.	 ->1	A->2	D->10	E->1	F->1	G->1	H->1	I->6	J->7	K->2	L->1	M->2	N->3	O->2	P->1	S->1	U->1	V->3	Å->1	
nd?	 ->1	.->1	F->1	J->1	
nda	 ->194	,->7	.->15	?->1	b->2	d->17	g->5	h->43	i->1	l->9	m->15	n->86	r->48	s->109	t->63	
ndb	a->9	e->1	u->1	
nde	 ->1738	!->9	"->1	(->1	,->117	.->141	:->37	;->4	?->4	b->11	f->13	h->1	k->10	l->92	m->6	n->385	r->942	s->129	t->458	v->8	
ndf	u->1	ä->4	ö->4	
ndg	ä->2	å->3	
ndi	 ->2	:->1	c->1	d->14	e->7	g->399	k->10	n->1	r->7	s->2	t->4	v->14	
ndk	u->1	
ndl	a->172	i->208	ä->75	ö->1	
ndm	e->3	ä->1	
ndn	a->4	i->74	
ndo	.->1	m->19	n->4	r->1	
ndp	e->1	r->1	u->103	
ndr	a->507	e->59	i->314	o->1	ä->2	
nds	 ->34	,->1	a->9	b->44	d->12	j->1	k->42	l->2	m->9	p->8	r->6	s->1	t->3	v->1	ä->1	
ndt	 ->6	,->1	e->1	
ndu	p->3	s->114	t->1	
ndv	a->26	i->41	
ndz	i->4	
ndä	r->1	
ndå	 ->56	,->1	.->1	
ndé	e->1	
ndö	v->1	
ne 	F->1	a->6	b->1	d->2	e->1	f->8	g->1	h->7	i->7	j->2	k->2	l->1	n->6	o->8	p->2	q->2	r->1	s->6	t->3	v->2	ä->2	å->1	
ne!	 ->1	
ne,	 ->9	
ne-	 ->1	A->2	M->1	s->1	
ne.	D->3	J->1	
ne:	 ->1	
nea	r->2	
neb	a->1	o->1	ä->108	ö->7	
ned	 ->21	.->2	e->9	g->2	l->5	m->3	o->1	r->3	s->7	v->13	
nee	x->1	
nef	a->6	f->3	i->5	
neg	a->26	
neh	a->3	å->78	ö->4	
nej	 ->2	,->2	.->1	
nek	a->13	
nel	a->1	e->1	i->2	l->281	n->2	s->1	t->1	u->1	
nem	a->4	
nen	 ->969	!->1	"->1	)->1	,->113	.->158	:->1	;->3	?->4	J->2	a->2	e->8	s->390	t->18	
neo	n->2	
nep	o->5	
ner	 ->480	"->1	,->52	-->10	.->58	;->1	?->5	N->2	a->99	e->22	g->111	h->46	i->64	l->14	n->208	s->32	ö->4	
nes	 ->27	,->1	e->2	i->8	m->2	r->1	s->1	t->1	
net	 ->18	,->6	.->12	a->1	e->6	i->1	t->3	ä->6	
neu	t->2	
nev	å->2	
nez	 ->1	u->1	
nfa	l->2	t->12	
nfe	d->1	k->2	r->170	s->1	
nfi	d->2	l->1	n->2	s->2	
nfl	i->16	y->13	
nfo	r->92	
nfr	a->15	e->1	i->1	o->1	å->4	
nfä	r->1	
nfö	r->226	
ng 	(->6	-->12	1->2	2->2	3->1	6->2	8->2	D->1	E->2	F->1	I->2	T->1	V->1	a->370	b->21	d->18	e->29	f->127	g->13	h->31	i->124	j->1	k->30	l->9	m->75	n->12	o->187	p->61	r->10	s->160	t->86	u->20	v->31	ä->48	å->5	ö->3	
ng!	J->1	
ng"	 ->2	,->2	.->2	
ng)	 ->4	.->1	N->1	
ng,	 ->215	
ng-	P->1	
ng.	 ->5	(->1	.->3	A->8	D->75	E->8	F->16	G->2	H->16	I->15	J->32	K->9	L->3	M->13	N->9	O->17	P->5	R->1	S->7	T->4	V->19	Ä->3	
ng:	 ->3	D->1	
ng;	 ->4	
ng?	D->2	H->1	J->1	O->1	T->1	Ä->1	
nga	 ->219	,->5	.->3	d->6	g->18	l->3	n->13	r->664	s->16	t->4	v->1	
ngb	r->1	
ngd	 ->19	a->1	e->12	o->15	p->4	r->1	y->1	
nge	 ->50	,->1	f->10	l->38	m->4	n->993	r->111	s->10	t->52	
ngf	a->15	l->1	o->21	r->2	u->1	ä->2	
ngg	å->2	
ngi	g->2	l->1	v->13	
ngk	ö->1	
ngl	e->2	i->37	
ngm	e->6	å->1	
ngn	a->8	i->44	
ngo	m->4	
ngp	o->2	
ngr	a->4	e->79	i->17	o->1	ä->1	
ngs	 ->10	-->12	a->30	b->27	c->13	d->4	e->3	f->321	g->6	h->2	i->21	k->190	l->73	m->27	n->7	o->12	p->109	r->37	s->81	t->25	u->7	v->45	y->2	ä->2	å->6	ö->1	
ngt	 ->41	,->1	.->3	a->1	e->8	g->11	i->4	o->5	v->4	
ngu	e->2	
ngv	a->6	
ngä	l->1	
ngå	 ->8	.->1	e->53	n->1	r->16	t->6	
ngö	r->3	
nha	m->1	n->48	s->1	
nhe	d->2	m->2	t->242	
nhi	l->1	
nho	 ->4	.->1	s->1	
nhu	n->1	
nhä	l->32	m->6	n->5	
nhå	l->55	r->1	
nhö	j->4	
ni 	1->6	2->2	a->25	b->10	d->7	e->4	f->15	g->5	h->24	i->15	j->3	k->17	l->3	m->3	n->8	o->8	p->3	r->5	s->33	t->7	u->5	v->24	ä->7	ö->1	
ni,	 ->16	
ni.	(->1	A->1	D->1	
nia	l->1	
nic	e->2	
nie	d->2	f->1	n->24	r->38	s->2	t->3	
nif	e->1	r->2	
nig	 ->3	a->5	h->12	t->1	
nik	 ->7	-->1	a->17	e->7	t->1	
nil	a->2	
nim	a->1	b->1	e->1	i->19	o->1	u->5	
nin	d->2	e->1	g->2448	s->1	v->1	
nio	 ->14	;->1	n->450	
nip	a->1	e->1	p->3	
nir	e->1	
nis	a->43	c->1	e->57	k->162	m->16	t->106	
nit	 ->6	,->1	.->1	e->14	i->106	o->1	s->8	t->15	u->2	z->1	ä->1	
niu	m->5	
niv	e->4	å->110	
nié	 ->1	
nj 	f->2	m->1	
nj.	D->1	
nje	 ->11	.->2	n->4	r->78	
njo	r->1	
nju	n->1	t->2	v->1	
njä	m->1	r->1	
njö	r->2	
nk 	b->1	e->1	h->1	p->1	r->1	t->1	u->1	v->1	
nk"	 ->1	
nk-	 ->1	
nk.	D->1	
nka	 ->42	,->1	.->2	l->9	n->288	r->18	s->3	t->1	
nkb	a->4	
nke	 ->48	,->2	b->1	f->1	g->1	l->48	n->25	p->1	r->52	s->1	
nkf	a->7	o->1	ö->1	
nki	r->1	t->2	
nkl	a->24	i->6	u->21	
nkn	a->4	i->15	y->1	
nko	.->1	l->1	m->19	n->6	p->1	
nkr	a->31	e->60	i->40	ä->1	
nks	 ->3	a->2	c->1	e->1	
nkt	 ->139	,->14	.->20	:->2	?->1	a->8	e->177	i->42	s->5	u->1	
nku	r->285	
nkä	n->1	
nkö	p->2	r->1	
nla	g->1	m->1	n->7	r->2	
nle	d->111	t->13	
nli	g->246	t->1	
nly	s->1	
nlä	g->32	m->5	n->8	
nlå	s->1	t->1	
nlö	p->5	s->1	
nma	n->1	r->26	
nmä	l->20	r->12	s->2	
nmö	t->2	
nn 	d->1	e->1	o->1	t->1	ä->1	
nn,	 ->2	
nn-	g->1	
nna	 ->926	,->4	.->12	?->1	b->1	d->6	g->9	k->2	l->1	m->1	n->111	r->31	s->58	t->116	
nnd	r->1	
nne	 ->22	!->1	,->5	.->2	b->117	d->1	f->6	h->85	l->5	n->58	r->199	s->28	t->9	v->2	
nnh	e->1	
nni	e->25	g->7	n->79	s->98	t->16	u->3	v->1	
nnl	a->3	i->2	y->1	ä->1	
nno	c->24	l->9	p->2	r->64	v->6	
nns	 ->338	,->3	.->7	a->4	k->1	
nnu	 ->75	.->4	;->1	
nny	t->2	
nnä	e->1	m->2	
no 	L->1	P->2	i->1	k->1	o->2	u->1	
no,	 ->2	
no.	J->1	O->1	
noc	k->24	
nod	l->3	
nog	 ->14	,->1	.->2	a->12	g->12	r->2	
noi	s->1	
nok	u->3	
nol	i->9	l->3	o->3	
nom	 ->545	,->3	.->6	a->2	b->7	d->6	e->8	f->161	g->16	i->286	l->2	r->1	s->18	t->1	
non	 ->4	,->1	.->1	?->1	e->1	y->5	
nop	o->17	r->2	
nor	 ->37	,->3	.->8	?->1	d->24	e->4	i->22	l->2	m->77	n->6	r->5	s->12	
nos	 ->4	!->1	,->2	
not	a->1	e->28	i->1	t->1	
nov	a->6	e->14	
now	-->1	
npa	s->14	
npo	r->2	
npr	i->2	o->1	ä->1	
npu	n->31	
npå	 ->1	
nr 	1->5	2->2	3->10	4->7	5->1	6->1	7->1	8->1	9->1	
nra	 ->11	d->1	r->1	s->1	
nre	 ->83	g->1	n->1	s->6	
nri	k->57	
nry	 ->1	m->1	
nrä	t->56	
nrå	d->1	
nrö	j->6	t->1	
ns 	-->1	2->2	B->3	E->3	G->1	H->1	I->1	S->1	V->1	X->1	a->84	b->66	c->2	d->97	e->94	f->135	g->30	h->26	i->103	j->7	k->50	l->33	m->111	n->38	o->97	p->51	r->94	s->146	t->49	u->60	v->52	y->9	ä->16	å->13	ö->15	
ns!	V->1	
ns,	 ->43	
ns-	 ->6	
ns.	D->12	E->2	F->1	I->1	J->3	L->1	M->3	O->1	S->1	V->1	
ns/	d->1	
ns:	 ->1	
ns;	 ->1	
ns?	.->1	E->1	J->1	
nsa	 ->14	,->1	d->27	f->2	k->1	m->223	n->4	r->14	s->5	t->66	v->2	
nsb	e->12	o->1	r->1	u->1	
nsc	h->9	
nsd	a->5	e->3	i->1	o->2	u->2	ö->1	
nse	 ->20	,->1	.->1	;->1	e->11	k->61	m->3	n->197	r->341	s->5	t->2	u->1	
nsf	o->1	r->9	u->1	ö->22	
nsg	r->1	
nsh	a->1	i->10	ä->2	
nsi	b->1	d->4	e->78	f->3	k->5	n->18	o->27	s->8	t->8	v->12	ä->1	
nsj	o->17	
nsk	 ->11	a->588	e->70	i->28	l->43	n->41	o->39	r->53	t->8	u->12	v->10	
nsl	a->45	e->19	i->22	o->8	u->29	ä->1	å->5	
nsm	e->5	i->2	o->1	y->8	ä->7	å->1	ö->1	
nsn	a->2	i->21	
nso	l->3	m->3	r->2	
nsp	a->2	e->13	i->3	l->2	o->187	r->19	
nsr	a->2	e->13	o->1	ä->43	
nss	a->7	c->1	e->1	i->1	k->4	t->23	v->1	y->6	
nst	 ->35	,->3	.->2	a->98	e->138	f->1	g->3	i->167	j->1	m->1	o->29	r->154	s->1	ä->86	å->1	
nsu	l->5	m->63	n->3	p->1	t->5	
nsv	a->311	e->1	i->10	ä->13	
nsy	n->85	
nsä	g->1	k->3	m->1	r->2	t->9	
nså	g->12	t->2	
nsö	k->10	v->13	
nt 	(->1	-->7	1->2	A->1	C->1	E->2	a->81	b->10	c->1	d->7	e->11	f->57	g->8	h->14	i->33	k->18	l->4	m->16	n->5	o->38	p->11	r->2	s->77	t->22	u->14	v->5	ä->7	å->1	ö->4	
nt!	"->1	
nt,	 ->41	
nt-	E->1	
nt.	 ->1	D->13	E->2	F->4	H->3	I->4	J->6	L->1	M->3	N->1	O->1	P->1	S->4	V->3	
nt:	 ->2	
nta	 ->122	,->1	.->2	b->4	d->1	g->79	i->1	k->17	l->77	m->2	n->28	r->109	s->27	t->28	v->1	
nte	 ->1584	!->2	,->15	.->14	:->1	?->2	g->42	k->3	l->14	m->27	n->62	r->358	s->1	t->480	x->1	
ntf	r->6	
nti	 ->19	!->3	,->3	-->3	.->3	a->3	b->1	d->1	e->29	f->21	k->4	l->3	m->3	n->83	o->41	q->1	s->12	t->13	
ntk	a->1	u->1	
ntl	i->249	
ntn	i->8	
nto	g->26	l->4	m->1	n->1	r->10	
ntp	o->2	r->1	
ntr	a->128	e->144	o->190	u->9	y->15	ä->63	å->1	
nts	 ->21	,->2	.->2	a->1	b->1	f->1	i->1	k->7	l->28	u->2	
ntt	i->1	
ntu	e->21	n->1	r->1	s->3	
ntv	a->1	e->2	ä->1	
nty	d->6	g->4	r->9	
ntä	k->5	r->2	
ntó	n->1	
ntö	r->3	
nu 	-->1	3->1	E->1	a->8	b->8	d->7	e->23	f->21	g->14	h->21	i->42	k->11	l->5	m->18	n->10	o->7	p->7	r->4	s->30	t->11	u->4	v->9	ä->17	å->1	
nu,	 ->6	
nu.	.->1	D->1	J->1	K->2	L->1	V->2	
nu:	 ->1	
nu;	 ->1	
nu?	J->1	
nua	r->16	
nuc	 ->1	
nue	r->2	
nuf	t->14	
nul	l->1	ä->1	
num	 ->4	.->1	e->5	m->2	
nun	n->1	
nup	p->4	
nus	 ->3	d->1	g->2	s->1	
nut	 ->3	.->3	e->14	n->2	p->1	s->1	t->2	v->1	
nuv	a->45	
nva	l->1	n->18	p->12	r->8	
nve	c->2	n->25	r->13	s->15	t->1	
nvi	k->5	n->12	s->41	t->1	
nvo	l->9	
nvä	g->23	n->199	r->1	
nvå	n->9	
ny 	b->1	e->1	f->4	g->1	h->1	i->2	k->8	l->3	m->1	o->2	p->2	r->2	s->6	t->1	u->1	v->3	
nya	 ->164	,->1	;->1	n->4	r->1	s->2	
nyb	a->39	i->2	
nyc	k->8	
nyd	a->1	
nye	 ->1	l->6	t->1	
nyf	a->1	ö->1	
nyh	e->13	
nyk	t->3	
nyl	i->30	
nym	 ->2	.->1	a->1	i->1	
nyn	a->6	
nyo	 ->1	n->3	
nyp	l->1	
nys	k->1	s->13	
nyt	a->5	e->2	n->1	s->1	t->122	
nyv	a->1	
nyå	r->1	
nz 	F->5	b->1	e->1	f->2	o->7	t->1	
nz)	(->1	.->1	
nz,	 ->3	
nzF	r->1	
nzb	e->1	
nze	s->1	
nzá	l->1	
nÄr	a->1	
näc	k->2	
näe	r->1	
näg	n->1	
näl	l->2	
näm	l->43	n->93	t->1	
när	 ->415	!->32	,->75	.->11	a->28	e->66	f->1	h->5	i->12	m->42	p->1	s->2	v->46	
näs	d->1	t->47	
nät	 ->5	.->1	e->4	s->1	t->1	v->11	
näv	a->1	
nå 	a->1	d->13	e->28	f->6	g->1	h->1	m->3	n->1	p->2	r->1	s->1	v->5	y->1	ä->1	å->1	ö->1	
nå,	 ->1	
nå.	 ->1	F->1	J->1	S->1	
nåb	a->2	
nåd	 ->1	a->1	d->6	
någ	o->358	r->147	
nål	a->5	
når	 ->15	i->2	
nås	 ->5	.->2	
nåt	t->20	
nço	i->1	
nèv	e->3	
nöd	b->1	e->1	i->13	s->1	v->124	
nöj	a->10	d->11	e->7	t->1	
nör	 ->1	,->1	s->2	
nös	t->19	
nöt	.->1	k->3	s->1	t->1	
növ	a->1	i->1	r->1	
o (	K->2	
o -	 ->3	
o 1	9->1	
o C	a->5	
o E	u->1	
o L	e->1	
o P	r->2	
o R	o->1	
o S	á->1	
o T	o->2	r->1	
o V	a->3	i->1	
o a	c->1	n->1	t->8	
o b	e->3	l->1	ä->1	
o d	e->1	i->1	å->1	
o e	t->1	
o f	a->2	r->2	u->1	ö->19	
o g	o->1	r->2	å->3	
o h	a->4	å->1	
o i	 ->11	n->1	
o k	a->2	o->1	v->1	ä->1	
o l	e->1	ä->1	
o m	e->2	i->7	å->4	
o n	ä->2	å->3	
o o	c->18	m->3	
o p	e->2	u->1	å->5	
o r	e->1	
o s	a->2	i->1	k->2	o->15	å->2	
o t	i->6	r->1	
o u	n->2	t->2	
o v	a->2	i->2	ä->1	
o ä	n->1	r->7	v->2	
o å	r->8	t->1	
o ö	p->1	v->1	
o!A	l->1	
o, 	A->1	H->1	T->1	W->1	a->2	d->5	e->3	f->2	h->2	i->2	k->1	m->3	o->6	s->10	t->2	v->2	ä->1	
o- 	o->1	
o-P	l->4	
o-a	f->1	n->1	
o-p	r->1	
o-r	å->1	
o. 	D->1	
o.-	 ->1	
o.A	t->1	v->1	
o.B	e->1	
o.D	e->5	ä->1	
o.E	u->1	
o.F	l->1	ö->3	
o.H	e->2	u->1	
o.J	a->5	
o.K	n->1	o->1	
o.L	å->1	
o.M	e->1	
o.N	ä->2	
o.O	c->1	m->2	r->1	
o.S	e->1	
o.T	r->1	y->1	
o.V	i->5	
o.m	.->7	
o/O	i->1	
o: 	v->1	
o; 	d->1	
o? 	D->1	
o?H	u->1	
oNä	s->1	
oU,	 ->1	
oU-	r->1	
oa 	f->1	o->1	s->1	
oac	c->31	
oad	 ->3	e->2	
oak	l->1	t->14	
oal	i->14	
oan	a->1	d->9	s->6	v->1	
oar	 ->5	d->1	e->1	
oat	e->1	
oav	b->2	s->10	
ob 	S->2	
oba	k->2	l->18	s->1	
obb	 ->2	,->2	y->12	
obe	b->1	f->1	g->5	h->2	r->60	s->5	t->1	
obi	l->7	n->1	
obj	e->1	
obl	e->184	i->14	
obo	d->3	
obs	e->2	
oc-	d->1	t->1	
oca	 ->1	
oce	d->1	n->94	s->109	
och	 ->4556	)->1	,->14	.->1	/->1	I->2	i->1	s->1	
oci	a->206	e->2	l->1	o->3	
ock	 ->75	"->1	,->8	.->3	a->9	b->1	e->5	h->3	s->589	u->5	
oco	,->1	
od 	a->9	b->2	d->4	e->3	f->19	h->1	i->9	j->2	k->2	l->1	m->5	n->1	o->2	p->4	r->2	s->9	t->8	u->1	v->2	ä->4	å->1	
od,	 ->5	
od.	D->1	F->1	V->1	
od?	-->1	
oda	 ->38	.->1	c->5	f->1	s->5	
odd	a->1	e->8	s->1	
ode	l->13	n->49	r->69	t->6	
odf	i->1	
odi	 ->17	,->1	.->2	;->1	f->5	g->4	n->1	s->22	
odj	u->2	
odk	ä->89	
odl	a->3	i->14	
odo	.->3	n->1	s->1	
ods	 ->30	,->1	.->4	;->1	N->1	e->2	
odt	a->38	o->2	y->6	
odu	c->31	g->1	k->53	
odw	i->1	
oeb	b->1	
oed	t->14	
oef	f->3	t->1	
oeg	e->5	
oek	 ->1	o->9	
oel	i->1	v->1	
oen	d->130	i->4	s->4	
oer	h->12	s->1	
oet	 ->1	i->1	t->6	
of 	-->1	a->1	e->2	f->5	h->2	i->3	k->1	l->1	o->2	s->4	t->1	u->1	ä->1	
of,	 ->4	
of.	D->2	E->1	J->1	
ofa	l->1	n->2	
ofd	r->1	
ofe	d->1	l->1	m->2	n->20	r->32	s->7	
off	e->93	i->5	r->16	
ofh	j->1	
ofi	 ->2	,->1	l->4	n->4	s->1	
ofo	b->1	
ofr	e->1	å->3	
ofs	i->1	t->3	
oft	 ->1	a->54	
ofu	l->2	
ofö	r->25	
og 	1->1	a->6	b->4	d->5	e->8	f->5	h->4	i->9	k->4	l->5	m->12	n->2	o->4	p->2	r->4	s->7	t->3	u->9	v->1	ä->1	å->1	ö->1	
og,	 ->3	
og.	D->2	F->2	H->1	J->2	M->2	N->1	S->1	
oga	 ->15	,->1	.->2	d->3	m->2	n->13	r->17	t->4	u->18	
ogb	e->1	
oge	 ->1	,->1	n->48	r->2	t->2	
ogg	r->12	
ogi	 ->4	.->2	k->8	n->1	s->34	
ogj	o->1	
ogk	u->1	
ogm	 ->1	a->1	
ogr	a->252	e->1	i->1	u->3	
ogs	 ->26	,->2	a->2	b->6	e->1	f->1	k->1	o->1	p->1	s->4	u->1	v->1	ä->2	
ogu	e->1	
ogy	n->1	
ogå	r->1	
ogö	r->9	
oha	n->3	
ohe	r->1	
ohj	a->1	ä->1	
oho	l->1	
ohä	m->1	
ohö	v->1	
oig	e->1	
oij	-->1	
oin	s->2	t->4	
oir	e->3	m->1	
ois	 ->1	e->1	k->1	s->1	t->2	
oja	l->7	
oje	k->64	
ojk	a->1	o->1	
ojo	s->1	
oju	s->6	
ojä	m->7	
ok 	a->1	d->1	f->2	g->1	h->1	i->1	m->1	o->9	s->4	t->1	ä->2	
ok,	 ->5	
ok.	D->1	H->1	J->1	T->1	V->1	
oka	 ->2	l->44	s->1	t->5	
oke	n->38	r->1	
oki	g->2	
okl	a->16	
oko	 ->5	l->26	n->3	r->1	
okr	a->138	e->2	i->2	ä->1	
oks	l->1	t->1	
okt	 ->5	o->8	
oku	l->3	m->46	n->3	s->5	
okä	n->2	
ol 	a->2	b->1	d->1	f->2	i->3	m->2	o->9	s->4	t->1	v->1	
ol,	 ->7	
ol-	 ->1	f->1	
ol.	D->1	E->2	H->1	K->1	M->1	
ol;	 ->1	
ola	 ->6	,->1	d->1	g->16	n->17	r->25	v->1	
olb	e->2	
old	a->2	i->5	
ole	 ->1	m->1	n->48	r->25	u->1	
olf	 ->2	e->4	r->1	s->3	ö->2	
oli	b->1	c->4	d->33	g->18	k->133	n->1	s->25	t->534	v->3	
olj	a->10	e->32	
olk	 ->14	,->1	.->8	a->17	e->21	f->1	g->2	h->9	l->1	n->57	o->7	p->10	r->5	s->6	v->2	
oll	 ->93	!->1	,->20	-->1	.->28	:->1	a->10	e->309	f->1	i->3	m->5	n->2	o->2	r->1	s->4	u->15	v->1	y->1	
olm	 ->1	,->1	.->1	
oln	 ->1	
olo	g->31	n->1	r->3	s->1	
olp	e->1	
ols	 ->3	a->1	b->1	f->2	i->1	k->5	p->1	s->1	t->1	u->1	v->1	
olt	 ->6	a->3	h->2	
olu	n->4	t->141	
olv	 ->1	e->10	
oly	c->48	m->5	
olz	m->2	
olä	m->5	
olö	s->2	
om 	"->7	-->10	1->5	2->3	3->6	4->4	5->1	6->1	A->9	B->12	C->4	D->7	E->99	F->9	G->8	H->7	I->6	J->4	K->6	L->8	M->4	N->1	O->1	P->9	R->3	S->8	T->12	V->1	W->3	a->528	b->217	c->6	d->680	e->339	f->395	g->160	h->369	i->289	j->155	k->302	l->133	m->300	n->152	o->117	p->103	r->231	s->391	t->156	u->157	v->458	y->4	Ö->4	ä->221	å->34	ö->33	
om!	T->1	
om"	.->1	
om)	 ->1	;->1	
om,	 ->58	
om-	 ->1	
om.	 ->2	A->1	D->10	E->2	H->2	I->1	J->7	M->4	N->1	O->1	S->2	V->3	
om/	r->1	
omI	.->1	
oma	d->1	g->1	n->3	r->30	t->19	
omb	 ->1	.->1	a->4	e->9	i->1	l->5	n->1	o->1	r->2	u->12	
omd	e->1	i->1	r->6	ö->2	
ome	d->21	n->24	r->10	s->1	t->2	u->4	
omf	a->83	l->1	o->4	å->2	ö->162	
omg	e->1	i->3	r->4	å->14	
omh	u->1	
omi	 ->20	,->2	.->3	?->1	e->8	n->41	s->242	
omk	r->15	
oml	a->1	i->18	o->2	ä->2	
omm	a->165	e->834	i->1253	o->3	u->33	ö->1	
omn	a->45	
omo	f->1	g->2	r->10	s->1	
omp	a->1	e->21	l->45	o->4	r->30	
omr	i->1	u->2	å->316	ö->42	
oms	 ->2	-->3	a->4	b->1	f->4	g->1	h->1	k->1	l->6	n->11	o->9	p->2	r->1	t->156	v->2	y->3	ä->8	
omt	a->1	ä->1	
omu	l->1	
omv	a->5	ä->12	
omá	n->1	
omä	s->1	
omå	l->3	
omé	 ->2	a->1	k->1	s->1	
omö	j->16	
on 	(->7	-->5	1->6	3->1	5->2	A->1	B->1	E->1	H->1	I->1	P->2	V->5	W->17	a->50	b->14	c->1	d->12	e->15	f->42	g->13	h->18	i->47	j->4	k->40	l->7	m->31	n->8	o->68	p->21	r->9	s->108	t->30	u->11	v->12	ä->12	å->5	ö->1	
on"	 ->1	
on)	 ->2	
on,	 ->72	
on-	 ->1	H->1	
on.	 ->4	1->1	A->1	B->1	D->22	E->3	F->5	G->1	H->7	I->7	J->14	K->2	L->1	M->4	N->2	O->3	S->5	T->2	U->1	V->16	Å->1	
on/	å->2	
on:	 ->3	
on;	 ->1	
on?	 ->2	D->1	J->1	K->3	V->1	Ä->1	
onN	ä->1	
ona	 ->26	d->7	k->1	l->158	n->2	p->2	r->8	s->3	t->6	z->2	
onb	e->1	l->15	
onc	e->40	i->2	k->14	
ond	 ->8	a->5	e->120	g->2	i->1	m->3	o->5	s->4	u->1	
one	 ->27	-->2	l->277	m->3	n->1516	r->591	t->8	
onf	e->172	i->4	l->16	r->1	
ong	e->1	i->2	r->1	s->1	
onh	u->1	
oni	 ->3	.->1	a->1	k->1	n->6	s->33	t->1	
onj	u->2	ä->1	
onk	r->58	u->285	
onl	a->1	i->34	
onm	ä->3	ö->2	
onn	a->1	ä->1	
ono	d->3	k->3	m->315	p->17	
onr	a->1	
ons	 ->11	-->4	a->12	b->2	d->8	e->68	f->23	h->9	i->13	k->14	l->12	m->7	n->2	o->4	p->12	r->17	s->17	t->122	u->75	v->1	ä->2	å->1	
ont	 ->2	.->1	a->29	e->17	i->63	o->7	r->193	
onv	e->29	i->4	
ony	m->5	
onz	á->1	
onä	r->248	
onå	r->1	
onö	d->11	
oo 	f->1	
ood	 ->1	f->1	s->1	w->1	
ooi	j->1	
ool	,->1	
oom	r->1	
oop	e->1	
oos	 ->1	
op 	a->1	b->1	d->1	f->1	o->2	p->1	s->2	t->1	u->1	ä->1	
op,	 ->6	
op-	s->1	
op.	D->1	I->1	J->1	S->1	
opa	 ->142	!->2	"->1	,->36	.->60	;->1	?->3	N->1	d->2	g->5	k->1	m->1	n->1	p->166	r->6	s->48	t->1	v->3	
ope	i->712	r->13	t->2	
opi	a->1	e->4	l->1	n->4	
opl	a->1	
opo	l->33	r->9	u->5	
opp	 ->16	,->1	.->1	a->107	e->19	l->7	m->12	n->12	o->7	
opr	a->1	o->7	
opt	i->8	
opu	l->7	
opy	r->1	
opå	 ->1	
opé	 ->1	e->9	
or 	-->3	F->1	M->2	T->3	a->100	b->23	c->1	d->31	e->12	f->41	g->7	h->19	i->59	j->26	k->7	l->4	m->27	n->6	o->88	p->24	r->6	s->110	t->26	u->24	v->21	ä->15	ö->2	
or)	 ->1	
or,	 ->83	
or.	 ->1	.->1	A->1	B->1	D->24	E->1	F->10	G->1	H->3	J->12	K->3	L->1	M->4	N->3	O->2	R->1	S->2	T->2	V->8	Ä->1	Ö->1	
or:	 ->4	
or;	 ->1	
or?	,->1	H->2	Ä->1	
ora	 ->158	,->2	.->3	?->1	d->5	l->8	n->1	r->4	t->33	
orb	e->2	i->1	r->15	
orc	e->1	y->4	
ord	 ->51	,->4	-->1	.->5	:->2	a->22	b->67	e->169	f->216	i->8	k->1	l->6	m->1	n->183	o->65	r->24	s->2	t->2	v->3	
ore	 ->30	a->5	b->1	d->1	g->1	l->1	n->69	r->50	s->1	t->3	
orf	ö->2	
org	 ->10	a->261	e->5	l->3	m->2	o->37	s->1	
orh	a->1	e->1	
ori	 ->6	a->10	e->31	g->2	k->7	m->5	n->10	s->51	t->106	u->10	
ork	 ->1	a->5	n->1	
orl	d->1	i->2	u->3	ä->1	
orm	 ->58	,->9	.->7	:->1	a->145	e->170	f->3	i->1	n->26	o->1	p->15	s->1	t->7	u->18	å->1	
orn	 ->22	)->1	,->12	.->10	?->1	a->99	e->1	o->2	s->4	
oro	 ->36	,->4	.->9	a->21	l->6	n->5	s->4	v->2	
orp	e->2	o->1	u->5	
orr	?->1	a->6	e->33	i->2	u->9	
ors	 ->54	,->7	.->11	a->37	b->1	d->8	e->7	i->1	k->44	l->3	t->3	ö->1	
ort	 ->262	)->1	,->26	-->3	.->21	:->1	?->1	N->1	a->9	b->3	d->1	e->131	f->100	g->6	i->9	k->2	l->1	m->2	n->2	o->15	p->2	s->143	u->100	v->1	y->1	
oru	m->6	
orv	 ->1	e->5	
orw	e->1	
orä	k->1	r->2	t->10	
orê	t->1	
orö	s->4	
os 	D->1	E->2	F->1	O->1	R->1	a->6	b->12	d->13	e->4	f->6	h->1	i->3	k->7	l->1	m->6	n->1	o->14	p->2	r->1	s->4	t->2	v->3	y->1	å->1	
os!	 ->1	
os,	 ->3	
osa	m->2	n->1	t->4	
ose	d->1	n->1	x->1	
osf	ä->1	
osi	o->1	t->87	v->1	
osj	u->1	
osk	e->3	o->3	r->1	v->1	y->1	
osl	a->1	ä->1	
osm	o->4	
osn	i->2	
oso	f->5	r->1	v->60	
osp	i->2	
oss	 ->289	,->15	.->18	:->1	?->2	a->2	e->2	i->3	n->1	t->1	
ost	 ->7	-->5	.->1	a->23	b->1	e->8	h->1	i->1	n->108	r->5	s->2	v->1	ä->4	
osv	.->6	
osy	n->1	s->4	
osä	k->12	t->5	
oså	r->1	
ot 	-->3	1->1	5->1	A->1	D->1	E->10	F->3	G->1	H->3	I->1	J->3	K->1	L->1	M->1	R->2	S->1	T->2	U->1	W->2	a->57	b->28	d->67	e->29	f->30	g->2	h->10	i->16	j->4	k->10	l->8	m->27	n->7	o->18	p->16	r->11	s->105	t->8	u->5	v->27	y->1	Ö->3	ä->3	å->2	ö->6	
ot!	 ->7	D->1	
ot,	 ->20	
ot.	 ->1	A->1	D->2	F->2	J->2	S->1	V->1	Ä->1	
ot?	N->1	
ota	 ->4	c->1	d->8	l->46	n->2	r->11	s->9	t->2	
otb	i->1	o->1	
ote	 ->1	k->6	l->1	n->36	r->38	s->10	t->8	
otf	u->1	ä->2	
otg	å->1	
oth	-->7	a->3	e->1	
oti	k->7	l->17	o->1	s->7	v->21	
otj	ä->1	
otn	i->17	
oto	 ->2	-->1	.->1	k->26	p->2	r->9	s->1	
otp	a->4	r->2	
otr	o->2	y->1	
ots	 ->64	a->23	p->2	t->16	v->17	y->1	ä->17	
ott	 ->54	,->11	.->11	a->27	e->147	g->1	i->1	l->5	m->1	n->4	o->1	s->33	
otu	l->1	m->1	r->1	s->1	
otv	e->6	i->3	
oty	d->4	
otä	n->1	
otå	l->1	t->3	
ou 	f->1	o->1	
ouc	h->12	
ouk	 ->1	
oul	a->1	o->5	
oum	b->4	
oun	c->1	d->6	
oup	 ->2	
our	a->8	g->5	i->1	l->6	n->3	s->1	
ous	e->1	k->1	
out	h->2	i->1	n->1	
oux	-->1	
ov 	a->16	f->4	i->2	k->1	n->1	o->7	p->9	s->3	t->8	
ov"	,->1	
ov,	 ->3	
ov.	 ->1	A->1	D->1	H->1	U->1	
ova	 ->2	d->4	k->1	n->10	r->2	t->13	
ove	m->11	n->7	r->11	t->38	
ovi	c->1	l->4	n->3	s->24	
ovj	e->1	
ovk	a->1	o->1	
ovo	 ->26	,->11	.->12	?->2	N->1	k->2	r->2	s->7	
ovs	i->1	k->2	m->5	t->1	
ovv	ä->2	
ovy	t->1	
ovä	c->3	d->2	l->1	n->1	r->15	s->1	
ovå	d->1	r->2	
ow 	t->1	
ow-	h->1	
owe	.->2	r->3	
owi	s->2	t->1	
own	 ->2	,->1	
ox 	o->1	s->1	
ox!	J->1	
ox,	 ->2	
oxa	l->5	
oxi	d->5	n->2	s->1	
oxn	i->1	
oya	l->1	
oyd	s->1	
oyo	l->2	
oäm	n->1	
oän	d->4	g->12	
oår	 ->1	
oön	s->1	
oöv	e->6	
p (	k->2	
p ,	 ->1	
p -	 ->3	
p C	a->1	
p E	u->1	
p J	ö->1	
p T	i->1	
p a	l->7	n->5	t->11	v->77	
p b	e->3	i->1	å->1	ö->2	
p d	e->44	o->1	ä->3	
p e	f->3	l->3	n->12	t->6	x->1	
p f	o->1	r->15	u->1	å->1	ö->21	
p g	e->2	r->2	
p h	a->7	e->1	u->1	ä->3	ö->1	
p i	 ->32	d->1	g->4	n->10	
p k	a->1	o->7	
p l	a->1	i->1	ä->3	
p m	a->1	e->11	o->4	å->2	
p n	a->1	i->1	y->1	ä->1	å->3	
p o	c->23	l->1	m->8	r->2	
p p	e->1	o->1	r->3	å->13	
p r	e->2	ä->3	å->1	ö->1	
p s	a->1	i->3	j->1	k->7	o->21	t->2	ä->2	å->2	
p t	i->18	o->1	r->1	v->1	y->2	
p u	n->3	p->1	t->8	
p v	a->4	i->4	ä->2	
p ä	n->3	r->11	v->1	
p ö	n->1	v->1	
p" 	f->1	
p"!	I->1	
p",	 ->2	
p, 	A->3	E->1	a->2	b->1	d->5	e->8	f->3	g->1	h->3	i->2	j->1	l->1	m->4	n->1	o->7	p->1	r->1	s->3	u->1	v->3	ä->1	
p-s	h->1	
p. 	S->1	s->1	t->1	
p..	(->1	
p.A	h->1	
p.D	a->1	e->15	
p.E	f->1	u->1	
p.F	a->1	
p.H	ä->1	
p.I	 ->3	n->1	
p.J	a->12	
p.M	e->1	
p.P	å->1	
p.S	j->1	l->1	o->1	
p.T	i->1	
p.V	i->8	
p.g	.->1	
p.Ä	n->1	v->1	
p: 	K->1	
p?H	u->1	
pa 	-->3	O->1	W->1	a->22	b->8	d->33	e->52	f->29	g->5	h->16	i->23	j->1	k->23	l->2	m->29	n->12	o->29	p->11	r->8	s->45	t->25	u->8	v->10	y->1	ä->12	å->1	ö->1	
pa!	A->1	F->1	
pa"	.->1	
pa,	 ->39	
pa.	.->2	1->1	D->15	E->3	F->3	H->6	I->2	J->8	K->1	M->3	N->1	O->1	P->1	R->1	T->2	U->1	V->10	Ä->1	
pa;	 ->1	
pa?	H->1	V->2	
paN	ä->1	
pac	i->5	k->5	
pad	 ->3	e->24	
pag	a->3	e->1	n->1	r->1	
pak	e->7	o->1	t->5	
pal	e->12	
pam	i->1	
pan	 ->2	,->1	d->64	e->1	i->8	j->7	s->12	t->1	
pap	a->166	p->5	
par	 ->74	.->3	a->26	c->1	e->11	i->4	k->14	l->558	n->1	s->1	t->148	å->1	
pas	 ->200	,->5	.->10	:->1	?->1	s->33	t->11	
pat	 ->14	.->1	:->1	e->1	i->13	j->1	r->1	s->9	
pav	a->3	
pay	a->2	
pba	c->1	
pbr	i->3	
pby	g->20	
pbä	r->1	
pbå	d->1	
pda	t->3	
pde	l->3	
pdr	a->22	
pe 	i->1	p->1	
pea	n->1	u->1	
pec	i->85	
ped	a->1	i->1	o->1	
peg	l->12	n->1	
peh	å->13	
pei	s->712	
pek	a->70	t->148	u->4	
pel	 ->77	,->7	.->5	:->3	;->1	a->46	e->2	l->1	n->1	p->1	r->5	v->28	
pen	 ->218	,->26	.->33	:->2	?->1	N->1	b->36	c->1	d->6	g->55	h->62	i->1	n->11	s->110	t->1	u->1	
per	 ->119	,->9	.->12	:->2	a->22	e->2	f->7	i->94	l->1	m->8	n->50	o->1	r->1	s->123	t->46	
pes	 ->2	k->1	s->2	t->5	
pet	 ->102	)->1	,->18	.->7	?->1	e->11	i->1	s->17	
pfa	l->1	n->1	t->51	
pfy	l->54	
pfö	d->1	l->10	r->13	
pgi	c->3	f->77	
pgo	d->1	
pgr	a->1	
pgå	 ->1	e->7	n->2	r->5	
pgö	r->2	
pha	r->1	
phe	r->3	t->4	
pho	v->13	
pht	a->1	
phä	n->1	v->5	
phå	l->3	
phö	j->1	r->9	
pia	 ->1	
pic	 ->1	e->1	
pie	l->8	n->3	r->1	
pil	l->1	o->4	
pin	 ->1	i->4	
pio	n->1	
pir	a->1	e->3	
pis	k->2	
pit	 ->2	a->27	e->6	u->2	
pja	k->1	
pka	y->11	
pko	l->1	m->6	
pkr	a->1	
pla	 ->1	c->17	d->1	n->132	r->2	s->8	t->45	
ple	m->11	n->12	t->17	v->17	x->4	
pli	c->13	g->104	k->33	m->5	n->17	t->4	v->1	
plo	m->11	s->2	
plu	n->1	r->1	s->2	
ply	s->4	
plä	d->2	
plå	d->11	g->1	n->3	
plö	s->4	t->4	
pma	n->58	
pmj	u->2	
pmu	n->21	
pmä	r->53	t->2	
pmö	t->12	
pna	 ->9	,->2	d->3	r->3	s->2	
pne	n->2	
pni	n->119	
pnå	 ->49	,->1	.->4	d->6	r->13	s->7	t->13	
po,	 ->1	
poe	t->1	
pok	 ->1	,->1	e->2	
pol	 ->15	,->3	-->1	.->2	;->1	a->1	e->2	f->3	i->557	k->1	s->4	
pon	d->1	e->12	s->2	t->4	
poo	l->1	
pop	u->7	
por	,->1	d->1	n->2	s->1	t->317	ä->2	
pos	 ->1	i->87	t->15	
pot	e->8	i->5	s->1	
pou	l->5	
poä	n->12	
pp 	(->2	-->2	E->1	T->1	a->24	b->4	d->42	e->21	f->25	g->3	h->12	i->30	k->7	l->5	m->9	n->5	o->11	p->16	r->6	s->18	t->16	u->9	v->7	ä->9	
pp,	 ->24	
pp.	.->1	A->1	D->5	F->1	J->7	M->1	P->1	V->3	Ä->2	
pp?	H->1	
ppa	 ->17	d->8	n->2	r->4	s->109	
ppb	a->1	r->3	y->20	ä->1	å->1	
ppd	a->3	e->3	r->22	
ppe	 ->1	h->13	l->1	n->178	r->70	t->35	
ppf	a->52	y->54	ö->24	
ppg	i->80	r->1	å->8	ö->2	
pph	e->4	o->13	ä->6	ö->10	
ppj	a->1	
ppk	o->7	
ppl	a->6	e->17	i->3	y->4	å->11	ö->4	
ppm	a->58	j->2	u->21	ä->55	ö->12	
ppn	a->16	i->17	å->93	
ppo	n->3	r->115	s->2	
ppr	e->54	i->6	o->5	u->1	y->1	ä->39	ö->5	
pps	 ->4	a->7	b->2	k->29	p->2	r->3	s->3	t->39	v->2	ä->3	
ppt	 ->5	a->10	e->3	i->1	o->2	r->10	ä->11	
ppu	n->1	
ppv	e->2	i->6	ä->2	
ppy	 ->1	
pra	c->1	g->1	k->33	n->1	t->5	x->8	
pre	c->43	f->3	j->4	l->3	m->10	n->5	p->52	r->1	s->81	
pri	c->3	d->20	k->6	l->3	m->1	n->195	o->38	s->28	v->28	
pro	b->174	c->201	d->76	f->10	g->238	j->62	k->1	m->22	n->1	p->19	s->1	t->37	v->18	
pru	n->19	s->1	
pry	c->1	
prä	c->2	g->5	k->1	n->1	t->36	
prå	k->24	n->2	
prö	r->5	v->15	
ps 	a->1	f->1	u->1	v->3	
ps-	 ->1	
ps.	J->1	M->1	
psa	m->4	t->3	v->2	
psb	e->4	r->1	y->1	
psd	i->1	
psf	r->1	
psi	n->15	s->1	
psk	a->23	h->1	j->4	o->5	ä->2	
psl	a->5	
psm	a->2	e->1	ä->16	å->1	
psn	i->11	
pso	n->1	r->1	
psp	e->2	o->2	r->3	å->2	
psr	a->1	e->11	ä->9	
pss	t->4	y->1	ä->2	
pst	o->4	ä->3	å->32	
psv	a->2	
psy	k->1	
psä	g->1	t->2	
pså	t->2	
pt 	b->2	d->2	e->2	f->1	i->3	k->1	o->1	s->2	t->2	u->5	v->1	ö->1	
pt.	D->1	H->1	
pta	 ->2	.->1	b->37	g->7	n->7	r->1	s->2	
pte	 ->6	m->15	n->4	r->45	s->2	t->3	
pti	k->3	l->1	m->7	o->14	s->5	
pto	g->4	m->1	
ptr	ä->10	
ptä	c->11	
pub	l->26	
pul	a->1	i->4	s->6	ä->2	
pum	p->2	
pun	d->4	k->342	
pur	i->1	
pus	 ->5	
pve	r->2	
pvi	g->1	l->1	s->5	
pvä	g->1	r->1	
py 	e->1	
pyr	a->1	i->1	
pän	n->11	
pär	r->3	
på 	-->5	1->4	2->4	3->3	4->1	5->3	7->2	8->3	9->2	A->3	B->7	C->2	E->18	F->1	G->2	H->1	I->9	M->1	O->1	P->1	R->3	T->1	V->2	a->205	b->40	c->3	d->314	e->224	f->96	g->106	h->23	i->26	j->7	k->50	l->34	m->77	n->64	o->38	p->23	r->49	s->126	t->50	u->16	v->90	y->1	z->1	Ö->2	ä->9	å->7	ö->8	
på,	 ->16	
på.	B->1	D->4	E->2	J->3	N->1	O->1	U->1	V->1	Ä->2	
på:	 ->3	
på?	.->1	J->1	
påb	j->1	ö->11	
påd	r->1	
påf	r->1	ö->4	
påg	i->3	å->18	
pål	a->1	e->1	i->1	ä->1	
påm	i->30	
påp	e->50	
pår	 ->4	,->2	a->4	e->1	n->2	
pås	k->7	t->21	
påt	a->9	r->3	v->4	
påv	e->37	i->3	
pé 	o->1	
pée	r->9	
pér	y->1	
pök	e->3	s->1	
qal	 ->2	
qua	 ->2	l->8	
que	 ->1	,->1	s->5	
qui	e->1	n->1	o->1	s->1	t->1	
quo	 ->1	,->1	
quq	a->2	
r "	K->1	a->2	f->1	i->1	k->1	n->1	ö->1	
r (	C->4	F->1	a->1	i->1	
r -	 ->86	,->1	
r 1	 ->2	,->2	/->1	0->4	2->2	3->1	5->2	6->1	7->3	9->72	
r 2	 ->1	0->64	5->1	6->1	7->2	8->1	9->3	
r 3	 ->1	-->1	0->2	1->1	2->2	3->3	5->2	6->1	7->1	8->1	9->1	
r 4	 ->1	0->4	1->1	2->1	3->1	4->1	5->1	6->1	
r 5	 ->3	,->1	0->2	
r 6	 ->1	0->1	
r 7	 ->2	.->1	3->1	5->1	6->1	
r 8	 ->1	0->4	1->1	
r 9	 ->1	0->2	7->2	
r A	g->1	l->8	m->2	n->1	r->1	z->1	
r B	N->2	S->1	a->13	e->6	i->1	o->5	r->6	
r C	E->1	S->1	e->2	o->5	
r D	a->3	e->1	o->1	u->1	
r E	C->1	G->7	M->2	U->18	g->1	h->1	k->1	l->1	r->3	u->112	v->3	x->1	
r F	N->3	P->2	a->1	i->1	l->1	o->2	r->2	ö->6	
r G	A->1	a->2	e->1	o->4	r->2	u->2	
r H	a->1	e->1	i->1	ä->2	
r I	 ->1	-->1	I->4	M->1	N->1	n->2	s->5	t->1	
r J	a->1	o->3	ö->2	
r K	a->3	i->11	o->3	u->3	v->1	y->1	
r L	a->10	e->1	i->1	o->2	u->1	y->2	
r M	a->4	e->1	o->17	
r N	a->1	e->1	i->3	o->1	
r O	F->1	L->2	r->1	s->1	
r P	P->1	V->1	a->23	o->10	r->2	
r R	E->1	a->2	e->2	h->1	o->1	u->1	å->1	
r S	a->2	c->6	e->5	h->1	k->1	o->2	p->1	w->1	y->2	ã->1	
r T	a->3	e->1	h->1	i->6	o->1	s->2	u->4	
r U	C->1	N->1	S->2	r->1	
r V	i->5	o->1	
r W	T->1	a->4	y->1	
r [	S->1	
r a	b->14	c->6	d->1	g->1	i->1	k->12	l->291	m->4	n->196	r->43	s->5	t->1979	u->1	v->252	
r b	a->44	e->269	i->47	j->1	l->43	o->18	r->53	u->22	y->9	ä->16	å->11	ö->30	
r c	a->10	e->4	h->2	i->8	o->2	
r d	a->18	e->2212	i->42	j->10	o->48	r->16	u->6	y->2	ä->105	å->29	ö->8	
r e	c->2	d->1	f->46	g->18	j->8	k->28	l->62	m->37	n->675	r->76	t->313	u->31	v->3	x->27	
r f	a->81	e->16	i->42	j->1	l->29	o->60	r->296	u->26	y->4	ä->2	å->53	ö->760	
r g	a->15	e->110	i->15	j->49	l->19	o->29	r->63	u->2	y->3	ä->8	å->28	ö->27	
r h	a->218	e->123	i->19	j->10	o->32	u->51	y->2	ä->55	å->14	ö->28	
r i	 ->552	.->1	a->1	b->3	c->2	d->7	f->6	g->13	h->4	k->1	l->4	m->1	n->717	r->1	s->2	t->6	v->1	
r j	a->285	o->17	u->59	ä->8	
r k	a->89	e->1	l->36	n->8	o->468	r->39	u->48	v->20	ä->23	ö->3	
r l	a->63	e->49	i->82	o->13	u->4	y->23	ä->69	å->37	ö->15	
r m	a->200	e->371	i->226	o->54	u->2	y->109	ä->32	å->95	ö->46	
r n	a->47	e->16	i->56	o->20	u->46	y->27	ä->110	å->110	ö->45	
r o	a->9	b->7	c->732	e->9	f->39	j->1	k->4	l->19	m->306	n->2	p->1	r->51	s->135	t->5	u->5	v->2	ö->1	
r p	a->62	e->48	l->15	o->34	r->88	u->10	å->334	
r r	a->17	e->179	i->30	o->8	u->6	y->1	ä->77	å->50	ö->26	
r s	a->121	e->78	i->218	j->33	k->172	l->19	m->9	n->15	o->644	p->30	t->210	u->6	v->30	y->43	ä->95	å->104	ö->4	
r t	.->3	a->382	e->11	i->439	j->15	o->17	r->70	u->7	v->40	y->36	ä->8	å->1	
r u	n->121	p->129	r->10	t->250	
r v	a->175	e->75	i->632	o->3	u->3	ä->77	å->90	
r y	n->1	p->1	r->2	t->16	
r Ö	V->1	s->7	
r ä	g->8	l->4	m->3	n->115	r->150	v->35	
r å	 ->2	k->1	l->1	r->36	s->6	t->59	
r ö	a->1	d->1	g->7	k->13	n->7	p->16	r->2	s->3	v->122	
r! 	1->1	A->1	B->2	C->1	D->20	E->10	F->8	G->2	H->1	I->9	J->26	K->1	L->4	M->1	N->4	O->1	P->2	S->3	T->5	U->2	V->11	Ä->3	Å->1	
r!"	D->1	O->1	
r!.	H->1	
r!D	e->7	
r!E	f->1	r->1	
r!J	a->5	
r!M	e->1	i->1	y->1	
r!T	i->1	
r!V	i->2	
r" 	h->1	m->2	o->1	s->2	
r")	,->1	
r",	 ->1	
r".	D->1	J->1	O->1	
r) 	B->1	V->1	o->3	
r).	)->1	
r)?	 ->1	
r)F	r->2	
r)J	a->1	
r)K	o->1	
r)T	a->1	
r, 	"->1	(->1	1->1	B->1	E->1	G->1	M->1	P->1	T->2	W->1	a->60	b->21	d->48	e->38	f->56	g->12	h->34	i->50	j->12	k->49	l->16	m->103	n->25	o->134	p->14	r->9	s->123	t->31	u->43	v->46	ä->37	å->7	ö->1	
r- 	o->4	s->1	
r-b	i->1	
r-k	o->1	
r-n	a->1	
r-p	r->11	
r-r	e->1	
r. 	(->1	A->1	D->7	E->5	F->1	H->1	J->2	M->3	N->1	S->2	T->1	V->2	i->1	Ä->1	
r.(	A->1	I->1	L->1	
r.)	 ->1	S->1	
r.-	 ->4	
r..	 ->4	(->3	.->2	H->1	V->1	
r.9	0->1	
r.A	l->4	m->1	n->1	t->4	v->4	
r.B	a->2	e->7	l->2	o->1	r->1	
r.C	S->1	
r.D	a->1	e->226	i->1	o->1	ä->14	å->2	
r.E	U->2	f->5	n->14	r->1	t->6	u->7	x->1	
r.F	P->1	e->1	o->1	r->13	å->1	ö->43	
r.G	e->7	ö->1	
r.H	a->1	e->25	u->3	ä->8	
r.I	 ->30	n->9	t->1	
r.J	a->119	
r.K	a->3	i->1	o->27	r->1	v->1	ä->1	
r.L	a->1	i->3	y->1	å->6	
r.M	a->6	e->29	i->4	y->1	ä->1	
r.N	a->4	i->2	u->1	y->1	ä->10	å->1	
r.O	b->1	c->8	m->17	r->2	
r.P	a->2	l->1	r->3	u->1	å->3	
r.R	a->1	e->5	i->1	ä->1	å->3	
r.S	a->5	e->2	k->1	l->2	o->7	t->5	å->5	
r.T	a->5	e->1	i->15	r->1	y->3	
r.U	n->7	t->1	
r.V	a->14	e->2	i->88	å->5	
r.k	o->1	
r.Ä	n->5	r->3	v->5	
r.Å	 ->2	
r.Ö	V->1	
r: 	"->1	A->1	D->3	F->3	I->1	K->1	O->1	P->1	V->2	a->4	d->8	e->2	f->3	h->1	i->1	k->1	n->1	o->2	t->1	u->1	v->5	Ä->1	
r; 	a->1	d->4	e->1	i->2	j->1	m->1	o->2	v->2	
r?,	 ->1	
r?-	 ->1	
r?.	 ->1	
r?B	o->1	
r?D	e->2	ä->1	
r?E	u->1	
r?F	r->2	
r?H	a->2	e->3	u->1	
r?I	 ->2	
r?J	a->3	
r?K	a->1	o->2	
r?M	e->2	
r?N	a->1	i->1	ä->1	
r?P	å->1	
r?S	o->1	
r?T	a->1	
r?V	e->1	i->2	
r?Ä	r->2	v->1	
rHe	r->1	
rJa	g->1	
rMe	d->1	
rNä	s->2	
ra 	"->2	-->6	1->4	2->2	5->2	7->1	A->1	B->1	D->1	E->18	F->2	I->3	J->1	L->3	R->2	T->2	a->228	b->86	c->4	d->288	e->305	f->265	g->80	h->71	i->107	j->6	k->181	l->69	m->217	n->83	o->175	p->137	r->77	s->291	t->126	u->69	v->114	y->7	Ö->3	ä->54	å->53	ö->28	
ra!	 ->1	M->1	
ra"	.->2	
ra,	 ->73	
ra.	 ->1	A->2	B->1	D->16	E->6	F->2	H->3	I->3	J->15	L->3	M->5	N->4	O->1	P->4	S->2	U->1	V->5	
ra:	 ->7	
ra;	 ->2	
ra?	A->1	D->1	J->1	
rab	b->50	e->5	i->6	l->1	r->1	s->2	v->1	
rac	a->3	k->1	o->1	
rad	 ->122	,->3	.->8	e->262	i->37	o->6	v->3	
rae	l->58	
raf	 ->1	a->1	f->41	i->23	r->2	t->149	
rag	 ->61	,->2	.->6	:->1	a->115	e->155	i->18	m->1	n->49	r->3	s->21	
rah	a->1	u->1	
rai	n->2	
rak	 ->10	,->1	.->3	?->1	a->4	e->3	i->1	o->5	r->1	s->3	t->94	
ral	 ->13	,->1	-->6	.->2	a->45	b->8	d->18	e->6	f->1	i->44	l->15	s->2	t->11	
ram	 ->293	,->28	.->29	?->2	a->18	e->62	f->146	g->53	h->24	i->1	k->11	l->21	m->109	n->2	p->25	r->1	s->50	t->117	u->1	v->4	å->22	ö->2	
ran	 ->37	,->4	-->1	.->6	?->2	a->1	b->8	c->5	d->812	g->6	i->3	k->43	l->2	n->10	o->1	s->237	t->108	v->22	z->3	ç->1	
rao	r->1	
rap	e->1	p->109	r->1	
rar	 ->433	!->21	,->31	.->13	:->1	;->1	a->1	b->2	e->47	k->4	l->1	n->17	s->1	t->3	v->5	
ras	 ->329	!->2	,->23	.->48	;->1	a->4	b->5	c->3	e->1	h->1	i->27	k->1	m->1	s->3	t->38	
rat	 ->126	,->14	.->14	;->1	a->10	e->102	i->257	o->9	s->45	t->2	u->53	ö->2	
rau	m->1	
rav	 ->48	,->4	.->6	?->1	a->3	e->48	t->1	
rax	 ->3	i->8	
ray	,->1	
raç	a->5	
rb,	 ->1	
rba	-->1	l->1	n->4	r->20	s->1	y->1	
rbe	d->1	g->1	h->6	l->3	m->1	r->35	s->2	t->576	
rbi	 ->1	f->2	g->6	h->1	l->1	n->22	s->7	
rbj	u->33	ö->1	
rbl	e->1	i->15	å->2	
rbr	i->15	o->1	u->1	y->5	ä->2	
rbu	d->26	n->12	
rbä	t->78	
rbö	l->1	r->11	
rce	 ->1	l->2	n->1	
rco	u->1	
rcy	k->4	
rd 	-->1	2->1	C->1	I->2	K->1	a->11	b->2	d->2	e->5	f->10	g->1	i->7	j->1	k->6	m->5	n->1	o->19	p->2	s->12	t->5	u->1	v->6	
rd)	,->1	
rd,	 ->18	
rd-	a->1	f->1	
rd.	B->1	D->6	E->1	H->1	I->1	J->1	U->1	V->2	
rd:	 ->2	
rd;	 ->3	
rda	 ->64	,->5	.->4	?->1	d->3	g->7	l->6	m->45	n->17	r->10	s->4	t->4	
rdb	r->57	ä->10	
rde	 ->137	,->3	-->2	.->8	a->1	d->2	f->7	g->3	l->47	m->1	n->64	r->294	s->18	t->27	u->1	
rdf	ö->223	
rdh	e->1	
rdi	g->41	n->1	r->2	s->13	t->1	
rdj	u->11	
rdk	u->1	
rdl	a->1	i->8	
rdm	å->1	
rdn	a->31	i->155	
rdo	 ->1	m->11	n->65	r->2	
rdr	a->182	e->1	i->19	ö->1	
rds	 ->1	-->1	b->1	k->1	l->3	m->2	o->1	p->7	s->3	t->3	u->1	v->1	
rdt	i->1	y->1	
rdu	b->2	n->1	
rdv	r->1	ä->2	
rdä	r->4	
rdö	m->20	r->1	
re 	-->5	1->2	2->2	3->1	4->1	A->1	B->1	D->2	E->2	H->1	K->1	a->64	b->46	c->1	d->30	e->38	f->127	g->21	h->35	i->59	j->3	k->61	l->11	m->121	n->18	o->74	p->42	r->21	s->127	t->51	u->33	v->40	ä->58	å->9	ö->11	
re!	S->1	
re"	 ->2	,->1	
re,	 ->88	
re-	A->1	
re.	 ->3	A->2	B->1	D->23	E->5	F->3	H->1	I->5	J->8	K->2	M->8	N->2	P->2	R->2	S->3	T->3	U->1	V->7	Ä->5	
re:	 ->2	
re?	D->1	K->1	O->1	V->1	
rea	 ->4	g->16	k->21	l->18	m->8	t->3	
reb	e->3	i->1	o->1	r->2	y->23	
rec	i->50	k->1	o->1	t->1	y->1	
red	 ->19	,->1	.->4	a->187	d->38	e->17	g->1	i->4	j->73	l->10	n->8	o->17	r->166	s->67	u->4	ö->2	
ree	-->2	.->1	l->4	
ref	a->20	e->7	l->7	o->134	t->13	u->1	ö->1	
reg	e->332	i->276	l->126	r->1	å->17	
reh	a->2	
rei	s->1	
rej	u->4	ä->3	
rek	e->1	i->6	l->17	o->75	r->1	t->284	v->1	
rel	a->27	e->10	i->34	l->56	s->28	ä->2	
rem	a->2	e->1	h->14	i->21	o->19	s->3	t->4	å->14	
ren	 ->220	)->2	,->41	.->39	;->1	?->3	a->48	d->44	g->5	h->24	i->22	k->8	l->9	o->3	s->556	t->58	z->19	ö->3	
rep	 ->1	a->57	n->1	p->25	r->26	u->18	
rer	 ->77	!->1	,->17	.->16	a->88	i->19	n->41	o->1	s->1	ö->1	
res	 ->22	,->3	a->22	e->57	i->10	k->28	l->104	o->105	p->96	s->144	t->42	u->161	ä->1	
ret	 ->113	,->11	.->19	:->1	a->249	e->14	i->4	o->3	r->85	s->16	t->17	
reu	r->1	s->1	t->4	
rev	 ->10	.->1	i->35	l->4	o->1	s->3	
rex	t->6	
rey	 ->3	e->3	
rez	,->1	
rfa	l->4	r->105	t->7	
rfe	k->7	
rfi	n->4	r->2	s->1	
rfj	o->1	
rfl	u->14	y->6	ö->1	
rfo	d->4	g->18	n->58	r->29	
rfr	y->1	å->13	
rfu	n->2	
rfä	k->1	r->3	
rfå	n->1	
rfö	l->10	r->358	
rg 	H->14	a->1	f->2	g->1	i->1	k->1	m->2	o->8	s->1	t->1	u->1	ö->1	
rg,	 ->6	
rg.	D->1	J->1	L->1	V->1	
rga	 ->1	d->1	n->98	r->171	v->2	
rge	 ->4	,->1	n->7	r->25	s->3	
rgh	.->1	
rgi	 ->13	,->2	-->1	.->5	a->7	b->3	c->1	e->4	f->7	i->1	k->39	m->2	n->10	o->2	p->7	s->13	v->8	z->5	ä->1	å->1	
rgl	i->3	ö->2	
rgm	ä->2	
rgn	e->1	
rgo	 ->1	n->37	t->1	
rgr	i->14	u->4	ä->4	
rgs	f->1	
rgu	m->17	
rgä	l->1	v->1	
rgå	 ->1	n->12	r->6	t->1	
rgö	r->17	
rha	n->98	s->3	v->1	
rhe	a->1	t->308	u->2	
rhi	n->31	s->1	
rho	l->4	p->12	
rhu	n->7	s->3	
rhä	m->2	n->3	
rhå	g->2	l->70	
rhö	g->2	l->4	r->12	
ri 	-->1	1->4	2->5	8->2	L->3	V->1	a->1	b->1	d->1	e->2	f->5	i->7	k->3	m->3	n->2	o->12	r->8	s->8	v->2	ä->2	ö->2	
ri!	H->1	
ri,	 ->21	
ri-	 ->10	
ri.	B->1	H->1	J->1	L->1	M->1	V->1	
ria	 ->32	,->4	.->2	l->23	n->3	s->3	t->5	
rib	e->4	l->6	u->1	
ric	h->6	i->2	k->7	
rid	 ->10	,->1	.->1	a->20	d->2	e->26	i->32	l->1	n->15	o->2	s->4	
rie	 ->1	-->1	f->1	l->21	n->41	r->60	s->1	t->13	
rif	e->6	i->2	r->6	t->30	
rig	 ->59	"->1	,->4	.->1	a->71	e->59	h->54	i->2	j->1	o->4	s->2	t->47	ö->5	
rih	a->2	e->116	
rik	 ->7	,->2	.->2	a->88	e->185	i->49	l->2	o->2	t->250	
ril	 ->3	.->1	a->2	i->1	j->1	o->1	
rim	i->28	l->23	m->1	s->8	å->1	
rin	 ->41	!->1	,->15	.->15	:->1	?->1	c->194	d->2	f->4	g->1193	h->6	i->1	n->1	o->7	r->15	s->18	t->6	ä->3	
rio	 ->2	d->86	r->40	t->3	
rip	a->37	e->19	i->2	l->6	n->1	o->3	s->1	
rir	r->1	
ris	 ->21	,->2	.->2	:->1	?->1	a->1	d->5	e->37	f->1	k->146	l->2	m->30	n->1	o->4	s->3	t->113	u->1	
rit	 ->74	a->18	e->185	i->52	l->1	o->17	r->1	t->24	
riu	m->12	t->1	
riv	a->57	b->1	e->43	i->27	k->3	n->9	s->15	
riä	r->4	
riè	r->1	
riö	s->8	
rja	 ->68	d->10	n->19	r->17	t->12	
rjd	e->1	
rje	 ->91	r->2	
rjn	i->4	
rk 	-->2	a->1	b->2	d->1	e->3	f->5	g->1	h->1	i->11	k->5	l->1	m->3	o->7	p->5	s->9	t->3	u->1	v->4	ä->2	
rk,	 ->7	
rk-	d->1	
rk.	B->1	D->3	F->1	J->1	S->1	V->1	
rk?	R->1	
rka	 ->91	,->5	.->1	d->2	n->36	p->1	r->131	s->30	t->24	
rkb	a->3	o->1	
rkd	a->1	
rke	 ->8	f->1	l->6	n->31	p->1	r->17	s->18	t->42	
rki	.->1	e->35	l->1	n->2	s->7	v->2	
rkk	i->2	
rkl	a->85	i->210	y->1	ä->1	
rkm	e->2	
rkn	a->191	i->38	
rko	g->1	l->1	m->8	n->3	p->1	r->4	t->7	v->1	
rkr	a->1	o->1	ä->1	
rks	 ->5	.->3	a->105	t->19	
rkt	 ->42	,->1	.->2	a->18	s->1	y->8	
rku	l->3	n->2	r->1	
rkä	n->42	
rkö	t->1	
rl 	H->1	o->1	v->3	
rl-	H->1	
rla	g->14	m->600	n->31	
rld	 ->2	,->2	.->1	e->37	s->17	
rle	d->2	g->2	k->2	v->10	
rli	g->420	k->46	n->9	s->2	t->10	v->21	
rlo	r->20	
rls	r->2	
rlu	n->3	s->10	
rly	s->2	
rlä	g->11	k->1	m->18	n->40	r->1	t->18	
rlå	t->15	
rlö	s->2	
rlø	n->2	
rm 	a->26	b->1	d->2	e->5	f->3	i->3	j->1	k->4	l->1	o->3	p->1	s->7	v->3	ä->1	ö->1	
rm,	 ->9	
rm-	e->1	
rm.	D->1	E->1	M->1	N->1	S->1	V->1	Ä->1	
rm:	 ->1	
rma	 ->29	.->1	c->1	d->5	j->1	k->1	l->11	n->18	r->43	s->16	t->84	
rme	d->52	l->17	n->26	r->134	
rmf	ä->1	ö->2	
rmi	d->12	n->12	s->2	
rmn	i->31	
rmo	,->1	d->14	n->19	r->1	u->1	
rmp	a->1	r->14	
rmr	a->2	
rms	i->2	t->2	
rmt	 ->19	
rmu	l->18	
rmy	n->15	
rmä	s->1	
rmå	 ->2	g->31	l->1	n->14	r->1	t->1	
rmé	 ->1	n->2	
rmö	g->1	t->2	
rn 	(->1	-->4	E->2	b->2	d->2	e->3	f->10	g->1	h->3	i->6	k->5	l->2	m->1	n->1	o->16	p->1	r->1	s->12	t->2	u->2	v->2	ä->3	
rn)	.->1	
rn,	 ->24	
rn-	 ->2	
rn.	)->1	.->1	D->8	F->3	H->2	J->2	K->1	M->1	O->1	V->1	Ö->1	
rn/	N->2	
rn?	A->1	
rna	 ->1405	!->3	"->3	,->221	.->269	/->1	:->3	;->4	?->12	H->1	d->1	g->1	l->2	m->1	n->6	r->6	s->219	t->94	
rnb	a->1	
rnd	 ->3	
rne	 ->1	,->1	a->1	d->2	k->8	n->8	r->4	t->11	
rnf	r->3	
rnh	i->1	
rni	e->14	n->27	s->24	t->1	v->1	é->1	
rnk	a->1	r->22	
rno	g->2	
rnp	o->2	r->2	u->2	
rns	 ->18	t->2	ä->3	
rnt	 ->4	.->1	e->3	u->1	
rnu	f->14	
rnv	a->8	ä->15	
rny	a->4	b->39	e->6	
rnä	t->1	
rnö	d->1	r->1	
ro 	-->2	1->1	E->1	a->4	b->2	d->2	f->11	h->1	i->6	l->1	m->2	n->5	o->6	p->6	s->12	t->3	u->1	v->1	ä->4	ö->1	
ro!	A->1	
ro,	 ->15	
ro-	r->1	
ro.	A->1	B->1	D->3	F->2	H->1	J->2	K->1	N->1	O->1	S->1	T->1	V->3	
roa	 ->3	d->5	k->12	n->10	r->5	t->1	
rob	l->183	
roc	e->204	k->1	
rod	a->9	d->9	e->2	i->28	u->84	
roe	d->14	k->5	n->127	
rof	 ->24	,->4	.->4	a->1	d->1	e->59	h->1	i->4	s->4	ö->1	
rog	 ->5	a->3	b->1	e->3	k->1	r->240	s->2	
roi	s->1	
roj	e->64	k->1	u->6	
rok	 ->6	,->3	i->2	l->1	r->2	
rol	,->1	.->1	e->1	i->18	l->246	ä->2	
rom	 ->2	,->1	a->1	e->10	i->22	r->3	s->6	
ron	 ->13	,->3	-->1	a->1	g->1	i->12	j->1	m->2	o->4	s->3	t->4	
roo	m->1	
rop	 ->3	,->1	.->1	a->477	e->713	o->25	p->2	r->1	å->1	é->10	
ror	 ->179	,->4	.->5	?->1	d->49	e->28	i->10	n->6	s->6	
ros	 ->4	a->1	e->1	k->3	m->4	s->4	t->4	
rot	.->1	a->13	e->13	f->1	h->1	n->17	o->26	s->64	t->62	u->2	
rou	k->1	p->1	x->1	
rov	 ->16	"->1	,->1	.->2	a->3	e->7	i->6	k->2	s->4	ä->18	
rpa	 ->6	c->5	r->3	s->3	
rpe	g->1	r->1	t->2	
rpl	a->1	i->21	
rpn	i->1	
rpo	l->21	p->1	s->2	
rpr	e->1	i->1	o->4	
rpt	 ->2	a->2	
rpu	s->5	
rpå	 ->2	
rqu	i->1	
rr 	A->1	B->10	C->3	E->2	F->1	G->2	H->2	J->1	K->6	L->1	M->1	N->1	P->8	R->1	S->5	W->1	a->1	b->3	d->4	e->2	f->8	g->2	h->6	i->5	k->85	l->15	m->2	n->1	o->7	p->3	r->12	s->4	t->320	v->3	ä->5	å->1	ö->1	
rr,	 ->4	
rr.	V->1	
rr?	V->1	
rra	 ->48	d->2	i->2	n->9	r->50	s->3	t->4	
rre	 ->85	,->1	c->1	f->1	g->6	k->27	n->285	p->3	r->5	s->6	y->3	z->1	
rrg	å->4	
rri	d->2	k->130	n->9	s->1	t->21	ä->4	
rro	g->2	n->1	r->11	
rru	m->2	p->7	
rrv	a->1	
rrä	d->1	n->4	t->2	
rrå	d->15	
rró	n->3	
rrö	r->4	s->1	
rs 	1->1	2->1	E->2	a->31	b->20	d->9	e->13	f->25	g->3	h->12	i->23	j->1	k->9	l->7	m->8	n->4	o->12	p->15	r->8	s->19	t->10	u->11	v->3	y->1	ä->3	å->2	ö->5	
rs,	 ->20	
rs-	b->1	
rs.	 ->1	.->1	D->9	H->1	J->3	M->1	N->1	O->1	T->1	U->1	V->4	
rsa	f->1	i->1	k->38	l->1	m->21	n->1	t->5	v->1	
rsb	e->5	r->1	u->1	
rsc	h->1	
rsd	a->8	
rse	 ->7	,->1	.->2	i->1	k->5	l->4	n->34	r->55	s->1	
rsf	r->47	u->4	ö->5	
rsh	i->1	
rsi	e->9	f->2	k->85	n->1	o->13	
rsk	a->43	i->163	j->1	n->35	o->3	r->25	t->1	u->2	ä->4	å->7	
rsl	a->495	i->1	u->1	
rsm	a->1	e->1	i->1	ä->1	å->1	
rso	m->197	n->113	r->1	t->1	
rsp	e->23	o->6	r->20	å->1	
rsr	a->2	
rss	k->2	l->1	
rst	 ->95	.->2	a->277	e->1	i->8	k->1	o->4	r->42	ä->72	å->104	ö->30	
rsu	m->9	n->3	
rsv	a->62	i->15	u->4	ä->7	å->2	
rsy	d->1	n->2	
rsä	k->59	l->5	m->10	n->2	t->35	
rså	g->1	t->1	
rsö	k->109	r->4	v->1	
rt 	-->6	C->1	D->1	E->5	F->1	G->1	a->151	b->24	d->28	e->42	f->72	g->14	h->15	i->37	k->22	l->11	m->37	n->14	o->65	p->35	r->8	s->101	t->20	u->28	v->16	y->2	Ö->1	ä->9	å->1	ö->3	
rt!	H->1	J->1	
rt)	 ->1	
rt,	 ->49	
rt-	 ->1	s->2	
rt.	 ->2	A->1	D->9	E->1	F->2	H->1	I->2	J->7	K->3	L->1	M->2	N->1	O->1	R->1	S->3	U->1	V->7	Ä->1	
rt:	 ->2	
rt?	J->1	
rtN	ä->1	
rta	 ->18	b->1	d->5	g->10	l->8	m->1	n->9	r->5	s->4	t->16	
rtb	e->2	i->1	
rtd	i->1	
rte	c->24	l->15	m->9	n->56	r->109	t->19	x->3	
rtf	a->97	e->1	r->1	ö->1	
rtg	r->4	å->5	
rth	e->1	u->1	y->1	
rti	 ->23	,->7	.->4	d->75	e->42	f->8	g->1	i->1	k->114	l->4	n->2	o->14	p->2	s->8	
rtj	u->1	ä->20	
rtk	o->19	
rtl	e->1	i->7	ä->1	
rtm	a->1	o->1	
rtn	e->28	i->2	ä->1	
rto	g->1	m->23	n->11	
rtp	l->1	r->2	
rtr	a->5	e->1	o->60	y->2	ä->10	ö->1	
rts	 ->52	,->6	.->6	a->13	e->6	i->6	k->1	m->2	o->2	s->3	ä->89	
rtu	g->97	n->2	s->3	t->2	
rtv	i->2	
rty	d->3	g->107	r->1	
rtz	 ->2	,->1	
rtä	c->1	n->2	
ru 	A->3	B->1	F->1	L->1	M->1	P->2	R->3	S->4	T->1	W->1	k->46	l->2	t->83	
ru,	 ->1	
rua	r->16	
rub	b->3	r->2	
ruc	k->2	
rue	r->5	
ruh	e->2	
rui	n->1	
ruk	 ->9	!->1	,->9	a->17	e->20	i->1	n->1	s->23	t->202	
rul	l->6	
rum	 ->40	!->1	,->5	.->4	e->55	p->2	
run	a->1	d->307	g->19	k->3	o->1	t->10	
rup	p->231	t->7	
rus	a->5	t->15	
rut	 ->2	.->1	a->2	b->3	e->5	g->1	i->10	o->15	s->64	t->4	v->4	ö->1	
ruv	a->1	i->15	
rv 	f->1	o->2	
rv,	 ->3	
rv.	"->1	B->1	E->1	
rva	 ->6	d->1	k->25	l->54	n->6	r->49	t->29	
rvb	r->1	
rve	c->1	n->13	r->28	t->5	
rvh	e->1	
rvi	c->7	d->9	n->74	r->12	s->11	
rvj	u->3	
rvl	i->2	
rvr	i->1	ä->1	
rvs	a->3	i->1	s->2	
rvt	 ->2	r->1	
rvu	n->3	
rvä	g->49	l->3	n->32	r->19	
rvå	n->6	
rwe	l->1	
ry 	F->1	o->1	
ry,	 ->1	
ry.	D->1	
ryc	k->105	
ryf	t->1	
ryg	g->16	t->3	
ryk	.->1	a->29	e->2	s->2	t->9	
rym	d->2	m->12	s->1	t->1	
ryo	s->1	
ryp	h->3	s->1	t->2	
ryr	 ->2	
rys	 ->1	a->2	k->2	n->1	s->21	
ryt	a->8	e->9	n->2	t->2	
rzw	a->1	
rä 	u->1	ö->1	
räc	k->153	
räd	 ->5	,->1	.->1	a->78	d->31	e->66	s->11	
räf	f->117	t->30	
räg	a->1	e->36	l->6	
räk	e->9	n->55	t->2	
räl	 ->2	,->1	
räm	b->1	d->1	e->1	j->62	l->35	m->5	s->48	
rän	 ->6	a->3	d->79	g->69	i->13	k->31	n->5	s->141	t->1	
räp	n->1	r->1	
rär	 ->1	t->1	
räs	c->2	k->1	
rät	a->1	o->1	t->754	
räv	a->68	d->4	e->45	i->1	s->55	t->2	
rå 	s->1	v->1	ä->1	
råd	 ->17	,->4	.->5	?->1	a->16	d->1	e->651	f->6	g->27	s->48	
råe	r->1	t->1	
råg	a->563	e->13	n->8	o->275	
råk	 ->5	.->1	a->10	e->4	i->3	l->3	o->2	r->30	t->1	
rål	d->3	k->1	n->3	s->1	
rån	 ->601	,->3	.->2	g->7	k->3	t->3	v->9	
råo	l->1	
råp	s->1	
rår	i->12	
rås	 ->2	
råt	 ->1	g->1	t->1	
råz	o->1	
réb	e->1	
réf	é->1	
rêt	s->1	
rín	c->1	
rón	 ->5	
röd	.->3	a->5	e->3	g->1	o->1	
rög	h->1	
röj	a->8	d->1	e->3	o->1	s->2	t->1	
rök	 ->1	,->1	s->1	
röm	 ->4	,->1	:->1	m->8	n->6	t->1	v->1	
rön	 ->2	a->16	b->1	i->1	t->1	
rör	 ->50	a->29	d->24	e->9	i->2	l->24	s->8	t->5	
rös	 ->3	a->3	k->3	t->183	
röt	 ->5	s->2	t->8	
röv	a->14	e->1	n->5	o->1	r->2	s->1	
s "	B->1	g->1	
s (	P->1	f->1	u->1	
s -	 ->20	,->1	
s 1	9->5	
s 2	 ->1	0->2	4->1	8->1	
s 3	,->1	
s 4	0->1	
s 8	0->1	
s A	d->1	l->1	
s B	N->3	a->3	l->1	
s C	E->1	
s D	a->1	e->3	
s E	G->2	U->2	u->13	
s F	P->1	
s G	e->1	i->1	o->1	
s H	e->1	
s I	s->1	
s L	e->1	
s M	i->1	
s O	z->1	
s P	a->1	
s R	E->1	u->1	
s S	O->1	j->2	p->3	
s V	D->1	i->1	
s W	i->1	u->1	
s X	X->1	
s a	b->3	d->1	g->3	k->1	l->48	m->3	n->99	r->41	t->174	u->4	v->288	x->1	
s b	a->8	e->143	i->9	l->15	o->8	r->9	u->15	y->4	ä->7	å->4	ö->1	
s c	e->7	i->1	o->1	
s d	a->22	e->204	i->26	j->1	o->13	r->2	u->2	ä->31	å->3	ö->5	
s e	f->24	g->18	k->30	l->23	m->8	n->124	r->3	t->43	u->3	v->1	x->12	
s f	a->25	e->4	i->11	j->1	l->16	o->27	r->113	u->21	y->4	å->10	ö->302	
s g	a->6	e->65	i->5	j->1	o->8	r->31	u->1	ä->3	å->4	ö->4	
s h	a->59	e->6	i->12	j->5	o->6	u->7	y->1	ä->34	å->7	ö->3	
s i	 ->299	d->4	g->4	h->1	k->2	l->2	m->1	n->225	r->1	
s j	a->11	o->2	u->20	ä->1	
s k	a->18	e->1	l->13	o->93	r->13	u->14	v->12	ä->5	ö->1	
s l	a->25	e->27	i->28	j->1	o->6	u->2	ä->12	å->1	ö->3	
s m	a->15	e->200	i->24	o->21	y->17	ä->6	å->41	ö->19	
s n	a->24	e->9	i->7	o->2	u->16	y->12	ä->22	å->33	ö->3	
s o	a->3	b->6	c->228	d->2	e->1	f->10	h->2	i->5	k->1	l->10	m->93	r->57	s->5	t->5	v->1	
s p	a->25	e->10	h->1	l->6	o->34	r->41	u->2	å->163	
s q	u->2	
s r	a->24	e->83	i->13	o->13	u->4	y->2	ä->51	å->4	ö->6	
s s	a->46	c->1	e->18	i->40	j->15	k->65	l->19	m->2	n->6	o->122	p->11	t->90	u->8	v->10	y->10	ä->26	å->24	ö->2	
s t	a->15	e->13	i->157	j->13	o->3	r->19	u->4	v->12	y->10	
s u	n->44	p->71	r->8	t->117	
s v	a->45	e->32	i->72	o->2	u->1	ä->41	å->4	
s y	r->2	t->19	
s ä	g->7	n->21	r->50	v->7	
s å	l->5	r->8	s->11	t->38	
s ö	d->5	g->2	k->5	m->2	n->2	p->2	r->3	v->38	
s! 	J->1	V->1	
s!D	e->1	
s!E	u->1	
s!F	ö->1	
s!G	e->1	
s!H	e->1	
s!V	i->1	
s".	D->1	J->1	K->1	
s) 	f->1	o->1	
s, 	1->1	E->1	L->1	M->1	S->1	T->1	W->1	a->18	b->6	d->16	e->20	f->23	g->4	h->8	i->14	j->4	k->7	l->1	m->32	n->9	o->52	p->7	r->1	s->32	t->6	u->11	v->15	ä->6	å->4	
s- 	f->1	o->42	
s-,	 ->1	
s-C	a->1	
s-J	ø->2	
s-b	e->2	i->1	
s-d	e->1	
s-f	ö->1	
s-i	n->2	
s-n	o->1	y->1	
s-p	r->1	
s-s	i->1	
s. 	1->2	D->3	E->2	M->2	P->1	W->1	a->11	d->4	e->3	f->3	g->1	h->2	i->5	j->1	m->4	n->1	o->2	p->1	s->1	v->2	
s.(	E->1	
s.)	Å->1	
s.-	 ->1	
s..	(->1	
s.A	l->3	n->2	t->1	
s.B	e->4	l->2	
s.C	e->1	
s.D	a->1	e->83	i->1	ä->12	å->4	
s.E	f->2	k->1	n->8	r->1	t->5	u->3	
s.F	a->1	l->2	r->7	ö->8	
s.G	e->4	r->1	
s.H	a->1	e->11	i->2	o->1	u->2	ä->1	
s.I	 ->12	n->3	
s.J	a->28	o->1	u->1	ä->1	
s.K	o->8	
s.L	a->1	e->1	å->2	
s.M	a->3	e->13	i->2	y->1	ä->1	å->1	
s.N	i->1	u->2	ä->4	å->1	
s.O	L->1	a->1	m->2	n->1	
s.P	a->3	e->1	r->2	å->2	
s.R	a->1	e->4	å->1	
s.S	a->3	e->1	l->5	n->1	o->2	å->1	
s.T	a->3	i->1	y->1	
s.U	n->4	t->2	
s.V	a->6	i->31	å->3	
s.Y	t->2	
s.k	.->4	
s.Ä	n->3	v->2	
s.Å	t->2	
s/d	e->1	
s/i	n->1	
s: 	a->2	e->1	f->1	h->1	k->1	v->1	
s; 	a->1	b->1	d->1	e->1	o->1	v->1	
s?.	 ->1	H->1	
s?D	e->1	
s?E	t->1	
s?F	r->1	
s?H	a->1	
s?I	 ->1	
s?J	a->1	o->1	
s?K	o->1	
s?O	c->1	
s?S	k->1	
s?T	i->1	
s?V	i->2	
s?Ä	r->1	
sNä	s->1	
sa 	(->1	-->1	1->1	2->3	3->1	P->1	R->1	a->56	b->29	c->1	d->28	e->9	f->66	g->15	h->18	i->31	k->32	l->19	m->48	n->5	o->47	p->61	r->33	s->65	t->34	u->22	v->25	ä->36	å->9	ö->3	
sa!	L->1	
sa,	 ->22	
sa.	.->1	A->1	B->2	D->6	E->1	F->2	H->1	I->2	J->3	K->1	M->4	R->1	S->1	U->1	Å->1	
sa?	P->1	
sab	e->3	l->1	o->8	
sac	a->1	e->3	
sad	 ->18	,->2	.->3	e->108	ö->1	
saf	e->1	f->2	t->1	
sag	 ->1	e->1	t->49	
sai	l->1	
sak	 ->39	,->2	.->5	:->1	a->20	e->60	f->1	k->2	l->11	n->39	o->2	p->1	r->1	t->9	
sal	a->1	e->2	i->1	m->1	t->1	u->1	
sam	 ->70	,->2	.->1	a->83	b->47	e->2	f->13	h->144	k->3	l->46	m->493	o->37	r->10	s->7	t->204	v->5	
san	 ->7	,->2	.->3	a->6	d->20	f->1	k->8	l->9	m->1	n->17	s->6	t->36	
sar	 ->87	!->1	,->4	.->2	b->27	e->5	g->1	n->1	t->3	
sas	 ->31	,->1	.->1	p->3	
sat	 ->42	,->1	.->5	e->1	i->46	o->3	s->141	t->65	
sau	r->1	
sav	b->1	g->8	i->1	t->15	v->1	
sba	n->2	r->5	s->2	
sbe	d->4	f->9	g->4	h->4	k->3	l->7	r->2	s->33	t->5	v->7	
sbi	d->2	l->7	s->2	
sbo	l->3	r->3	u->5	
sbr	i->2	o->2	u->16	
sbu	d->3	r->1	s->1	t->1	
sby	g->44	
sbå	d->1	
sbö	r->12	
sca	y->6	
sce	n->15	r->1	
sch	 ->4	!->1	.->1	?->1	a->1	e->23	h->1	l->4	w->1	
sci	e->1	p->14	s->12	
sco	r->1	
scy	k->3	
sda	g->15	
sde	b->3	l->14	p->1	
sdi	g->2	k->5	m->1	r->7	
sdo	k->6	m->4	
sdr	a->4	ä->1	
sdu	g->5	k->1	
sdö	m->2	
se 	(->1	-->3	G->1	a->54	b->2	d->17	e->7	f->33	g->3	h->10	i->11	j->3	k->7	l->1	m->22	n->5	o->29	p->12	r->3	s->28	t->71	u->6	v->15	ä->4	ö->14	
se"	,->1	
se,	 ->19	
se-	 ->1	N->1	
se.	B->1	D->6	E->4	F->1	J->3	K->1	L->1	M->4	N->1	O->1	S->2	V->3	
se;	 ->1	
se?	E->1	
sea	k->1	
seb	a->1	y->1	
sed	 ->1	a->104	d->5	e->1	
see	n->60	
sef	f->7	u->11	
seg	 ->1	d->1	e->4	l->13	r->3	
seh	i->1	
sei	l->1	s->2	
sek	e->4	l->2	o->26	r->16	t->91	u->3	v->61	
sel	 ->15	!->2	,->5	-->3	.->3	b->1	e->3	f->1	l->3	o->1	s->103	ö->3	
sem	e->7	i->4	ö->1	
sen	 ->285	!->1	,->44	.->84	;->1	?->2	N->2	a->116	b->3	d->9	f->1	h->4	i->13	l->3	r->1	s->31	t->91	
seo	m->1	
sep	a->1	t->15	
ser	 ->544	!->1	,->40	.->43	:->1	?->3	a->163	b->15	i->102	l->13	n->140	s->1	v->23	
ses	 ->22	.->1	i->5	s->6	
set	 ->32	,->1	.->3	a->1	i->1	s->1	t->69	ê->2	
seu	r->1	t->1	
sev	i->2	ä->14	
sew	i->1	
sex	 ->17	,->1	i->1	m->1	p->1	t->1	u->3	v->1	
sfa	k->1	l->6	r->2	s->6	t->11	
sfe	l->2	
sfi	e->31	n->1	s->3	
sfl	a->15	o->2	y->1	
sfo	n->22	r->8	s->1	
sfr	i->60	ä->4	å->45	
sfu	l->16	n->2	
sfä	r->1	s->1	
sfå	n->1	
sfö	r->292	
sga	r->3	s->4	
sge	m->1	
sgi	l->1	v->16	
sgr	a->5	e->2	u->11	ä->3	
sgy	n->7	
sgå	 ->2	s->1	
sgö	r->1	
sh 	P->2	
sh,	 ->1	
sha	l->1	n->15	t->1	u->1	v->1	
she	m->1	r->1	t->51	
shi	n->14	p->1	
shj	ä->2	
sho	p->1	t->1	
shu	s->2	
shä	m->2	n->1	
shå	l->1	
sia	s->3	t->2	
sib	i->1	
sid	a->78	e->11	i->35	k->1	o->7	u->1	
sie	l->37	n->7	r->50	
sif	f->22	i->14	u->1	
sig	 ->369	,->8	.->18	;->1	a->16	n->16	t->14	
sik	 ->2	e->3	t->219	
sil	 ->1	a->2	i->1	v->3	
sim	i->2	m->1	u->2	
sin	 ->169	.->1	a->138	d->8	e->3	f->3	g->20	i->9	n->8	o->1	r->4	s->22	t->4	
sio	n->1299	
sis	 ->4	,->1	k->98	m->15	t->77	
sit	e->1	i->90	l->3	r->1	t->107	u->126	
siv	 ->8	.->1	a->8	e->17	t->11	
siä	r->2	
sjo	v->17	
sju	 ->5	,->1	k->13	n->13	r->2	t->2	
sjä	l->173	t->19	
sjö	f->8	m->2	n->5	s->4	t->1	v->1	
sk 	-->1	T->1	a->20	b->21	c->2	d->15	e->3	f->19	g->8	h->8	i->13	j->5	k->37	l->17	m->15	n->19	o->27	p->28	r->20	s->30	t->10	u->23	v->4	ä->1	å->13	ö->3	
sk,	 ->7	
sk-	b->1	f->1	i->1	s->1	
sk.	 ->1	D->1	H->4	I->3	J->1	M->1	O->1	V->1	
ska	 ->1579	,->18	.->12	:->2	b->1	d->82	f->26	k->2	l->679	m->10	n->54	p->667	r->49	s->17	t->80	
skb	e->8	
ske	 ->96	!->1	)->2	,->6	.->2	d->15	k->1	l->3	m->7	n->18	o->2	p->17	r->79	s->1	t->23	v->2	
skf	a->1	r->1	y->1	ö->1	
skh	a->6	e->1	
ski	c->17	e->2	f->6	l->259	n->10	p->12	s->8	
skj	u->31	
skk	a->1	o->2	
skl	a->25	i->45	
skn	i->78	
sko	a->2	e->1	f->2	g->38	h->3	l->13	m->46	n->170	p->3	r->84	s->11	t->166	u->1	v->2	
skr	a->61	e->9	i->140	o->42	ä->27	
skt	 ->256	!->1	,->7	.->12	a->1	
sku	g->3	l->508	n->1	p->1	r->8	s->62	t->84	
skv	a->8	o->3	ä->13	
sky	 ->1	d->108	f->1	h->1	l->34	m->1	n->15	v->1	
skä	l->52	m->4	n->5	r->17	
skå	d->10	l->1	r->1	
skö	n->1	p->1	r->7	t->23	v->1	
sla	 ->18	"->1	,->2	.->1	d->1	g->623	k->1	m->1	n->21	p->3	r->5	t->1	v->2	
sle	d->39	n->2	r->1	s->5	
sli	b->1	e->1	g->158	n->5	p->2	r->1	s->48	t->1	v->14	
slo	 ->1	,->2	b->1	g->20	l->1	m->1	p->2	r->5	t->1	v->1	
slu	k->3	m->5	n->1	s->2	t->521	
sly	c->18	
slä	c->3	g->9	k->4	m->2	n->35	p->21	
slå	 ->33	d->1	e->1	n->1	r->47	s->27	
slö	j->6	s->58	t->3	
sm 	-->1	e->3	f->1	h->1	i->1	m->1	o->18	p->2	s->6	u->1	ä->2	ö->1	
sm,	 ->11	
sm.	D->7	F->1	H->1	I->2	J->1	M->1	N->1	O->2	V->4	
sm?	V->1	
sma	j->1	k->5	n->16	r->15	s->2	t->1	
sme	d->116	k->2	n->22	r->9	t->6	
smi	d->3	l->5	n->16	s->2	t->3	
smo	d->2	l->1	m->5	n->1	t->1	
smu	g->1	l->1	s->1	t->3	
smy	n->31	
smä	d->1	l->1	n->33	r->4	s->12	
små	 ->53	,->2	.->1	f->5	g->1	l->12	n->4	s->1	
smö	j->4	n->1	t->2	
sna	 ->13	,->2	b->71	c->2	d->4	r->72	t->9	
sne	d->13	
sni	e->2	n->108	t->15	v->33	
sno	r->7	
sny	c->1	h->1	
snä	l->1	t->3	v->1	
snå	l->5	r->1	
snö	j->3	v->1	
so 	e->1	f->1	i->1	o->1	ä->2	
so,	 ->1	
so-	 ->1	
soc	h->1	i->207	
sod	l->1	
soe	f->1	
sof	f->2	i->5	t->1	
sol	a->1	d->2	e->7	i->33	l->1	s->1	u->140	y->1	
som	 ->3643	,->22	g->1	l->3	m->3	r->41	s->1	
son	 ->13	,->1	.->1	a->25	e->46	g->1	i->5	l->34	s->1	t->3	
sop	a->1	
sor	 ->8	,->4	.->2	b->1	d->36	e->1	g->24	i->4	n->1	t->8	
sos	 ->2	,->1	k->1	ä->2	
sot	 ->1	
sov	j->1	o->60	å->3	
sp"	,->1	
sp.	 ->2	
spa	k->8	n->12	r->21	t->2	
spe	c->85	g->12	k->152	l->56	n->13	r->19	t->2	
spi	c->1	l->1	n->1	r->3	s->1	
spl	a->43	i->11	
spo	,->1	l->128	n->7	r->110	s->5	t->1	
spr	a->1	i->103	o->105	u->19	å->26	
spu	n->18	
spä	n->11	r->3	
spå	f->1	r->13	
spö	k->4	
squ	e->1	i->1	
sra	d->1	e->58	m->8	p->6	
sre	a->1	d->2	f->2	g->39	k->5	l->1	p->6	s->10	
sri	k->17	l->1	s->3	
sro	l->1	
sru	b->1	h->2	m->1	n->2	t->1	
sry	c->1	m->2	
srä	d->1	t->61	
srå	d->23	
srö	r->2	
ss 	-->1	a->49	b->11	d->24	e->24	f->34	g->9	h->9	i->42	k->10	l->6	m->30	n->11	o->45	p->22	r->11	s->55	t->25	u->13	v->19	y->1	ä->13	å->16	ö->6	
ss"	.->1	
ss)	 ->1	
ss,	 ->24	
ss.	A->1	D->8	E->3	F->2	H->2	J->4	M->2	N->2	S->1	V->7	Ä->2	
ss:	 ->1	
ss?	.->1	J->1	V->1	
ssa	 ->516	!->1	,->4	.->8	b->8	d->9	g->2	k->1	l->1	m->14	n->25	r->9	s->7	t->1	v->1	
ssb	e->5	r->10	
ssc	h->1	
sse	 ->21	,->5	-->1	.->3	?->1	d->1	k->19	l->128	n->125	r->49	t->7	
ssf	a->1	o->2	ö->4	
ssg	y->7	
ssh	e->4	u->1	ä->1	
ssi	d->1	f->12	g->32	l->3	m->2	n->1	o->1223	s->7	t->4	v->12	
ssj	ö->1	
ssk	a->6	e->3	i->11	o->2	r->8	y->5	ä->3	ö->6	
ssl	a->14	y->18	ö->2	
ssm	e->4	
ssn	a->28	i->7	ö->3	
sso	 ->5	,->1	c->1	n->1	r->9	
ssp	e->1	r->2	
ssr	e->3	ä->2	
sst	 ->8	a->316	e->5	i->1	o->1	r->25	y->7	ä->49	å->1	ê->1	ö->31	
ssu	e->1	p->2	s->1	t->61	
ssv	ä->4	å->1	
ssy	n->2	s->57	
ssä	k->66	l->7	n->1	t->10	
st 	-->3	1->3	2->1	3->2	4->1	5->1	7->1	9->1	D->1	E->3	I->1	M->1	P->1	a->47	b->13	c->1	d->40	e->23	f->46	g->16	h->24	i->43	j->2	k->25	l->14	m->34	n->28	o->51	p->45	r->14	s->52	t->31	u->17	v->48	ä->11	å->5	ö->4	
st!	D->1	T->1	
st,	 ->26	
st-	 ->1	b->5	
st.	 ->1	A->1	D->3	E->1	F->2	G->1	J->3	K->2	M->2	N->2	V->4	Ä->1	
st:	 ->1	
st?	N->1	V->1	
sta	 ->513	,->16	.->14	:->5	;->2	?->1	N->1	a->1	b->25	c->1	d->96	g->62	i->22	k->7	l->6	m->1	n->183	r->105	s->8	t->624	u->1	v->2	
stb	a->4	e->2	i->1	l->1	r->1	
std	e->11	
ste	 ->850	,->4	.->3	:->1	d->4	e->6	f->7	g->67	i->1	k->2	l->9	m->229	n->72	p->1	r->505	s->5	t->4	u->9	x->3	
stf	l->1	u->1	ä->8	ö->8	
stg	r->3	ö->3	
sth	a->1	o->3	ä->1	å->1	
sti	a->1	c->9	d->14	e->1	f->128	g->19	k->6	l->61	m->11	n->28	o->1	p->1	s->93	t->165	
stj	ä->9	
stk	l->1	o->1	u->2	ä->1	
stl	a->3	i->3	ä->3	
stm	a->2	y->3	ä->2	
stn	a->109	i->72	ä->2	
sto	 ->2	d->16	l->103	m->2	n->27	p->20	r->380	w->3	
stp	a->5	
str	a->164	e->28	i->172	o->97	u->247	y->35	ä->131	å->6	ö->23	
sts	 ->2	.->2	a->2	e->2	l->21	t->51	v->1	
stt	o->1	y->2	
stu	 ->1	d->14	g->1	l->1	m->1	n->17	r->2	t->2	
stv	a->1	e->1	i->4	ä->1	
sty	c->5	m->3	r->53	
stä	d->21	l->426	m->226	n->126	r->51	t->1	v->2	
stå	 ->65	,->3	.->2	:->1	d->2	e->46	l->41	n->226	r->183	s->6	t->30	
stê	t->1	
stö	d->427	l->1	r->137	t->19	
sua	l->1	
sub	j->1	s->27	v->10	
suc	c->5	
sud	d->1	
sue	l->2	
sug	a->1	
sul	 ->2	.->1	e->3	t->121	
sum	 ->1	b->1	e->61	m->20	t->2	
sun	d->11	e->1	
sup	p->6	r->1	
sur	d->1	s->50	t->2	
sus	 ->3	e->1	p->1	
sut	a->3	b->15	o->61	r->5	s->6	t->2	v->3	ö->1	
suv	e->17	
sv.	 ->3	,->1	?->1	S->1	
sva	g->44	l->1	n->2	r->466	t->2	
sve	k->2	n->3	p->3	r->7	
svi	k->8	l->22	n->16	s->32	
svu	n->4	
svä	g->1	l->2	m->7	n->2	r->29	s->6	t->1	v->1	
svå	g->2	n->1	r->95	
swa	g->1	
syd	d->1	e->1	k->1	v->1	ö->1	
syf	t->74	
syk	o->1	
syl	 ->4	,->2	-->1	.->3	b->1	f->2	r->2	s->6	
sym	b->9	p->9	
syn	 ->83	,->2	.->4	;->1	a->4	d->8	e->9	l->8	n->52	o->1	p->29	s->7	t->4	v->12	
syr	a->3	i->8	
sys	 ->1	s->109	t->191	
säg	:->1	a->180	e->81	n->2	s->5	
säk	e->321	r->64	t->15	
säl	j->8	l->12	
säm	n->2	r->15	s->5	
sän	d->22	k->8	
sär	 ->3	a->1	b->1	e->4	k->1	s->156	
säs	o->1	
sät	e->1	t->682	
så 	"->1	-->2	1->1	E->4	F->1	M->1	a->211	b->43	d->35	e->41	f->66	g->23	h->41	i->55	j->2	k->61	l->34	m->92	n->18	o->17	p->23	r->12	s->153	t->42	u->23	v->69	z->1	ä->36	å->3	ö->4	
så,	 ->18	
så.	 ->1	D->2	I->2	J->1	N->1	O->1	P->1	
så:	 ->1	
såd	a->163	
såg	 ->18	s->4	v->1	
såh	ä->1	
sål	d->2	e->40	u->4	
sån	g->3	
sår	b->3	e->1	
sås	o->32	
såt	e->2	g->12	i->1	
såv	i->3	ä->40	
sí 	ä->1	
söd	a->1	e->1	r->6	
sök	 ->11	,->2	a->60	e->26	n->24	t->20	
sön	d->7	e->1	
sör	j->16	
söv	e->15	n->1	
t "	E->1	K->4	O->1	P->1	e->4	k->1	o->1	r->2	
t (	5->1	8->2	9->1	B->2	C->1	E->2	F->1	I->2	S->1	a->1	d->1	f->2	h->1	i->2	k->1	t->2	Ö->1	
t ,	 ->1	
t -	 ->89	,->2	e->1	
t 1	 ->2	,->1	0->2	1->1	2->1	3->1	8->1	9->19	
t 2	 ->2	0->1	1->1	2->1	3->1	5->2	6->1	7->1	
t 3	 ->2	9->1	
t 4	 ->2	0->3	8->1	
t 5	 ->1	,->2	0->1	
t 6	 ->1	
t 7	 ->1	0->3	
t 8	 ->1	0->1	8->2	
t 9	 ->1	0->1	3->1	4->1	5->1	8->1	
t :	 ->1	
t A	B->1	d->1	i->1	k->1	l->4	m->3	s->1	u->1	
t B	N->1	a->3	e->2	o->1	r->3	
t C	E->1	a->2	l->1	
t D	 ->1	a->6	e->1	u->2	
t E	G->12	I->1	K->1	L->1	U->22	l->1	q->8	r->3	u->111	v->1	
t F	E->1	N->2	P->3	l->4	r->3	ö->5	
t G	a->1	o->1	r->5	
t H	a->4	e->1	
t I	 ->1	C->1	N->1	n->2	r->1	s->4	t->3	
t J	o->3	ö->3	
t K	a->1	i->1	o->4	u->3	y->2	
t L	a->1	e->2	
t M	a->2	i->2	o->4	ü->1	
t N	a->1	
t O	L->3	
t P	a->1	e->1	o->6	
t R	I->2	a->5	o->1	
t S	E->1	a->2	c->1	j->2	o->2	t->3	u->1	v->1	
t T	V->1	h->3	i->1	o->3	u->14	
t U	N->1	
t V	a->1	e->1	o->1	ä->1	
t W	a->2	u->1	
t a	b->8	c->12	d->7	g->16	i->1	k->18	l->119	m->6	n->331	r->123	s->3	t->816	v->599	
t b	a->49	e->439	i->69	l->86	o->23	r->76	u->11	y->21	ä->30	å->8	ö->60	
t c	a->1	e->7	h->2	i->8	
t d	)->1	a->27	e->1341	i->83	j->7	o->27	r->43	u->2	y->6	ä->44	å->18	ö->13	
t e	)->1	-->1	d->1	f->62	g->35	k->24	l->43	m->9	n->341	p->1	r->53	t->123	u->48	v->5	x->58	
t f	.->1	a->164	e->27	i->229	j->4	l->34	o->69	r->298	u->37	y->4	ä->3	å->134	ö->1241	
t g	a->32	e->211	i->8	j->7	l->20	o->95	r->49	y->6	ä->224	å->48	ö->141	
t h	a->414	e->39	i->25	j->20	o->38	u->31	y->3	ä->103	å->41	ö->52	
t i	 ->500	.->1	a->1	b->6	c->4	d->9	f->15	g->10	l->4	m->6	n->630	r->8	s->4	t->4	
t j	a->109	o->6	u->28	ä->9	
t k	a->125	e->1	l->56	n->7	o->492	r->93	u->87	v->21	y->1	ä->26	ö->7	
t l	a->80	e->40	i->65	j->2	o->13	u->7	y->23	ä->122	å->29	ö->32	
t m	a->259	e->450	i->197	o->90	u->6	y->102	ä->18	å->155	ö->57	
t n	a->22	e->19	i->58	o->30	r->1	u->52	y->63	ä->88	å->70	ö->35	
t o	a->13	b->9	c->724	d->1	e->5	f->27	g->2	k->4	l->17	m->322	n->6	p->8	r->60	s->55	t->8	v->2	ä->1	ö->2	
t p	a->108	e->43	i->1	l->24	o->135	r->143	u->5	å->326	
t r	a->18	e->172	i->50	o->2	u->13	y->4	ä->67	å->53	ö->58	
t s	.->1	a->154	e->148	i->118	j->30	k->392	l->46	m->4	n->21	o->543	p->45	t->436	u->9	v->56	y->72	ä->283	å->130	ö->7	
t t	.->1	a->192	e->14	h->1	i->407	j->5	o->17	r->62	u->6	v->27	y->44	ä->23	å->3	
t u	l->1	n->140	p->181	r->26	t->319	
t v	a->228	e->70	i->828	o->13	r->1	ä->102	å->48	
t w	o->1	
t y	p->1	t->34	
t z	o->1	
t Ö	s->6	
t ä	c->1	g->24	m->8	n->97	r->885	v->39	
t å	 ->3	k->1	l->7	r->35	s->7	t->89	v->1	
t ö	d->3	g->5	k->30	l->1	m->1	n->8	p->13	s->15	v->113	
t! 	D->2	J->2	N->1	S->1	V->1	
t!"	J->1	
t!(	P->1	
t!.	 ->1	(->1	
t!D	e->1	ä->1	
t!H	e->3	
t!J	a->1	
t!K	u->1	
t!L	e->1	
t!M	e->1	
t!N	ä->1	
t!P	r->1	
t!T	v->1	
t" 	(->1	g->1	m->1	o->1	ä->1	
t",	 ->4	
t".	E->1	J->1	
t) 	(->1	C->1	h->2	p->1	s->1	t->1	
t),	 ->3	
t).	D->1	H->2	L->1	
t)N	ä->1	
t, 	"->1	C->1	D->1	E->2	G->1	H->1	I->3	J->1	L->1	O->1	P->1	S->2	W->1	Z->1	a->43	b->20	c->1	d->61	e->59	f->67	g->15	h->50	i->50	j->9	k->36	l->11	m->89	n->21	o->137	p->16	r->11	s->140	t->24	u->39	v->63	ä->33	å->4	ö->2	
t- 	o->3	
t-E	x->1	
t-a	n->5	
t-b	e->5	
t-f	r->1	
t-s	t->2	
t. 	(->1	7->2	A->1	D->18	E->1	F->1	H->2	I->3	J->1	K->1	M->1	O->1	S->1	V->3	a->1	
t.(	A->1	F->1	P->3	
t.)	A->1	B->2	F->1	R->1	
t.-	 ->1	
t..	 ->2	(->1	.->2	H->1	
t.1	9->1	
t.A	c->1	l->5	n->2	r->2	t->2	v->9	
t.B	e->5	i->1	l->1	o->1	r->1	å->2	
t.D	a->1	e->242	i->3	ä->17	å->5	
t.E	G->1	f->7	k->1	n->18	r->1	t->6	u->10	
t.F	P->1	e->1	i->1	l->2	r->22	ö->41	
t.G	e->4	i->1	r->2	
t.H	a->5	e->49	i->1	u->5	ä->7	
t.I	 ->44	b->1	n->5	
t.J	a->147	u->2	
t.K	o->18	r->1	u->2	ä->2	
t.L	a->1	i->2	ä->1	å->11	
t.M	a->16	e->52	i->13	o->4	å->1	
t.N	a->5	i->7	u->8	ä->11	å->1	ö->1	
t.O	K->1	b->1	c->12	f->1	m->16	r->3	
t.P	P->1	a->8	l->1	o->1	r->4	u->1	å->7	
t.R	a->1	e->3	i->1	ä->1	
t.S	a->3	e->1	k->3	l->6	o->6	t->8	y->1	å->10	
t.T	a->7	h->1	i->4	r->3	u->1	v->1	y->3	
t.U	n->5	r->1	t->3	
t.V	a->23	i->90	ä->1	å->3	
t.e	x->20	
t.o	.->7	
t.Ä	n->3	r->1	v->7	
t.Å	 ->3	r->2	t->1	
t.Ö	k->1	s->1	v->1	
t: 	"->4	E->1	F->1	H->1	J->2	U->2	V->1	a->1	d->5	e->2	f->2	h->1	j->2	k->1	m->1	o->2	s->1	t->1	u->1	v->2	ö->1	
t; 	D->1	a->2	d->5	e->1	f->2	u->1	å->1	
t? 	M->1	R->1	
t?.	 ->2	(->2	
t?A	n->1	t->1	v->1	
t?D	e->4	
t?E	t->1	u->1	
t?H	e->1	u->2	
t?I	 ->1	
t?J	a->4	o->1	
t?K	o->1	ä->1	
t?N	e->3	i->2	ä->1	
t?O	c->1	m->1	
t?R	I->1	
t?S	k->2	
t?T	ä->1	
t?U	t->1	
t?V	a->1	i->4	
t?Ä	r->1	
tBe	t->1	
tJa	g->1	
tNä	s->1	
ta 	-->8	1->1	A->2	E->10	F->1	J->1	M->1	N->1	S->2	a->117	b->131	c->3	d->174	e->123	f->242	g->63	h->116	i->129	j->2	k->75	l->29	m->172	n->39	o->149	p->186	r->68	s->287	t->68	u->116	v->71	y->2	Ö->2	ä->194	å->24	ö->16	
ta!	D->1	F->1	
ta,	 ->82	
ta.	 ->3	(->1	)->1	-->1	.->2	A->1	B->2	C->1	D->28	E->6	F->3	G->1	H->4	I->7	J->12	K->1	M->7	N->2	O->4	P->3	S->7	T->2	V->16	Ä->1	
ta:	 ->6	
ta;	 ->2	
ta?	D->1	J->1	N->1	V->1	
taN	ä->1	
taa	f->1	
tab	 ->1	a->1	e->38	i->24	l->26	r->3	u->2	
tac	k->149	
tad	 ->17	,->2	.->25	e->86	g->29	i->8	k->24	m->2	s->4	t->1	
taf	r->10	
tag	 ->73	,->20	.->21	?->1	a->172	b->15	e->91	i->100	l->5	n->23	s->35	
tai	n->26	
tak	 ->1	,->2	a->5	e->3	l->1	t->26	u->1	
tal	 ->122	"->1	,->6	-->3	.->11	:->1	F->1	a->375	b->2	e->80	f->5	i->45	j->35	l->14	m->418	n->15	o->2	r->4	s->37	t->9	v->1	y->2	
tam	e->9	i->2	p->1	
tan	 ->372	,->10	.->17	;->1	?->1	a->1	b->1	d->183	e->8	f->32	k->101	n->24	o->1	s->71	t->18	v->1	
tap	o->1	p->8	
tar	 ->349	,->6	.->9	b->32	e->69	h->1	i->39	k->62	l->2	m->10	n->19	t->16	v->1	
tas	 ->176	,->10	.->15	i->3	k->1	p->2	t->101	ä->1	
tat	 ->172	,->16	.->30	:->2	?->2	e->414	i->58	l->101	o->1	s->79	t->8	u->13	ö->6	ü->1	
tau	e->1	n->3	r->1	
tav	 ->2	l->8	
tax	-->3	e->1	
tba	l->2	n->4	r->3	s->2	
tbe	f->2	h->1	s->4	t->7	v->1	
tbi	l->65	
tbl	o->1	
tbo	k->53	l->1	
tbr	a->1	e->4	i->1	
tbu	d->4	r->1	
tby	g->3	t->17	
tc.	 ->3	D->1	E->1	
tc?	A->1	
tch	a->1	e->1	
tde	l->3	m->11	r->1	
tdi	k->1	r->1	
te 	(->2	-->9	1->1	B->1	E->12	F->2	I->1	J->1	O->1	Q->1	a->197	b->195	c->5	d->128	e->80	f->193	g->116	h->189	i->101	j->14	k->146	l->79	m->142	n->66	o->87	p->81	r->75	s->223	t->128	u->92	v->170	ä->101	å->29	ö->22	
te!	D->1	M->1	
te,	 ->38	
te-	 ->1	L->1	
te.	 ->1	.->1	A->2	B->1	D->10	F->3	H->3	I->1	J->5	K->1	L->3	M->3	N->1	O->1	P->1	R->2	S->2	U->1	V->6	Å->3	
te:	 ->2	
te?	F->1	H->2	I->1	S->1	
tea	t->1	u->3	
teb	a->1	e->14	o->1	
tec	k->47	
ted	e->3	t->4	
tee	n->8	r->1	
tef	e->1	r->3	ö->6	
teg	 ->55	,->3	.->2	e->7	i->63	o->8	r->42	å->1	
tei	n->3	
tek	e->2	n->52	o->1	t->4	
tel	 ->6	a->2	e->7	i->1	l->27	n->1	s->31	t->1	ä->4	
tem	 ->75	,->9	.->11	:->1	a->19	b->15	e->90	o->27	p->6	ä->37	
ten	 ->828	!->4	"->4	)->3	,->112	.->167	:->2	;->2	?->2	F->1	H->1	N->1	a->10	b->4	d->17	e->19	f->2	h->3	k->1	l->1	p->1	r->2	s->164	t->17	v->8	
teo	r->2	
tep	o->1	r->1	
ter	 ->1017	!->15	"->2	)->2	,->114	-->3	.->153	:->3	;->2	?->4	H->1	a->537	b->4	d->42	e->1	f->27	g->16	h->9	i->178	k->8	l->64	m->14	n->713	o->1	p->4	r->178	s->289	t->17	u->34	v->83	å->1	
tes	 ->16	,->1	-->1	.->4	a->1	e->3	g->3	i->3	l->19	s->12	t->17	y->1	
tet	 ->812	!->1	"->2	,->91	-->1	.->94	:->4	?->5	e->76	i->2	s->156	
teu	r->9	
tex	t->45	
tfa	l->7	r->90	s->3	t->2	
tfe	d->1	
tfl	a->1	e->1	i->1	y->1	
tfo	r->42	
tfr	a->1	å->16	
tfu	l->15	
tfä	l->8	r->20	s->2	
tfå	n->1	
tfö	l->12	r->114	
tga	v->1	
tgi	c->1	f->16	l->8	v->2	
tgj	o->4	
tgr	u->7	
tgä	r->245	
tgå	 ->4	.->2	e->14	n->18	r->8	v->1	
tgö	r->63	
th 	S->1	h->1	n->1	o->1	
th,	 ->1	
th-	B->7	
tha	n->2	r->3	v->1	
the	 ->3	n->6	r->2	t->5	
thi	e->2	
tho	m->3	
thu	 ->1	s->7	
thy	 ->1	
thä	l->1	r->4	
thå	l->11	
thö	r->1	
ti 	-->1	a->1	d->2	f->10	g->1	h->4	i->9	k->3	m->2	o->12	p->2	s->9	t->2	u->1	v->1	å->1	
ti!	 ->3	
ti"	 ->1	
ti,	 ->14	
ti-	g->1	i->1	r->1	
ti.	.->1	D->3	E->2	F->1	H->3	I->1	J->1	K->2	M->1	V->1	
tia	l->3	n->1	t->80	
tib	e->11	
tic	a->1	e->4	h->1	k->5	
tid	 ->196	,->16	.->15	:->1	a->23	e->124	i->152	l->4	n->6	p->10	s->55	t->6	
tie	-->1	b->1	d->2	l->11	m->3	n->4	r->38	t->33	u->1	ä->2	
tif	a->3	i->36	o->3	r->18	t->128	
tig	 ->109	,->8	.->11	?->1	a->227	d->12	e->4	g->1	h->182	i->2	l->4	m->1	t->197	
tih	o->1	
tii	n->1	
tik	 ->127	!->1	"->1	,->31	.->25	?->2	a->11	e->255	l->15	o->7	r->3	s->1	
til	 ->3	a->1	e->2	i->1	l->2685	
tim	a->11	e->6	i->10	m->11	t->4	u->11	ö->1	
tin	 ->15	,->2	.->5	a->15	d->2	e->13	g->96	i->4	k->3	m->1	n->2	o->5	r->2	s->13	u->2	v->1	
tio	 ->15	e->1	f->1	n->1254	p->3	s->1	t->7	
tip	e->1	r->2	
tiq	u->2	
tir	e->1	
tis	 ->7	,->1	.->1	d->2	e->22	h->1	k->588	m->7	p->1	t->9	y->1	
tit	 ->7	a->4	e->9	i->7	r->1	s->8	t->22	u->159	y->5	
tiv	 ->211	,->23	.->23	:->2	;->1	?->2	a->133	b->1	e->144	f->4	i->42	l->2	r->5	t->114	
tiö	s->12	
tja	 ->18	d->4	n->9	r->3	s->6	t->2	
tjo	c->2	
tju	g->4	s->1	
tjä	m->8	n->173	r->3	
tka	n->1	s->15	t->1	
tkl	a->1	
tko	m->21	n->18	s->2	
tkr	a->1	i->1	ä->3	
tku	b->1	s->2	
tkv	ä->1	
tkä	l->1	
tkö	t->3	
tla	g->1	n->21	
tle	 ->3	.->1	k->1	r->6	v->1	
tli	g->530	n->76	s->2	
tlo	v->3	
tlä	g->4	m->2	n->16	
tlå	t->2	
tlö	s->5	
tma	k->1	n->22	r->2	t->1	
tme	d->2	r->1	
tmi	n->27	s->1	
tmo	n->1	
tmy	n->4	
tmä	n->2	r->32	s->1	t->1	
tmå	l->1	
tna	 ->35	,->3	.->6	d->109	r->8	s->3	
tne	 ->2	n->3	r->28	s->1	t->6	
tni	n->648	s->14	
tnj	u->1	
tny	t->42	
tnä	m->8	t->1	
to 	-->1	a->1	f->3	h->2	i->1	k->1	o->2	s->2	t->1	v->1	ö->1	
to-	a->1	p->1	
to.	J->1	V->1	
to/	O->1	
toa	k->1	n->1	
tob	a->3	e->9	
toc	k->3	
tod	 ->28	e->16	o->1	
tog	 ->42	a->2	e->2	s->22	
tok	o->26	
tol	 ->7	.->2	a->25	e->64	i->4	k->26	p->1	s->13	t->11	v->1	
tom	 ->99	!->1	)->1	,->5	.->1	a->8	e->6	f->1	m->1	o->7	r->8	s->2	
ton	 ->33	,->1	-->1	.->3	/->2	?->1	a->46	d->3	e->30	g->1	h->1	i->1	s->4	v->4	å->1	
top	-->1	i->1	p->31	r->2	
tor	 ->127	,->10	.->8	a->177	b->15	c->4	d->3	e->45	f->2	g->1	h->2	i->92	k->3	l->1	m->29	n->55	p->3	s->17	t->44	v->4	
tos	 ->14	
tot	a->34	
tow	n->3	
tox	i->1	
tpa	r->9	
tpe	k->1	n->1	r->10	
tpl	a->4	å->2	
tpo	l->3	s->10	
tpr	a->1	e->1	i->1	o->4	ä->1	
tpu	n->3	
tra	 ->73	,->1	d->26	f->50	g->10	k->36	l->79	m->5	n->151	o->1	p->3	r->33	s->20	t->112	u->1	v->2	x->3	
tre	 ->133	,->5	.->6	:->1	a->11	c->1	d->80	g->2	k->1	l->1	m->31	n->1	p->5	r->31	s->126	t->8	v->3	
tri	 ->11	,->3	-->1	b->1	c->7	d->23	e->8	f->4	k->44	l->3	n->104	o->2	p->2	s->3	
tro	 ->12	.->1	a->12	d->9	e->58	f->90	g->2	j->1	l->192	n->14	p->2	r->151	s->2	t->54	u->1	v->19	
tru	e->5	k->187	m->63	n->4	p->3	s->9	t->1	
try	c->101	g->8	k->34	m->11	p->1	
trä	 ->2	c->32	d->161	f->117	n->69	p->1	s->1	t->15	v->32	
trå	d->4	e->1	k->3	l->5	n->2	
trö	g->1	j->1	k->3	m->19	s->4	t->2	
ts 	"->2	(->1	-->9	8->1	B->1	E->1	L->1	S->2	a->126	b->34	c->2	d->50	e->17	f->101	g->39	h->23	i->64	k->13	l->14	m->42	n->12	o->67	p->34	r->24	s->51	t->46	u->45	v->16	y->3	ä->9	å->5	ö->4	
ts!	F->1	
ts,	 ->48	
ts-	 ->12	b->1	
ts.	A->1	B->1	D->20	E->6	F->1	H->2	I->1	J->5	K->3	M->2	N->1	R->2	S->4	T->1	V->3	Ä->1	
ts:	 ->1	
ts?	F->1	K->1	
tsa	 ->7	k->5	m->25	n->12	r->9	s->7	t->87	v->2	
tsb	a->4	e->12	u->1	ö->5	
tsc	e->2	h->4	
tsd	e->1	o->4	
tse	 ->11	.->1	d->4	e->1	k->2	l->5	n->31	r->81	s->3	t->4	
tsf	a->11	i->1	l->15	o->3	r->10	å->1	ö->12	
tsg	a->3	i->8	r->8	
tsh	a->2	j->2	
tsi	f->2	g->1	k->5	n->5	t->2	
tsk	a->7	i->10	l->2	o->167	r->9	u->1	y->8	
tsl	a->20	e->28	i->138	o->4	ä->15	å->17	ö->43	
tsm	a->15	e->4	i->2	y->10	ä->2	å->2	
tsn	i->10	o->6	ä->1	
tso	f->2	l->1	m->6	r->16	s->5	
tsp	a->5	e->2	l->11	o->7	r->87	å->2	
tsr	a->3	e->6	i->1	u->3	ä->4	å->18	
tss	a->1	e->5	i->2	k->5	p->1	t->34	y->23	ä->21	
tst	a->52	i->50	j->1	r->34	y->3	ä->55	å->13	ö->3	
tsu	g->1	t->7	
tsv	a->19	e->2	i->5	ä->4	
tsy	n->1	s->1	
tsä	g->10	k->8	t->152	
tså	 ->61	,->2	g->3	t->2	
tt 	"->2	(->2	-->11	1->3	2->2	4->1	5->1	7->1	8->2	9->1	A->4	B->6	C->1	D->3	E->107	F->7	G->1	H->1	I->7	J->3	K->3	M->2	N->1	O->3	P->3	R->3	S->3	T->16	V->1	a->443	b->426	c->5	d->1136	e->280	f->652	g->352	h->231	i->305	j->101	k->399	l->215	m->498	n->153	o->204	p->265	r->207	s->784	t->349	u->333	v->648	w->1	y->19	z->1	ä->103	å->83	ö->91	
tt,	 ->85	
tt.	 ->3	.->2	A->2	B->1	D->30	E->3	F->7	H->9	I->4	J->13	K->3	L->4	M->12	N->3	O->3	P->4	S->4	T->1	U->1	V->7	Ä->3	
tt:	 ->6	
tt?	A->1	D->1	O->1	S->1	V->1	
ttB	e->1	
tta	 ->1218	!->2	,->47	.->85	:->1	?->1	c->3	d->24	g->18	l->98	n->70	r->87	s->59	t->35	v->7	
tte	 ->27	,->1	-->2	b->15	d->1	f->3	g->1	i->2	l->5	n->227	p->1	r->236	s->10	t->163	
ttf	r->1	u->1	ä->7	ö->1	
ttg	ö->1	
tth	å->9	
tti	 ->1	c->1	d->1	g->169	l->47	n->2	o->2	s->16	t->6	
ttj	a->41	ä->25	
ttk	r->1	v->1	
ttl	a->5	e->4	i->2	
ttm	ä->1	å->1	
ttn	a->15	e->11	i->287	
tto	 ->2	-->1	a->1	l->1	n->9	r->3	
ttr	a->105	e->79	i->21	y->72	ä->5	
tts	 ->37	,->3	-->1	.->7	a->4	b->6	d->1	f->2	h->2	i->2	k->9	l->135	m->2	o->8	p->4	r->3	s->53	t->4	v->4	
ttv	i->75	
tty	s->2	
ttä	n->1	
tté	 ->10	e->4	f->2	n->41	s->2	
ttö	m->5	
tu 	m->21	
tua	l->1	t->129	
tud	 ->1	e->5	i->9	
tue	l->55	r->3	
tuf	f->2	
tug	a->26	i->70	o->1	u->1	
tul	a->6	e->33	l->4	
tum	 ->75	,->3	.->4	e->3	m->3	
tun	c->1	d->17	g->18	i->2	n->5	
tur	 ->67	,->19	-->2	.->10	?->1	a->9	b->1	e->136	f->61	h->1	i->25	k->22	l->102	m->1	n->2	o->2	p->20	r->1	s->8	u->3	v->1	å->1	
tus	 ->4	.->1	?->1	e->17	f->1	i->3	
tut	i->158	s->12	v->2	
tva	k->1	l->1	p->1	r->3	
tve	c->238	k->29	r->30	t->7	
tvi	d->107	k->6	l->2	n->33	s->215	v->43	
tvu	n->11	
tvä	n->1	r->51	t->5	
två	 ->122	.->1	:->2	h->1	n->6	
ty 	E->1	d->4	i->1	n->2	p->2	v->2	ä->1	
ty-	p->1	
tyc	k->94	
tyd	 ->4	.->1	a->17	d->3	e->97	i->11	l->124	
tyg	 ->35	)->1	,->3	.->4	;->1	?->1	a->37	e->25	s->13	
tym	p->3	
tyn	a->1	g->10	
typ	 ->20	,->2	.->2	e->16	f->1	g->1	
tyr	 ->1	.->1	a->20	e->16	k->17	n->7	s->2	
tys	k->25	t->3	
tyv	ä->30	
tz 	i->1	o->1	s->1	
tz,	 ->1	
tz.	 ->1	
tzi	d->2	
täc	k->31	
täd	a->2	e->19	
täk	t->5	
täl	l->426	
täm	d->19	l->3	m->187	n->2	p->2	s->1	t->16	
tän	 ->1	d->114	g->11	k->377	
täp	p->4	
tär	 ->6	,->1	.->1	a->11	e->4	k->51	t->2	
tät	a->2	e->2	h->1	
täv	 ->1	j->1	l->3	
tå 	a->16	d->3	e->1	f->21	h->2	i->5	k->4	n->2	o->3	s->1	t->1	u->2	v->4	
tå,	 ->3	
tå.	F->1	J->1	
tå:	 ->1	
tåd	d->2	
tåe	l->14	n->32	
tåg	 ->1	,->1	e->1	k->1	o->1	
tål	 ->1	a->2	f->5	g->1	i->27	s->6	v->5	
tån	d->226	
tår	 ->177	,->3	.->3	e->10	
tås	 ->6	
tåt	"->1	g->3	t->30	
té 	-->2	e->1	f->3	h->1	m->1	s->2	
tée	r->4	
téf	ö->2	
tén	 ->23	,->4	.->2	?->1	s->11	
tés	y->2	
têt	e->3	
tón	i->1	
töd	 ->160	,->14	.->38	;->1	?->1	d->2	e->122	j->72	m->2	n->1	p->1	r->2	s->13	å->5	
tök	a->11	n->1	
töl	d->1	
töm	d->1	m->4	t->1	
tör	 ->5	,->1	a->5	d->3	e->31	i->2	n->5	r->75	s->41	t->3	
töt	a->3	e->2	f->1	t->13	
töv	a->15	e->21	n->1	
tür	k->1	
u -	 ->1	
u 3	4->1	
u A	h->2	n->1	
u B	e->1	
u E	g->1	r->1	
u F	r->1	
u L	y->1	
u M	c->1	o->1	
u P	e->1	l->1	
u R	e->3	
u S	c->3	u->1	
u T	h->1	
u W	a->1	
u a	b->1	l->6	n->4	t->8	v->2	
u b	a->3	e->6	l->4	
u c	o->1	
u d	e->6	i->3	u->1	ä->1	å->1	ö->1	
u e	f->1	g->1	m->1	n->13	t->8	u->1	
u f	a->2	i->4	l->1	r->3	å->4	ö->17	
u g	e->5	ä->3	å->4	ö->3	
u h	a->19	o->1	ä->1	å->3	ö->5	
u i	 ->4	g->1	n->50	s->1	
u k	a->7	o->52	
u l	e->2	i->1	y->1	ä->4	
u m	e->35	i->3	o->1	ä->1	å->10	
u n	u->1	ä->8	å->1	
u o	c->14	f->3	m->1	
u p	a->1	l->1	o->1	r->2	u->1	å->5	
u r	e->3	u->1	å->2	ö->1	
u s	a->6	e->2	i->2	k->7	l->1	m->1	o->2	p->1	t->14	v->1	ä->2	å->2	
u t	a->88	i->5	y->3	
u u	n->1	p->3	t->1	
u v	a->1	e->3	i->7	ä->1	
u ä	l->1	n->8	r->24	
u å	t->2	
u",	 ->1	
u, 	L->1	a->1	e->3	h->1	i->1	m->2	o->2	p->1	s->3	u->1	å->1	ö->1	
u-l	ä->1	
u..	T->1	
u.D	e->1	
u.E	t->1	
u.J	a->1	
u.K	o->2	
u.L	å->1	
u.V	i->2	
u: 	g->1	
u; 	i->1	
u?J	a->1	
uMe	d->1	
ua 	n->2	
uad	e->1	
ual	 ->6	"->1	,->1	i->3	
uan	z->1	
uar	i->32	
uat	e->1	i->129	
ubb	a->3	e->6	l->11	
ube	t->1	
ubi	k->2	
ubj	e->1	
ubl	a->1	i->33	
ubr	i->2	
ubs	i->23	t->4	
ubv	e->12	
uc 	s->1	
ucc	e->5	
uce	n->22	r->13	
uch	n->12	
uck	a->3	i->1	n->1	o->2	
uct	o->1	
ud 	7->1	B->2	e->1	f->5	m->9	o->4	r->1	t->9	v->1	ä->1	
ud,	 ->4	
ud.	D->2	V->1	
uda	 ->15	k->2	n->10	p->1	r->1	s->2	
udd	a->2	e->3	h->1	i->2	
ude	 ->1	n->3	r->19	t->14	u->1	
udf	r->4	ö->1	
udg	e->107	
udi	c->1	e->9	k->3	s->1	t->1	
udl	i->3	
udm	å->2	
udn	a->2	i->1	
udo	r->1	
udr	e->3	o->3	
uds	 ->2	a->16	f->3	i->3	k->10	m->10	p->1	t->4	y->1	
udu	p->1	
ue 	k->1	
ue,	 ->2	
uec	e->1	
uei	r->1	
uel	a->1	l->67	
uen	,->1	
uer	 ->3	,->1	a->8	l->2	n->1	
ues	 ->4	"->1	a->1	
uff	 ->1	a->1	
ufm	a->1	
uft	 ->1	.->1	b->1	e->1	i->11	o->1	
ufö	r->1	
uga	,->1	l->26	r->1	
uge	n->2	r->1	
ugg	 ->3	a->2	b->1	e->1	l->1	
ugi	s->70	
ugl	i->6	
ugn	 ->1	a->5	
ugo	 ->2	f->1	n->1	r->1	s->1	
ugu	e->1	
uha	m->1	
uhe	 ->1	,->1	
uhn	e->1	
uie	r->1	
uig	o->1	
uin	e->1	s->1	
uio	l->1	
uis	e->3	i->1	
uit	a->1	
uiz	 ->1	
uk 	a->2	m->1	o->5	p->1	s->1	
uk!	A->1	
uk,	 ->9	
uk.	J->1	
uka	 ->1	,->1	d->2	r->17	s->5	
ukd	o->1	
uke	n->1	t->19	
ukf	ö->1	
ukh	u->7	
uki	t->1	
ukn	i->3	
uks	e->1	f->2	l->1	o->2	p->9	r->2	s->6	
ukt	 ->7	,->1	.->1	a->12	b->2	e->17	i->62	o->6	s->2	u->153	ö->3	
ukv	å->3	
ul 	f->1	o->2	s->1	
ul.	V->1	
ula	 ->2	.->1	d->1	n->5	r->2	t->14	
uld	a->2	b->1	e->3	
ule	n->1	r->64	
ulf	-->2	e->1	k->1	
ulg	a->1	
uli	 ->8	,->2	s->5	
ulk	l->1	
ull	 ->28	,->3	.->6	a->29	b->3	e->486	f->4	g->3	h->1	i->1	k->6	o->5	s->44	t->43	v->2	ä->2	
ulo	r->1	s->5	
uls	 ->2	e->4	k->1	
ult	 ->2	a->111	b->1	e->29	h->6	i->10	r->2	u->146	
ulz	 ->3	
ulä	g->1	r->3	
um 	-->1	a->59	b->1	d->1	e->2	f->11	h->3	i->22	m->4	o->12	p->4	s->8	u->2	v->1	y->1	ä->5	å->2	
um!	D->1	M->1	
um,	 ->12	
um.	 ->1	A->2	D->4	H->1	I->1	L->1	M->1	O->1	P->1	R->1	S->1	V->2	Ä->1	
uma	n->6	r->1	t->1	
umb	a->1	ä->4	
ume	n->176	r->6	t->6	
umg	ä->1	
umh	e->3	
uml	e->1	
umm	a->9	e->8	i->1	o->8	
ump	 ->3	.->1	a->3	e->2	n->3	
umr	a->1	
umt	 ->1	a->1	i->2	
umu	l->2	
umä	n->1	
umö	r->2	
un 	s->1	
un.	D->1	
una	 ->2	l->3	n->1	
unc	 ->1	h->1	i->1	
und	 ->119	,->2	.->3	?->1	a->104	b->1	e->585	f->4	g->3	i->6	k->1	l->90	n->4	o->1	p->2	r->36	s->11	t->1	v->65	ä->1	
une	r->11	
ung	 ->9	.->3	a->24	d->14	e->71	f->1	l->13	m->6	n->6	r->1	s->1	t->2	
unh	a->1	
uni	 ->12	c->2	k->18	l->2	o->437	s->3	t->1	v->4	
unk	a->4	e->3	i->2	l->1	n->4	t->377	
unn	a->259	e->6	i->22	l->2	o->1	
uno	 ->1	
uns	k->17	
unt	 ->4	.->1	a->7	l->8	o->2	p->1	r->21	
uo 	s->1	
uo,	 ->1	
up 	,->1	d->1	ö->1	
upa	 ->5	,->1	d->1	n->1	r->1	s->3	t->3	
upe	r->3	t->5	
upg	å->7	
upn	i->5	
upp	 ->252	,->20	.->19	?->1	b->26	d->27	e->168	f->129	g->88	h->29	k->7	l->25	m->136	n->93	o->1	r->110	s->84	t->34	u->1	v->8	
upr	a->1	
ups	i->1	k->1	
upt	 ->7	i->7	
upé	r->1	
uqa	l->2	
ur 	-->2	2->20	E->4	U->1	a->5	b->15	d->49	e->16	f->15	g->4	h->6	i->6	j->1	k->17	l->11	m->36	n->5	o->10	p->9	r->1	s->56	t->5	u->9	v->34	ä->6	
ur,	 ->21	
ur-	 ->4	
ur.	D->4	F->1	H->1	K->1	N->1	O->1	R->1	T->1	V->3	
ur?	M->1	
ura	 ->6	,->2	.->1	k->1	l->1	n->12	r->9	s->1	t->5	
urb	a->1	e->1	
urd	 ->1	
ure	l->40	n->55	r->43	s->1	t->2	
urf	o->63	ö->2	
urg	 ->6	,->4	.->4	a->1	h->1	
urh	i->1	o->4	
uri	.->1	d->30	e->2	s->41	t->2	
urk	-->1	a->15	i->41	m->2	
url	a->6	i->104	
urm	i->1	ä->1	
urn	a->3	e->1	ä->1	ö->1	
uro	 ->16	!->1	,->8	-->1	.->8	d->5	f->1	j->6	m->2	n->7	o->1	p->1207	s->4	
urp	o->16	r->4	
urr	e->287	
urs	 ->5	,->1	.->1	b->1	e->61	f->1	k->4	p->20	s->1	t->4	ä->15	
urt	 ->2	z->3	
uru	t->3	v->15	
urv	a->13	e->1	i->1	
urå	t->1	
us 	1->1	2->1	a->2	b->3	e->2	f->2	h->1	j->5	k->2	o->3	p->1	q->2	s->2	t->2	u->1	ä->1	
us,	 ->5	
us-	b->1	
us.	D->2	E->1	G->1	H->1	I->1	
us?	O->1	
usa	 ->1	l->2	r->2	
usc	h->1	
usd	i->1	
use	"->1	f->3	n->19	r->3	t->11	w->1	
usf	ö->1	
usg	a->4	r->2	
ush	 ->1	,->1	å->1	
usi	a->3	k->4	o->8	v->20	
usk	.->1	o->1	
usl	ä->1	
usp	"->1	e->1	
usq	u->1	
uss	a->5	e->3	i->62	l->2	
ust	 ->101	,->1	.->3	:->1	a->4	b->3	e->39	i->10	l->2	m->3	n->5	o->2	r->117	v->1	
usu	l->6	
usí	 ->1	
usö	v->1	
ut 	-->1	1->1	8->2	9->1	T->1	a->15	b->7	d->8	e->8	f->20	g->2	h->7	i->20	k->5	l->4	m->11	n->14	o->32	p->30	r->3	s->24	t->5	u->6	v->3	ä->4	å->1	ö->5	
ut,	 ->34	
ut.	 ->2	(->1	)->1	D->9	F->4	G->1	I->1	J->5	K->1	N->2	O->1	S->2	T->1	V->2	Ä->1	
ut:	 ->1	
ut;	 ->1	
ut?	.->1	E->1	
uta	 ->55	,->5	b->3	d->30	f->10	l->2	n->357	p->1	r->50	s->13	t->14	u->3	
utb	a->1	e->8	i->60	r->4	u->4	y->20	
utd	e->1	
ute	 ->4	a->3	l->3	n->21	r->104	s->23	t->57	
utf	a->4	l->2	o->40	r->7	ä->13	ö->46	
utg	a->1	i->25	j->4	å->29	ö->59	
uth	a->1	e->1	ä->4	
uti	e->1	f->16	k->1	n->8	o->260	q->1	t->11	
utj	ä->5	
utk	a->16	o->4	r->3	
utl	a->5	i->72	o->3	ä->7	å->2	ö->2	
utm	a->20	y->1	ä->32	
utn	a->17	i->41	y->41	ä->4	
uto	/->1	m->100	p->1	r->1	
utp	e->2	l->2	r->2	u->1	
utr	a->2	e->13	i->19	o->7	u->4	y->11	ä->2	
uts	 ->6	-->1	a->65	c->2	e->17	f->12	i->2	k->157	l->24	p->4	r->1	t->43	u->1	ä->63	å->3	
utt	a->100	e->2	i->2	j->24	n->2	o->5	r->73	ö->5	
utv	a->4	e->241	i->107	ä->32	
uty	p->1	
utä	n->5	
utå	t->1	
utö	k->12	v->30	
uum	 ->1	t->1	
uva	 ->1	r->46	
uve	l->2	r->19	
uvi	d->15	
uvr	i->1	
uvu	d->54	
ux,	 ->2	
ux-	a->1	
uxe	m->6	
uxh	a->1	
uxi	t->1	
uxn	a->2	
uyu	 ->2	
v "	p->1	r->2	
v (	K->1	
v -	 ->9	
v 1	4->1	9->3	
v 2	0->1	
v 4	0->1	1->1	
v 5	 ->1	4->1	
v 8	 ->1	
v 9	3->1	4->2	6->5	
v A	h->2	m->2	r->1	
v B	N->6	S->1	a->2	e->8	o->1	r->2	
v C	a->1	
v D	a->2	e->1	i->2	u->1	ü->1	
v E	G->1	U->17	n->1	r->1	u->70	x->2	
v F	N->1	P->2	l->1	ö->8	
v G	a->1	e->2	r->3	
v H	a->1	e->1	i->1	
v I	s->2	
v J	a->1	e->1	o->2	
v K	i->3	o->10	u->1	
v L	a->3	i->1	ö->1	
v M	a->2	c->1	o->1	
v O	L->3	s->1	z->1	
v P	a->2	o->1	é->1	
v R	a->1	i->1	
v S	a->1	c->6	
v T	a->1	e->1	h->4	i->1	o->1	
v U	N->1	
v V	a->2	ä->1	
v W	a->1	i->1	y->1	
v a	c->1	d->2	g->1	l->36	n->31	p->2	r->40	s->1	t->70	v->29	
v b	a->3	e->42	i->15	l->4	o->3	r->10	u->8	y->2	å->2	ö->3	
v c	e->2	i->6	o->1	
v d	a->6	e->561	i->29	j->2	o->12	r->1	ä->2	
v e	f->5	g->2	k->12	n->114	r->18	t->52	u->7	v->1	x->8	
v f	a->49	i->6	j->2	l->16	o->8	r->36	u->5	y->1	ä->1	å->5	ö->125	
v g	a->3	e->32	i->3	l->1	o->2	r->11	ö->1	
v h	a->20	e->7	i->5	j->1	o->1	u->8	ä->2	ö->3	
v i	 ->15	b->1	c->3	d->2	m->5	n->37	
v j	o->5	u->4	ä->2	
v k	a->13	l->4	n->1	o->119	r->5	u->5	v->7	ä->8	
v l	a->21	e->12	i->16	o->5	ä->5	å->1	ö->2	
v m	a->18	e->31	i->40	o->6	y->3	ä->7	å->8	ö->1	
v n	a->14	i->1	o->1	y->13	ä->2	å->6	ö->2	
v o	a->3	b->4	c->29	f->5	k->1	l->14	m->33	n->1	p->1	r->11	s->12	t->2	u->1	v->1	
v p	a->22	e->12	i->1	o->9	r->37	å->33	
v r	a->6	e->33	i->8	o->2	y->1	ä->12	å->12	ö->1	
v s	a->16	c->1	e->10	i->25	j->3	k->23	l->2	m->2	n->1	o->46	p->2	t->81	u->4	v->2	y->24	ä->15	å->15	
v t	a->4	e->8	i->40	j->28	o->2	r->13	u->6	v->2	y->2	ä->1	
v u	n->30	p->6	t->37	
v v	a->23	e->10	i->26	o->4	ä->20	å->24	
v y	t->5	
v Ö	s->2	
v ä	l->1	m->1	n->6	r->9	
v å	l->1	r->8	s->1	t->16	
v ö	b->1	d->1	k->4	p->4	s->2	v->4	
v",	 ->1	
v, 	9->1	a->3	b->1	d->5	e->3	f->1	h->4	i->1	j->1	l->1	m->5	n->2	o->8	s->8	t->2	u->1	ä->2	
v. 	D->1	M->1	V->2	m->1	
v."	D->1	
v.(	S->1	
v.,	 ->1	
v..	 ->2	H->1	
v.?	A->1	
v.A	t->1	v->2	
v.B	a->1	l->1	
v.D	e->11	ä->1	å->1	
v.E	f->1	n->2	r->1	
v.F	r->1	ö->4	
v.H	e->1	
v.I	 ->2	n->1	
v.J	a->2	
v.K	o->1	
v.L	å->1	
v.M	e->3	
v.O	L->1	m->1	
v.R	i->1	å->1	
v.S	v->1	å->1	
v.U	p->1	
v.V	i->3	
v.Y	t->1	
v: 	F->1	v->1	
v; 	a->1	
v?F	ö->1	
v?N	e->1	
v?V	i->1	
va 	4->1	E->2	a->18	b->14	c->1	d->23	e->28	f->16	g->5	h->6	i->15	j->1	k->21	l->5	m->8	n->5	o->18	p->15	r->12	s->20	t->18	u->7	v->33	ä->2	å->8	ö->3	
va,	 ->9	
va.	A->1	D->1	H->1	L->1	N->1	O->1	V->2	
va?	N->1	
vac	k->9	
vad	 ->238	?->1	e->12	
vag	 ->3	a->30	h->12	n->3	t->1	
vak	a->19	i->1	n->14	s->9	t->8	u->2	
val	 ->35	,->3	.->5	;->1	a->3	b->1	d->34	e->13	f->5	i->51	k->4	l->2	r->1	s->1	t->61	u->23	
van	 ->41	,->1	.->2	a->2	c->1	d->64	h->2	i->1	l->12	n->2	o->3	p->1	s->15	t->18	
vap	e->26	n->2	
var	 ->351	,->30	.->43	;->1	?->1	a->580	d->5	e->147	f->39	g->1	h->3	i->136	j->84	k->15	l->63	m->15	n->30	o->10	p->1	r->1	s->119	t->10	v->8	
vas	 ->23	,->2	.->6	t->1	
vat	 ->13	.->2	a->18	e->1	i->19	s->6	t->49	ö->1	
vav	t->7	
vbe	s->3	t->1	
vbi	o->1	
vbo	r->1	
vbr	i->1	o->4	u->2	y->3	ö->6	
vbä	r->1	
vda	 ->7	d->3	r->12	t->5	
vde	 ->5	,->1	l->8	s->2	
vdv	u->1	
ve 	(->2	1->1	E->1	a->2	b->4	d->4	e->3	f->1	k->4	l->2	m->3	p->3	r->3	s->1	t->2	ä->1	
ve,	 ->2	
ve-	 ->1	p->2	
veN	ä->1	
veb	r->1	
vec	 ->1	k->289	
ved	e->13	
vek	 ->2	a->24	h->4	l->1	o->1	s->5	
vel	 ->26	,->2	a->10	e->2	s->9	
vem	 ->17	b->11	s->1	
ven	 ->363	,->4	.->9	:->1	e->3	h->4	s->50	t->90	
vep	 ->1	e->1	s->1	t->1	
ver	 ->396	,->8	.->14	a->43	b->10	c->1	d->14	e->77	f->23	g->47	h->5	i->23	k->588	l->35	m->2	n->5	o->1	p->1	r->4	s->96	t->57	v->72	y->1	ä->17	
ves	 ->2	t->18	
vet	 ->236	"->1	,->28	.->26	a->32	e->105	n->17	s->13	t->5	v->27	y->7	
veu	r->1	
vfa	l->25	
vfo	l->1	
vfö	r->8	
vga	s->1	v->1	
vge	 ->3	r->5	s->1	t->1	
vgi	c->4	f->4	v->1	
vgj	o->4	
vgr	ä->4	
vgå	.->1	e->1	n->3	r->1	t->1	
vgö	r->61	
vhe	t->1	
vhj	ä->4	
vhä	n->2	
vhå	l->1	
vi 	-->3	1->1	5->1	E->2	I->1	L->1	P->1	a->128	b->108	d->56	e->44	f->97	g->52	h->175	i->194	j->11	k->123	l->27	m->90	n->35	o->44	p->15	r->28	s->161	t->62	u->38	v->74	y->1	ä->47	å->7	ö->8	
vi,	 ->16	
vi.	V->1	
vi?	.->1	
via	 ->12	n->1	
vic	 ->1	e->20	k->3	
vid	 ->217	,->2	.->2	a->58	d->5	e->22	g->109	h->5	l->1	m->1	s->1	t->64	u->8	
vie	n->2	r->1	
vif	t->1	
vig	 ->1	l->1	t->3	v->1	ö->1	
vik	a->35	e->14	i->1	l->4	n->1	t->365	
vil	 ->5	-->1	a->6	b->2	d->1	e->6	f->2	i->3	j->229	k->317	l->633	r->1	s->5	t->2	
vin	 ->2	d->5	g->32	i->1	k->12	n->161	s->15	
vir	k->3	r->13	
vis	 ->237	)->1	,->17	.->9	a->235	b->17	d->1	e->20	f->3	h->3	i->24	k->4	m->1	n->14	o->5	s->196	t->27	u->3	
vit	 ->39	.->1	b->50	e->39	s->10	t->7	
viv	e->33	l->10	
vja	s->1	
vje	t->1	
vju	 ->2	a->1	
vka	r->1	
vkl	a->21	
vko	n->1	s->1	
vkr	a->3	ä->1	
vku	n->1	
vla	 ->5	"->2	.->1	d->4	g->1	n->1	r->6	t->2	
vle	d->2	
vli	g->10	n->1	s->2	v->1	
vlo	p->1	
vlä	g->10	
vlå	d->1	
vma	t->1	
vmi	l->1	
vna	 ->9	d->16	
vni	n->36	
vo 	(->2	T->1	a->1	b->1	f->3	h->1	i->1	k->2	m->1	o->7	t->1	u->1	v->1	ä->3	
vo,	 ->11	
vo.	-->1	A->1	D->2	E->1	F->1	H->1	K->1	L->1	M->1	O->1	V->1	
vo?	 ->1	H->1	
voN	ä->1	
vof	f->1	
vok	a->5	o->1	r->1	
vol	u->5	v->9	y->4	
von	 ->18	
vor	 ->1	.->1	d->2	e->29	i->1	
vos	 ->7	
vot	 ->4	!->1	,->1	e->13	u->1	
voå	r->1	
vpl	å->1	
vpr	i->1	
vra	d->1	k->10	n->1	p->1	r->1	s->1	
vre	d->1	g->2	
vri	d->14	g->66	k->1	è->1	
vru	n->1	
vrä	k->1	n->2	t->5	
vs 	a->6	b->1	d->14	e->20	f->10	g->1	h->3	i->13	k->1	m->4	n->1	o->4	p->2	r->1	s->10	u->3	v->4	ä->1	ö->1	
vs,	 ->10	
vs.	 ->45	A->1	D->3	E->2	F->1	I->1	R->1	S->2	V->1	
vs?	T->1	
vsa	k->4	r->3	t->4	
vsc	y->3	
vsd	u->2	
vse	 ->1	d->3	e->47	r->15	s->1	t->14	v->14	
vsf	o->1	ö->1	
vsi	d->2	k->38	n->1	
vsk	a->19	e->5	i->1	o->3	r->3	v->5	y->2	
vsl	a->2	o->2	u->74	ä->2	å->3	ö->6	
vsm	a->2	e->88	i->5	ä->3	
vsn	i->4	
vso	m->1	
vsp	e->5	
vss	t->2	
vst	a->2	e->1	o->2	y->7	ä->11	å->26	
vsu	p->1	
vsv	a->1	i->1	
vsä	g->1	k->1	t->4	
vt 	-->1	a->11	b->4	d->4	e->4	f->8	h->3	i->9	k->4	m->4	n->1	o->17	p->6	r->4	s->33	t->7	u->2	v->1	y->1	ä->1	å->4	ö->1	
vt,	 ->7	
vt.	 ->1	D->2	E->1	I->1	P->1	Ä->1	
vta	l->89	r->1	
vti	d->1	m->2	
vtr	u->1	
vts	 ->2	.->1	
vtv	i->1	
vud	 ->9	a->7	d->3	e->1	f->5	l->2	m->2	r->3	s->21	u->1	
vul	e->1	s->1	
vun	d->1	g->11	n->11	
vux	i->1	n->2	
vva	k->6	
vve	c->8	r->2	
vvi	k->8	s->15	
vvä	g->5	r->2	
vyt	t->1	
väc	k->23	
väd	e->2	j->9	r->1	
väg	 ->33	,->16	.->9	N->1	a->55	b->1	d->3	e->27	g->3	l->5	m->1	n->17	r->23	s->7	t->2	
väk	a->1	t->2	
väl	 ->100	,->2	.->3	b->1	d->23	f->9	g->3	j->22	k->54	l->11	m->4	s->8	t->4	u->3	v->4	
väm	l->15	m->3	n->4	t->1	
vän	 ->1	d->341	l->15	n->3	s->16	t->88	
väp	n->2	
vär	d->168	e->1	l->61	n->3	p->2	r->49	s->9	t->41	v->7	
väs	e->36	t->4	
vät	s->1	t->5	
väv	a->2	n->4	t->1	
väx	a->9	e->10	l->4	t->32	
vå 	-->1	a->13	b->3	d->3	e->7	f->28	g->4	h->3	i->7	j->1	k->4	l->2	m->12	n->3	o->9	p->14	r->2	s->21	t->8	u->6	v->7	y->1	ä->3	å->8	
vå,	 ->13	
vå.	A->1	B->2	D->7	F->1	G->1	H->2	J->4	M->1	N->1	P->1	V->1	
vå:	 ->2	
vå;	 ->1	
vå?	S->1	
våd	l->1	
våe	r->14	
våg	 ->2	a->6	e->2	l->1	r->3	
våh	u->1	
vål	d->12	l->1	
vån	 ->8	.->4	a->17	g->7	i->2	
vår	 ->145	,->1	a->175	b->2	d->8	e->2	i->31	l->2	s->2	t->134	ö->1	
vö,	 ->1	
vö.	D->1	
vön	 ->1	
vör	d->1	
w Y	o->1	
w f	ö->1	
w t	i->1	
w, 	s->1	
w-h	o->1	
w.M	e->1	
wag	e->1	
wal	d->1	e->1	
wan	 ->1	
war	z->1	
we.	E->1	V->1	
web	b->1	
wei	z->1	
wel	l->1	
wer	 ->1	,->2	
wie	s->1	
wil	l->1	
wis	 ->2	
wit	t->1	z->1	
wn 	a->1	ä->1	
wn,	 ->1	
wob	o->3	
woo	d->3	
wor	s->1	
x a	l->1	n->4	v->2	
x e	f->1	u->1	
x f	l->1	
x i	n->1	
x m	i->1	å->10	
x o	c->1	
x p	l->1	o->1	
x s	a->1	
x t	i->1	u->1	
x ö	v->1	
x!J	a->1	
x, 	j->1	n->2	s->2	
x-a	f->1	
x-f	r->3	
x. 	E->1	F->1	N->1	U->1	a->2	d->2	e->1	i->1	k->2	m->2	n->2	o->1	p->1	u->1	v->1	
x.D	e->1	
x.J	a->1	
xa 	e->1	u->2	
xa,	 ->1	
xa.	H->1	M->1	
xak	t->18	
xal	 ->2	a->1	t->2	
xam	e->6	i->10	
xan	?->1	d->8	
xas	 ->7	
xat	 ->1	
xbe	l->1	
xce	p->6	
xel	k->1	r->1	v->2	
xem	b->6	p->118	
xen	 ->1	
xer	 ->6	,->1	i->1	
xfi	c->1	
xha	v->1	
xib	e->11	i->10	l->6	
xid	 ->4	u->1	
xik	o->1	
xil	r->1	t->1	
xim	a->6	e->2	i->1	
xin	 ->1	k->1	
xis	 ->5	.->2	e->1	k->1	m->1	t->19	
xit	 ->1	
xkl	u->3	
xla	n->1	r->2	
xli	n->2	
xmå	n->1	
xna	 ->1	.->1	
xni	n->1	
xon	 ->3	
xor	.->1	
xpa	n->6	
xpe	d->1	r->46	
xpl	i->1	o->2	
xpo	n->2	r->4	
xt 	a->2	f->1	i->1	k->1	l->1	o->7	s->6	ä->1	
xt,	 ->7	
xt.	K->1	M->1	O->1	
xtb	r->1	
xte	n->25	r->19	
xth	u->7	
xto	n->1	
xtr	a->7	e->30	
xts	k->3	
xue	l->3	
xup	é->1	
xvä	r->1	
xxo	n->3	
y -	 ->1	
y C	a->3	
y E	u->1	
y F	o->1	
y b	i->1	
y d	e->4	
y e	n->2	u->1	
y f	a->1	o->1	ö->6	
y g	r->1	
y h	a->2	ä->1	
y i	 ->1	n->3	
y k	e->1	o->3	u->3	v->1	
y l	a->1	e->1	i->1	
y m	y->1	
y n	a->1	ä->1	
y o	c->3	l->1	
y p	e->2	å->2	
y r	ö->2	
y s	e->1	i->1	o->1	p->1	t->1	y->2	
y t	y->1	
y u	n->1	p->1	
y v	a->1	e->1	i->6	
y ä	r->1	
y å	t->1	
y! 	G->1	
y, 	H->1	J->1	a->1	d->1	h->1	k->2	s->2	
y-p	r->1	
y.A	n->1	
y.D	e->1	
y.V	i->2	
yDe	 ->1	
ya 	"->1	8->1	E->3	Z->2	a->12	b->14	d->5	e->2	f->10	g->3	i->4	j->1	k->17	l->7	m->17	n->2	o->6	p->13	r->17	s->7	t->8	u->3	v->4	ä->2	å->6	
ya,	 ->1	
ya;	 ->1	
yab	e->1	u->2	
yag	o->4	
yal	 ->1	
yan	d->1	n->2	s->3	
yar	 ->1	b->1	
yas	 ->1	t->1	
yav	t->1	
yba	r->39	
ybe	t->2	
ybi	l->3	
yck	 ->24	,->2	.->1	a->112	b->1	e->552	l->34	n->5	o->17	s->20	t->21	ö->5	
ycl	i->1	
yd 	g->1	i->1	s->1	t->1	
yd.	S->1	
yda	 ->3	f->2	n->18	
ydd	 ->34	)->1	,->3	.->6	a->32	e->21	s->16	
yde	l->76	r->27	u->1	
ydi	g->11	
ydk	o->1	u->1	
ydl	i->125	
ydo	s->2	
yds	 ->1	
ydv	ä->1	
ydö	s->1	
ye 	P->1	o->1	
ye-	a->2	
yed	 ->2	
yel	s->6	
yen	s->1	
yer	 ->2	.->1	n->1	
yet	a->1	
yfa	l->1	s->1	
yft	 ->2	a->43	e->46	o->3	
yfö	r->2	
yg 	d->1	f->5	i->4	m->3	n->1	o->3	s->15	u->3	
yg)	,->1	
yg,	 ->4	
yg.	E->1	F->1	V->2	
yg;	 ->1	
yg?	D->1	
yga	 ->11	d->21	n->6	r->1	
ygb	l->1	
ygd	 ->2	.->2	e->31	s->10	
yge	l->5	n->13	r->1	t->8	
ygg	a->63	d->4	e->16	h->6	n->19	o->1	r->1	s->3	t->5	
ygi	e->2	
ygk	r->1	
ygn	i->1	
ygp	l->4	
ygr	u->2	
ygs	a->4	b->1	i->1	s->9	t->1	ä->1	
ygt	 ->3	r->2	
yhe	t->13	
yhu	n->1	
yhö	g->1	
yis	t->2	
yk.	H->1	
yka	 ->25	,->2	s->4	
yke	l->3	r->7	
ykl	a->4	
yko	l->1	
yks	 ->2	
ykt	a->2	b->1	e->12	i->13	r->1	
yl 	g->1	o->3	
yl,	 ->2	
yl-	 ->1	
yl.	D->1	J->1	V->1	
yla	.->1	n->1	
ylb	e->1	
yld	i->29	
ylf	ö->2	
yli	b->1	g->31	k->3	
yll	a->39	d->1	e->21	n->1	r->1	s->4	t->4	
ylr	ä->2	
yls	ö->6	
ym 	a->1	m->1	o->1	s->1	
ym.	D->1	
yma	 ->1	s->1	
ymb	o->9	
ymd	 ->1	e->1	
yme	n->1	r->1	
ymi	t->1	
ymm	a->1	e->17	
ymp	a->9	i->2	n->2	t->1	
ymr	a->10	
yms	 ->1	
ymt	 ->1	s->1	
yn 	-->1	a->2	g->1	h->1	i->2	l->1	o->5	p->4	t->65	v->1	ä->2	å->1	
yn,	 ->2	
yn.	A->1	E->1	S->2	
yn;	 ->1	
yna	 ->1	m->5	n->1	s->3	z->6	
ynd	 ->4	a->14	e->1	i->164	r->1	s->4	
yne	n->6	r->2	s->1	
yng	a->1	d->6	e->1	r->1	s->3	
ynl	i->8	
ynn	,->1	a->18	e->56	s->3	
yno	n->1	
ynp	u->29	
yns	 ->1	t->2	ä->4	
ynt	 ->2	,->1	e->1	
ynv	i->12	
yo 	s->1	
yol	a->2	
yon	 ->2	,->1	
yos	t->1	
yot	o->7	
yp 	C->1	a->18	f->1	
yp,	 ->2	
yp.	D->1	E->1	
ype	n->12	r->5	
ypf	a->1	
ypg	o->1	
yph	å->3	
ypl	a->1	
ypo	t->2	
ypp	a->1	e->1	
yps	.->1	
ypt	e->2	o->2	
yr 	a->1	e->1	f->1	h->1	j->1	
yr.	E->1	
yra	 ->37	,->1	:->1	m->1	n->4	r->7	s->2	
yrd	 ->1	
yre	 ->1	,->1	g->1	k->3	l->7	n->1	t->3	
yri	e->28	g->1	s->4	
yrk	a->16	e->20	o->3	
yrn	e->2	i->7	
yrs	 ->2	
yrt	 ->1	.->1	i->4	
yrå	 ->2	e->1	k->30	n->3	
ys 	-->1	a->16	b->3	d->1	f->3	g->1	i->1	j->1	o->3	s->1	v->1	
ys,	 ->4	
ys-	d->1	
ys.	D->2	F->1	G->1	H->1	
ys?	D->1	I->1	
ysa	 ->10	n->4	t->2	
yse	n->5	r->23	
ysi	s->9	
ysk	 ->1	a->23	l->22	t->2	
ysn	i->5	
yss	 ->10	,->2	.->1	a->2	e->127	l->10	n->29	
yst	 ->5	e->192	r->1	
yta	 ->13	.->1	n->13	s->1	
yte	 ->10	,->1	l->3	r->9	t->6	
yti	s->1	
ytl	i->2	
ytn	i->3	
yts	 ->1	
ytt	 ->42	,->3	.->4	a->31	e->91	i->13	j->41	n->4	o->2	r->43	s->1	
yu 	i->1	s->1	
yva	l->1	
yve	r->2	
yvä	r->40	
ywo	o->1	
yxf	i->1	
yår	s->1	
z F	i->3	l->2	
z G	o->1	
z a	n->1	
z b	e->1	
z d	y->1	
z e	l->1	n->1	t->1	
z f	r->1	å->1	ö->2	
z h	a->1	
z i	 ->1	
z o	c->8	m->1	
z s	a->2	o->2	
z t	o->2	
z)(	T->1	
z).	H->1	
z, 	G->1	L->3	b->1	i->1	p->1	t->1	u->1	
z-k	a->3	
z. 	E->1	
zFr	u->1	
za 	o->1	
za,	 ->1	
za.	D->1	S->1	
zak	s->1	
zar	e->2	
zbe	k->2	t->1	
zen	.->1	
zes	-->1	
zid	a->2	
zig	e->4	
zio	-->4	
zis	m->8	t->13	
zji	k->5	
zma	n->2	
zon	 ->4	e->3	i->1	
zor	e->2	
zqu	i->1	
zue	l->1	
zwa	l->1	
zál	e->1	
º C	.->1	
Ämn	a->1	
Än 	e->3	
Änd	a->1	r->14	å->5	
Änn	u->3	
Änt	l->1	
Är 	I->1	d->19	h->1	i->1	k->2	r->1	s->1	v->1	
Ära	d->6	
Äve	n->46	
Å E	D->1	
Å P	S->1	
Å a	n->10	
Å e	n->2	
Å k	o->1	
Å s	o->1	
ÅDS	K->1	
ÅGO	R->1	
År 	1->4	2->1	
Åre	t->1	
Årl	i->1	
Åta	g->1	
Åte	r->4	
Åtg	ä->5	
Île	-->1	
Ö (	Ö->2	
Ö f	ö->1	
Ö h	ä->1	
Ö i	n->1	
Ö m	i->1	
Ö o	c->3	m->1	
Ö s	o->1	
Ö v	i->1	
Ö ä	r->1	
Ö) 	s->1	
Ö).	J->1	
Ö-l	e->1	
Ö-m	e->1	
Ö:s	 ->4	
ÖST	N->2	
ÖVP	 ->5	)->1	
Ögo	n->2	
Öka	d->1	
Öpp	e->1	
Öst	e->86	t->2	
Öve	r->2	
Övr	i->1	
ále	z->1	
án,	 ->1	
ánc	h->1	
ão 	T->2	
ä u	t->1	
ä ö	v->1	
äck	 ->3	a->37	e->38	h->1	l->78	n->32	o->1	s->9	t->18	v->3	
äd 	b->1	f->1	h->2	u->1	
äd,	 ->1	
äd.	D->1	
äda	 ->11	,->1	n->10	r->57	t->1	
ädd	 ->5	,->1	a->14	e->7	n->4	
äde	 ->15	.->3	H->1	P->1	l->6	n->4	r->58	s->11	t->12	
ädj	a->17	e->7	
ädr	e->1	
äds	 ->8	l->9	
äer	;->1	
äff	a->115	l->2	
äft	a->30	e->1	i->1	
äg 	[->1	a->8	b->1	e->6	f->2	g->2	h->2	i->2	k->1	m->3	o->2	s->1	t->1	ä->1	å->1	
äg,	 ->16	
äg.	A->1	B->1	D->1	E->1	J->1	M->2	O->1	V->1	
äg:	 ->1	
ägN	ä->1	
äga	 ->185	,->16	.->3	:->4	g->6	n->13	r->43	s->5	
ägb	y->1	
ägd	 ->2	a->1	e->1	
äge	 ->9	,->1	.->2	l->8	n->32	r->125	s->3	t->19	
ägg	 ->22	"->1	,->1	.->1	a->180	e->43	i->3	n->27	s->21	
ägl	a->5	e->5	i->2	
ägm	ä->1	
ägn	a->53	e->1	i->2	
ägr	a->22	e->11	ö->1	
ägs	 ->7	e->6	k->2	n->7	o->1	t->1	
ägt	 ->11	
äka	r->6	
äke	m->1	n->9	r->324	
äkn	a->40	e->2	i->14	
äkr	a->40	i->24	
äkt	 ->7	.->1	a->12	e->5	i->3	s->6	
äl 	-->2	6->1	S->1	a->11	b->4	d->7	e->4	f->11	g->3	h->7	i->16	k->5	l->1	m->9	n->1	o->4	p->3	r->3	s->16	t->8	u->10	v->4	ä->5	å->1	ö->1	
äl,	 ->5	
äl.	A->1	D->1	F->3	J->2	M->1	S->1	
äla	 ->2	n->1	
älb	e->1	
äld	 ->1	a->1	i->23	r->7	
äle	n->5	r->2	t->9	
älf	t->3	u->1	ä->8	
älg	r->2	ö->1	
älh	a->1	
äli	g->1	
älj	a->22	e->5	n->3	
älk	l->1	o->50	ä->3	
äll	 ->2	,->2	.->2	?->1	a->178	b->1	d->80	e->604	i->56	n->71	o->39	s->37	t->26	
älm	e->2	å->2	
äln	i->12	
älp	 ->48	,->2	.->5	a->41	e->5	l->1	s->1	t->3	v->1	
äls	 ->2	a->24	i->1	k->2	n->2	o->8	t->7	
ält	 ->6	a->2	e->15	n->1	s->1	
älu	t->3	
älv	 ->39	,->5	.->4	a->70	b->5	f->3	h->1	k->21	n->3	p->1	s->16	t->5	ä->1	
ämb	e->8	
ämd	 ->6	a->9	e->5	h->1	
äme	l->1	
ämf	ö->18	
ämj	a->62	
ämk	a->2	
äml	i->109	
ämm	a->36	e->161	i->4	
ämn	 ->1	,->1	.->1	a->121	d->26	e->34	i->17	s->9	t->19	v->2	
ämp	a->136	e->1	l->61	n->80	
ämr	a->10	e->5	
äms	 ->1	i->1	t->77	
ämt	 ->17	,->3	.->1	a->7	n->1	s->1	
ämv	i->2	
än 	1->6	2->2	3->2	E->1	F->1	W->1	a->17	b->2	d->22	e->36	f->13	g->4	h->4	i->17	j->1	k->6	l->4	m->14	n->9	o->16	p->7	r->6	s->23	t->11	u->2	v->18	ä->4	å->8	
än,	 ->2	
än.	I->1	J->2	T->1	
än;	 ->1	
äna	 ->7	d->1	r->16	
änd	 ->9	,->2	.->1	a->142	b->9	e->325	i->232	l->6	n->64	p->6	r->368	s->46	å->53	
änf	ö->1	
äng	 ->5	.->1	a->27	b->1	d->30	e->56	i->3	l->23	n->44	r->62	s->5	t->15	
änh	e->47	
äni	e->1	n->1	t->12	
änk	 ->3	a->329	b->4	e->42	l->5	n->15	s->5	t->20	
änl	i->15	
änn	a->115	e->111	i->108	s->4	u->77	y->2	
äns	 ->6	a->62	c->2	e->42	f->2	k->50	l->50	n->12	o->1	p->1	t->138	v->1	y->72	ö->12	
änt	 ->50	,->3	.->2	:->1	a->97	l->20	n->7	s->13	
änv	i->35	
äpa	d->1	
äpn	a->2	i->1	
äpp	 ->2	,->1	.->1	a->9	e->6	h->1	s->1	t->3	
äpr	o->1	
är 	"->1	-->13	1->5	2->2	3->1	5->1	7->1	8->1	A->1	B->9	C->1	D->1	E->17	F->2	K->5	L->1	M->14	N->1	P->20	R->2	S->2	V->4	W->2	a->314	b->140	c->4	d->651	e->399	f->227	g->55	h->88	i->251	j->70	k->103	l->63	m->207	n->126	o->119	p->68	r->61	s->199	t->91	u->60	v->234	y->12	Ö->1	ä->34	å->5	ö->37	
är!	 ->29	.->1	D->1	E->1	J->1	
är,	 ->115	
är.	 ->3	.->1	D->10	E->2	F->4	G->1	H->1	I->1	J->11	K->1	R->1	S->3	V->8	k->1	
är:	 ->5	
är;	 ->1	
är?	D->1	H->1	J->1	
ära	 ->139	,->2	.->1	d->22	n->28	r->3	s->6	v->4	
ärb	e->1	
ärd	 ->27	,->8	.->6	;->2	a->37	e->331	i->41	l->3	o->7	s->16	
äre	 ->1	f->12	m->19	n->74	r->35	t->1	
ärf	r->1	ö->280	
ärg	,->2	a->1	
ärh	e->5	ä->1	
äri	 ->2	b->6	f->2	g->19	n->12	
ärj	a->2	
ärk	a->32	b->3	e->22	i->1	l->5	n->19	s->59	t->41	
ärl	 ->1	d->58	e->3	i->21	
ärm	a->36	e->50	i->10	n->5	
ärn	-->2	a->42	e->8	f->2	i->4	k->23	p->4	s->4	t->3	v->23	
äro	 ->1	a->1	m->1	s->1	
ärp	a->8	e->1	l->1	n->1	o->2	t->2	å->2	
ärr	 ->37	,->2	.->1	a->6	e->9	ä->1	ö->4	
ärs	 ->6	k->159	m->1	t->8	y->1	
ärt	 ->31	,->5	.->4	a->21	i->2	l->7	o->17	s->1	
äru	t->1	
ärv	 ->1	a->55	b->1	h->1	i->6	l->1	s->3	t->2	
äs 	t->1	u->1	y->1	
äsa	 ->3	
äsb	a->2	
äsc	h->2	
äsd	u->1	
äse	n->36	r->6	
äsf	r->1	
äsk	.->1	u->1	
äsn	i->2	
äso	n->1	
äss	i->31	
äst	 ->12	a->122	b->4	e->14	k->1	m->1	n->2	r->3	s->1	v->1	
ät 	d->1	k->1	m->1	o->2	s->5	
ät.	 ->1	
äta	 ->2	,->1	r->2	s->2	
äte	.->1	n->4	r->2	t->2	
äth	e->1	
äti	g->1	
äto	r->1	
äts	k->1	t->1	
ätt	 ->303	,->37	.->57	:->2	?->4	a->266	e->202	f->9	h->9	i->124	l->1	m->1	n->214	r->153	s->220	v->74	ä->1	
ätv	e->11	
äv 	m->1	
äva	 ->38	d->4	n->17	r->5	s->13	t->1	
ävd	a->27	e->4	v->1	
äve	n->275	r->46	s->1	
ävi	g->1	
ävj	a->1	
ävl	a->2	i->1	
ävn	a->4	i->10	
ävs	 ->52	,->3	.->2	
ävt	 ->2	s->2	
ävu	l->2	
äxa	 ->1	.->2	n->7	t->1	
äxe	l->3	r->7	
äxl	a->2	i->2	
äxo	r->1	
äxt	 ->7	,->2	.->2	b->1	e->10	h->7	s->3	
å "	m->1	
å -	 ->8	
å 1	0->2	3->2	4->1	9->1	
å 2	0->3	2->1	4->1	
å 3	3->1	4->1	7->1	
å 4	0->1	
å 5	 ->1	0->2	
å 7	,->1	5->1	
å 8	0->2	6->1	
å 9	0->1	5->1	
å A	l->2	s->1	t->1	
å B	S->1	a->5	e->1	
å C	E->1	S->1	
å D	a->1	
å E	G->4	U->4	r->2	u->18	
å F	l->1	ö->1	
å G	e->1	o->2	
å H	o->1	
å I	S->1	n->6	r->1	s->1	
å K	i->1	
å M	a->1	o->1	
å O	l->1	
å P	P->1	a->1	
å R	i->2	o->1	
å T	y->1	
å V	ä->2	
å a	b->1	c->1	k->4	l->42	m->1	n->41	r->15	s->3	t->353	v->26	
å b	a->11	e->38	i->7	l->11	o->10	r->12	y->2	ä->13	å->3	ö->10	
å c	e->1	i->1	r->1	
å d	a->10	e->398	i->4	j->7	o->2	r->2	u->4	y->1	ä->3	å->1	
å e	f->7	g->3	k->6	l->4	m->1	n->153	r->8	t->173	u->14	x->3	
å f	a->21	e->4	i->14	l->5	o->8	r->56	u->3	y->2	ä->6	å->12	ö->136	
å g	a->3	e->28	i->1	l->2	o->4	r->87	ä->4	å->9	ö->7	
å h	a->29	e->14	i->1	j->6	o->4	u->20	ä->8	å->1	ö->3	
å i	 ->50	a->1	c->1	d->1	g->5	h->1	l->2	m->1	n->80	r->1	t->1	
å j	a->8	o->2	u->3	ä->3	
å k	a->42	l->8	n->1	o->82	r->7	u->3	v->5	ä->3	ö->2	
å l	a->17	i->10	o->5	y->1	ä->34	å->24	ö->1	
å m	a->18	e->53	i->38	o->7	y->43	ä->2	å->46	ö->10	
å n	a->4	e->2	o->7	y->29	ä->15	å->32	ö->4	
å o	a->2	b->3	c->55	e->1	f->6	g->1	l->6	m->34	n->2	r->6	s->7	
å p	a->7	e->8	l->11	o->5	r->16	u->9	å->23	
å r	a->3	e->36	i->6	y->2	ä->17	å->10	ö->3	
å s	a->40	e->29	i->39	j->3	k->37	l->3	m->8	n->31	o->40	p->12	t->49	u->2	v->5	y->5	ä->41	å->31	
å t	a->36	e->4	i->67	j->1	o->11	r->17	v->8	y->3	ä->3	
å u	n->17	p->21	t->24	
å v	a->44	e->23	i->89	r->1	ä->38	å->26	
å y	t->3	
å z	i->2	
å Ö	s->2	
å ä	g->1	n->12	r->44	v->3	
å å	h->1	r->8	s->1	t->12	
å ö	k->2	n->2	p->6	v->6	
å, 	a->4	b->2	d->1	e->3	f->7	g->1	h->3	i->2	l->1	m->7	n->4	o->13	r->3	s->4	t->1	v->2	ä->1	
å. 	D->2	
å..	.->1	
å.A	t->2	
å.B	e->1	i->1	r->1	
å.D	e->13	o->1	ä->2	
å.E	n->1	u->2	
å.F	P->1	r->1	ö->2	
å.G	e->1	r->1	
å.H	e->2	
å.I	 ->1	n->1	
å.J	a->8	u->1	ä->1	
å.M	e->1	
å.N	i->1	o->1	ä->2	
å.O	c->1	m->1	r->1	
å.P	å->2	
å.S	l->1	o->1	
å.U	n->1	
å.V	i->4	
å.Ä	r->2	
å: 	a->1	d->2	f->2	Ö->1	å->1	
å; 	d->1	
å?.	 ->1	
å?I	n->1	
å?J	a->1	
å?S	e->1	
åba	r->2	
åbe	r->1	
åbj	u->1	
åbö	r->11	
åd 	(->1	-->1	a->2	b->1	f->3	i->1	n->1	o->5	s->3	
åd,	 ->4	
åd.	D->1	J->1	K->1	L->1	M->1	
åd?	Ä->1	
åda	 ->39	,->1	d->3	n->170	r->4	
ådd	 ->1	a->4	e->4	
åde	 ->103	,->14	.->23	:->1	;->1	?->1	f->1	n->134	r->36	t->416	
ådf	r->6	
ådg	i->26	ö->1	
ådl	i->7	
ådn	i->1	
ådr	a->1	
åds	b->1	k->20	l->3	m->3	o->20	r->1	t->1	
åel	i->6	s->8	
åen	d->136	
åer	 ->6	,->3	.->4	:->1	n->1	
ået	.->1	
åfr	e->1	
åfö	l->4	r->6	
åg 	I->1	a->18	d->6	e->2	h->1	i->2	n->3	o->1	r->1	s->3	t->1	u->2	Ö->1	ä->1	
åg,	 ->1	
åg.	E->1	
åga	 ->256	!->1	,->26	.->42	:->7	?->1	d->8	n->211	r->25	s->20	t->7	v->1	
åge	k->1	l->3	n->1	r->2	s->10	t->3	
ågi	c->3	
ågk	r->2	
ågl	a->6	ä->1	
ågn	i->8	
ågo	l->1	n->167	r->278	t->193	
ågr	a->149	u->3	ä->1	
ågs	 ->2	.->2	
ågt	 ->2	
ågv	e->1	
ågå	 ->1	e->6	r->10	t->1	
åhu	n->1	
åhä	n->6	r->1	
åhö	r->1	
åja	,->1	
åk 	f->1	p->3	t->1	
åk.	 ->1	
åka	 ->1	r->9	
åke	t->4	
åki	g->3	
åkl	a->37	i->3	
åko	m->2	
åkr	a->30	
åkt	a->1	e->1	
ål 	(->1	1->16	2->10	5->2	a->4	b->2	e->1	f->20	g->1	h->2	i->7	j->1	l->1	n->1	o->8	p->2	r->1	s->15	t->1	u->2	ä->4	
ål,	 ->17	
ål-	2->1	
ål.	B->1	D->3	E->1	F->1	H->2	I->2	J->1	K->1	M->2	N->2	Ä->1	
ål:	 ->2	
åla	 ->2	,->1	g->4	m->2	r->3	
åld	 ->2	e->14	r->3	s->6	t->2	
åle	d->44	n->18	t->30	
ålf	ö->5	
ålg	e->1	
åli	g->27	n->29	t->1	
ålk	a->1	
åll	 ->19	,->5	.->7	:->1	?->1	a->182	b->25	e->122	i->23	n->67	s->22	
ålm	e->1	
åln	i->3	
åls	d->1	e->7	k->1	s->1	t->1	ä->17	
ålu	n->4	
ålv	e->5	
ålä	g->6	
åmi	n->30	
ån 	(->21	-->2	1->7	2->1	3->1	5->3	8->1	9->1	A->10	B->5	C->3	D->2	E->29	F->6	G->4	H->2	I->5	J->1	K->5	L->3	M->1	N->3	O->1	P->7	R->1	S->6	T->6	U->2	V->1	W->2	a->36	b->14	d->99	e->43	f->45	g->4	h->7	i->3	j->4	k->37	l->9	m->23	n->6	o->23	p->21	r->17	s->27	t->25	u->22	v->19	Ö->1	ä->1	å->1	ö->4	
ån,	 ->4	
ån.	D->4	H->1	Ä->1	
åna	 ->4	d->74	n->2	r->12	s->1	
ånb	o->1	
ånd	 ->54	,->8	.->10	?->2	a->8	e->31	i->1	p->97	s->19	
åne	r->2	
ång	 ->147	"->1	,->11	.->14	a->178	d->1	e->73	f->19	k->1	l->1	m->1	n->2	r->3	s->73	t->52	v->6	å->1	
åni	n->7	
ånk	o->3	
åns	p->1	
ånt	a->2	o->1	
ånv	a->8	ä->1	
åny	o->1	
åol	j->1	
åpe	k->50	
åps	l->1	
år 	-->1	1->19	2->33	B->1	M->1	O->1	a->58	b->18	d->65	e->49	f->59	g->28	h->18	i->121	j->14	k->29	l->14	m->39	n->11	o->27	p->31	r->15	s->70	t->41	u->29	v->45	y->1	ä->8	å->9	ö->5	
år"	.->1	
år)	?->1	
år,	 ->32	
år.	 ->2	D->12	E->1	F->2	H->4	I->2	J->4	K->1	L->2	M->1	O->1	R->1	S->1	T->1	V->6	Ä->1	
år?	N->1	S->1	
åra	 ->179	,->1	n->1	r->5	s->1	t->1	
årb	a->3	e->2	
ård	 ->6	)->1	,->2	a->16	e->1	n->2	s->4	
åre	n->40	t->45	
årh	u->7	
åri	g->45	n->1	
årk	l->1	ö->1	
årl	i->8	ö->2	
årn	i->2	
års	 ->11	a->1	b->2	p->2	r->2	s->2	t->1	
årt	 ->146	,->3	.->1	a->1	i->1	u->3	
årö	v->1	
ås 	a->4	b->3	d->3	e->2	f->4	g->3	i->15	k->1	m->1	o->1	p->1	s->1	t->2	u->1	v->1	
ås,	 ->1	
ås.	D->1	F->1	L->1	
ås:	 ->1	
åsa	m->3	t->1	
åse	r->3	
åsi	k->50	
åsk	a->1	y->7	å->2	
åso	m->34	
åss	 ->1	
åst	 ->1	a->27	e->696	r->1	å->21	
åsy	f->5	
åt 	E->1	F->1	a->8	b->1	d->27	e->8	f->2	g->1	h->1	i->11	j->1	k->5	l->1	m->59	n->2	o->28	p->2	r->4	s->6	t->3	u->1	v->2	Ö->1	ä->3	å->1	
åt"	,->1	
åt,	 ->5	
åt.	D->3	F->1	H->1	J->1	K->1	N->1	V->1	
åta	 ->44	g->34	l->24	n->4	r->10	s->6	
åte	 ->1	n->7	r->278	t->1	
åtf	ö->12	
åtg	ä->240	å->1	
åti	l->1	t->3	
åtl	i->5	
åtm	i->27	
åtn	a->6	j->1	
åtr	y->3	
åts	 ->4	a->2	k->3	t->3	
ått	 ->127	,->2	.->7	a->5	f->1	o->4	s->9	
åtv	i->4	
åva	r->2	
åve	r->37	
åvi	d->3	l->1	s->3	
åvo	r->2	
åvä	l->41	
åzo	n->1	
ça 	M->5	
çoi	s->1	
ère	 ->1	
ète	 ->1	
ève	 ->1	,->1	k->1	
é -	 ->3	
é a	t->2	v->1	
é e	l->1	
é f	ö->3	
é h	a->1	
é j	a->1	
é k	o->1	
é m	e->1	
é o	c->3	m->1	
é p	e->1	
é s	o->5	
é u	t->1	
é ä	r->1	
é, 	m->1	
éav	t->1	
ébe	t->1	
ébé	 ->1	
éch	a->1	
ée,	 ->1	
éer	 ->10	,->3	.->1	n->7	
éfé	r->1	
éfö	r->2	
éko	n->1	
én 	(->2	a->6	b->3	f->3	i->1	k->1	l->1	m->1	o->15	s->2	v->2	ä->1	
én,	 ->5	
én.	H->1	M->1	W->1	
én?	V->1	
éns	 ->11	
ére	n->1	
éry	s->1	
és 	R->1	
ésy	s->2	
éta	i->1	
éun	i->2	
ête	 ->3	
êts	 ->1	
í ä	r->1	
íez	 ->1	
ínc	i->1	
ón 	C->2	i->1	t->1	v->1	
óni	o->1	
ône	-->1	
ö f	ö->2	
ö i	 ->2	
ö k	a->1	
ö m	o->1	
ö s	a->1	o->1	
ö v	i->1	
ö!D	e->1	
ö, 	f->8	h->1	l->1	s->1	u->1	
ö- 	o->2	
ö.D	e->3	å->1	
ö.M	e->1	
ö.U	n->1	
ö.V	i->1	
öan	p->1	s->2	
öar	 ->1	n->5	
öav	t->1	
öbe	l->1	s->2	
öbl	e->2	
öbo	 ->1	
öbr	o->1	
öck	e->3	
öd 	-->2	a->5	b->1	d->3	e->3	f->27	g->1	h->2	i->12	k->5	l->1	m->5	o->18	p->7	s->20	t->43	v->6	ä->2	å->2	ö->1	
öd,	 ->14	
öd.	"->1	-->1	.->1	A->2	D->12	E->1	F->2	H->5	I->2	J->3	M->2	N->1	O->1	R->1	S->1	T->1	U->1	V->2	Ä->2	Å->2	
öd;	 ->1	
öd?	-->1	
öda	 ->6	"->1	,->1	d->3	n->5	s->2	t->1	
ödb	e->1	
ödd	.->1	e->3	
öde	 ->2	,->4	.->1	?->1	l->6	m->1	n->34	p->1	r->63	s->4	t->34	
ödf	ö->1	
ödg	r->1	
ödi	g->13	n->1	r->1	
ödj	a->71	e->1	
ödm	e->1	o->1	
ödn	i->2	
ödo	r->1	s->1	ä->1	
ödp	o->1	
ödr	a->9	
öds	 ->10	d->1	f->1	i->1	p->1	y->4	
ödv	ä->125	
ödå	t->5	
öen	d->1	
öer	 ->3	n->1	
öfa	k->1	r->9	
öfr	å->4	
öft	e->11	
öfö	r->4	
ög 	a->1	b->1	f->1	g->6	i->1	k->1	n->2	p->2	s->6	
ög,	 ->1	
öga	 ->16	,->1	.->1	k->1	t->1	
öge	 ->2	l->1	r->31	
ögh	e->3	
ögl	j->1	
ögn	a->1	i->3	
ögo	n->19	
ögr	a->1	e->19	
ögs	k->1	t->28	
ögt	 ->9	,->1	.->1	e->2	i->4	
öin	f->1	
öja	 ->17	.->1	d->1	k->2	n->2	r->4	s->3	
öjd	 ->7	a->9	e->6	p->2	
öje	 ->4	l->1	r->5	t->2	v->3	
öjl	i->309	
öjn	i->2	
öjo	r->1	
öjs	 ->1	m->2	
öjt	 ->2	s->2	
ök 	a->4	b->1	i->5	o->1	s->1	
ök,	 ->3	
öka	 ->76	,->1	.->3	d->37	n->11	r->22	s->11	t->27	
öke	 ->1	.->1	n->2	r->21	t->4	
ökm	o->1	
ökn	i->43	
öko	n->6	
ökr	a->8	
öks	,->1	b->1	t->1	
ökt	 ->14	e->6	
ökv	a->1	
öl 	n->1	o->1	
öl,	 ->1	
öla	g->1	r->1	
öld	 ->1	,->1	b->1	g->1	
ölj	a->91	d->44	e->20	n->10	s->5	t->4	
öll	 ->20	.->1	s->4	
öln	 ->2	
öm 	a->2	b->1	i->1	t->1	
öm,	 ->1	
öm:	 ->1	
öma	 ->26	,->1	.->1	n->7	s->2	
ömb	a->1	
ömd	,->2	e->2	
öme	.->1	r->9	s->1	
ömi	n->1	
öml	i->2	
ömm	a->23	e->9	
ömn	i->34	
öms	 ->3	e->5	k->1	
ömt	 ->10	s->2	å->1	
ömv	ä->1	
ömä	n->2	s->11	
ömå	l->3	
ön 	N->1	e->2	f->2	h->1	i->1	o->6	p->1	s->2	t->1	v->2	ä->1	
ön!	D->1	
ön,	 ->9	
ön.	D->3	E->1	F->1	J->1	L->1	M->1	U->1	V->2	
öna	 ->13	/->1	r->2	s->3	
önb	o->1	
önd	e->7	
öne	-->1	a->1	n->3	r->2	
önh	e->1	
öni	t->1	
önk	 ->3	.->1	
öno	r->2	
öns	 ->2	a->5	g->1	k->69	t->3	
önt	 ->2	a->3	
öom	r->4	
öov	ä->1	
öp 	a->2	
öpa	 ->3	n->6	r->4	
öpe	n->1	r->14	
öpk	r->1	
öpo	l->8	
öpp	e->79	n->20	
öpr	o->4	
öps	b->1	l->1	
öpt	 ->6	e->3	
öpå	v->1	
ör 	"->6	-->7	1->17	2->7	3->2	5->2	7->2	8->1	A->4	B->6	C->2	D->3	E->75	F->5	G->2	H->1	I->4	K->7	L->2	M->1	O->1	P->4	S->3	T->8	V->1	W->2	a->1015	b->96	c->7	d->718	e->273	f->155	g->59	h->102	i->86	j->32	k->173	l->66	m->213	n->98	o->118	p->81	r->110	s->248	t->114	u->121	v->177	y->4	Ö->2	ä->39	å->39	ö->52	
ör"	.->1	
ör,	 ->32	
ör.	 ->2	(->1	.->1	D->7	E->1	F->1	H->1	J->1	K->1	M->3	V->5	
ör:	 ->3	
ör;	 ->1	
ör?	D->1	F->2	I->1	Ä->1	
öra	 ->459	,->9	.->18	?->1	k->1	l->1	n->396	r->3	s->84	
örb	a->14	e->33	i->32	j->14	l->15	r->5	u->38	ä->78	
örd	 ->6	,->1	.->2	a->50	e->82	h->1	j->11	n->1	o->4	r->165	u->3	ä->4	ö->20	
öre	 ->27	b->26	d->168	f->21	g->26	h->1	k->22	l->48	m->13	n->85	r->23	s->164	t->273	
örf	a->84	i->1	j->1	l->18	o->18	r->5	ä->3	å->1	ö->5	
örg	 ->14	l->2	r->3	ä->1	
örh	a->95	i->31	o->12	å->56	ö->1	
öri	g->21	n->21	r->1	
örj	a->124	d->1	e->2	n->4	
örk	 ->1	a->9	l->77	n->3	o->2	r->1	u->2	
örl	a->3	e->2	i->116	o->20	u->10	ä->6	å->4	
örm	e->5	i->3	o->12	y->1	å->48	ö->1	
örn	 ->2	a->1	e->10	i->7	s->1	u->14	y->49	
öro	l->2	n->3	r->78	
örp	a->6	l->21	
örr	 ->4	,->2	a->45	e->83	g->3	i->1	ä->5	å->1	
örs	 ->54	,->7	.->9	a->12	e->33	i->67	k->13	l->492	o->6	p->1	t->462	u->9	v->83	ä->60	å->1	ö->65	
ört	 ->58	,->3	.->2	e->3	i->6	j->21	n->1	r->66	s->34	v->1	y->3	ä->1	
öru	n->1	t->84	
örv	a->56	e->22	i->21	r->1	ä->54	å->6	
örä	n->74	
örå	d->1	l->3	
örö	d->5	r->2	v->3	
ös 	-->1	d->2	e->1	k->1	o->2	p->1	r->1	s->2	u->1	
ös,	 ->1	
ös.	D->1	
ösa	 ->50	,->4	.->4	r->3	s->6	
öse	k->1	r->4	s->1	
ösg	ö->1	
ösh	e->44	
ösi	d->1	
ösk	a->2	e->3	y->11	ä->2	
ösn	i->52	
ösr	y->1	
öss	 ->3	)->1	o->1	
öst	 ->31	,->3	.->2	a->97	b->1	e->81	f->7	l->1	n->57	r->6	s->1	t->1	u->2	v->3	ö->1	
ösy	n->6	
öt 	9->1	a->1	d->1	h->1	l->1	t->4	v->1	
öt.	D->1	
öta	 ->17	n->1	r->1	s->1	
öte	 ->13	b->1	n->4	r->90	s->6	t->21	
ötf	å->1	
ötk	ö->3	
ötr	a->1	
öts	 ->6	.->1	e->5	k->1	l->4	
ött	 ->16	.->3	a->4	e->11	k->1	r->1	s->4	
öut	s->1	
öva	 ->26	d->2	n->1	r->7	s->9	t->2	
övd	e->2	
öve	r->747	
övi	t->1	
övl	a->1	i->1	
övn	i->12	
övo	å->1	
övr	a->3	i->65	
övs	 ->20	,->2	.->5	k->1	t->1	
övt	 ->3	s->1	
övä	n->7	r->3	
öw 	f->1	
öy 	-->1	
ööw	 ->1	
øn,	 ->2	
ørg	e->2	
ühr	k->1	
ünc	h->1	
ürk	d->1	
üss	e->4	
